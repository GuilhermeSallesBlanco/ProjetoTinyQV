// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Sun Jan 11 17:38:13 2026
//
// Verilog Description of module tinyQV_top
//

module tinyQV_top (clk, rst_n, ui_in, uo_out) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(8[8:18])
    input clk;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    input rst_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(10[20:25])
    input [7:0]ui_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    output [7:0]uo_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    wire GND_net, VCC_net, rst_n_c, ui_in_c_7, ui_in_c_6, ui_in_c_5, 
        ui_in_c_4, ui_in_c_3, ui_in_c_2, ui_in_c_1, ui_in_c_0, uo_out_c_7, 
        uo_out_c_6, uo_out_c_5, uo_out_c_4, uo_out_c_3, uo_out_c_2, 
        uo_out_c_1, uo_out_c_0, rst_reg_n;
    wire [3:0]qspi_data_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(34[16:28])
    wire [3:0]qspi_data_oe;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(36[16:28])
    
    wire qspi_ram_a_select, qspi_ram_b_select;
    wire [27:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    wire [31:0]data_to_write;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(56[17:30])
    wire [31:0]data_from_read;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(59[16:30])
    wire [3:0]debug_rd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(75[16:24])
    
    wire debug_uart_txd;
    wire [7:6]gpio_out_sel;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(79[16:28])
    wire [3:0]connect_peripheral;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(81[15:33])
    
    wire debug_register_data;
    wire [3:0]debug_rd_r;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(85[15:25])
    
    wire debug_uart_tx_start;
    wire [7:0]peri_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(95[16:24])
    wire [31:0]peri_data_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(96[17:30])
    wire [7:0]ui_in_sync0;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(101[15:26])
    wire [7:0]ui_in_sync;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(102[15:25])
    wire [7:0]time_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(238[15:25])
    wire [3:0]qspi_data_in_3__N_1;
    wire [3:0]qspi_data_out_3__N_5;
    wire [1:0]gpio_out_sel_7__N_13;
    wire [24:0]addr_adj_3354;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(23[16:20])
    
    wire n39;
    wire [31:0]addr_24__N_228;
    wire [31:0]writing_N_164;
    
    wire n57, debug_instr_valid, debug_stop_txn;
    wire [23:1]instr_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(56[15:25])
    wire [1:0]qv_data_write_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(64[15:30])
    wire [1:0]qv_data_read_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(65[15:29])
    
    wire rst_reg_n_adj_3302, data_out_hold, data_ready_r, clk_c_enable_341, 
        clk_c_enable_66, n24289, clk_c_enable_340, clk_c_enable_342, 
        n24253, n2, n3, n3_adj_3303, n2_adj_3304, n24288, n24287, 
        n24252, n27757, n24286, n24285, clk_c_enable_143, n24284, 
        n24251, n24250, n28957, n31883, n17920;
    wire [7:0]\uo_out_from_user_peri[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(59[17:38])
    wire [12:0]baud_divider_adj_3410;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(36[31:43])
    
    wire n24283, n48, n24249, led_state, n32622, n4251, n33, n54, 
        n4501, n30, n51;
    wire [4:0]\gpio_out_func_sel[0] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    wire [4:0]\gpio_out_func_sel[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    wire [4:0]\gpio_out_func_sel[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    wire [4:0]\gpio_out_func_sel[3] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    wire [4:0]\gpio_out_func_sel[4] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    wire [4:0]\gpio_out_func_sel[5] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    wire [4:0]\gpio_out_func_sel[6] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    wire [4:0]\gpio_out_func_sel[7] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    
    wire n4503, data_ready_r_N_2823, n48_adj_3305, n44, n24282, n45, 
        n32548, n24281;
    wire [31:0]data_from_peri_31__N_2415;
    
    wire n31795, n57_adj_3306, n42, clk_c_enable_208;
    wire [31:0]data_from_user_peri_1__31__N_2455;
    
    wire n6142, n24248, n6218, n39_adj_3307;
    wire [12:0]cycle_counter;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(43[25:38])
    wire [3:0]fsm_state;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(47[11:20])
    
    wire next_bit, n36, n33_adj_3308, n24224, n40, uart_txd_N_3005, 
        n30_adj_3309;
    wire [31:0]instr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(47[17:22])
    
    wire n8880;
    wire [31:0]imm;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(100[16:19])
    wire [2:1]instr_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(113[15:24])
    wire [3:0]rd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(119[15:17])
    wire [31:0]pc;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(128[17:19])
    wire [31:0]next_pc_for_core;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(129[17:33])
    wire [23:1]return_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(135[17:28])
    wire [3:1]instr_write_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(152[15:33])
    
    wire was_early_branch;
    wire [15:0]\instr_data[0] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]\instr_data[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]\instr_data[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]\instr_data[3] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [23:1]early_branch_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[17:34])
    
    wire n29831, n10672, n34285, n24280, n54_adj_3310, n32615, n51_adj_3311, 
        n26838, n45_adj_3312, n60, n8109, n24247, n24223, n24216, 
        n24246, n15569, n26692, n24275, n32614, n66, n8854, n66_adj_3313, 
        n24274, n7, n32610, n24273, clk_c_enable_50, n10944;
    wire [20:0]pc_23__N_911;
    
    wire n24221, n24272;
    wire [22:0]instr_addr_23__N_318;
    
    wire qspi_write_done, data_stall, instr_active_N_2106, n24271, n32524, 
        n31796, n8177, n31794, n31793, n31792, n31791, n31790, 
        n31789, continue_txn_N_2131, data_stall_N_2158, n29, n26870, 
        n16810, n16811;
    wire [7:0]uart_rx_buf_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(98[15:31])
    
    wire n24270, n765, n32544, n24244, n24222, n24215, n2191, 
        n2150, n2211, n2594, n24269, n24268, n2130, n2196;
    wire [1:0]cycle;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(58[15:20])
    wire [3:0]mul_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(138[16:23])
    
    wire n6220, instr_complete_N_1647, n24267, n24316, n29631, n24266, 
        n24217, n24315, n24243, n24314, n24242, n24313, n24241, 
        n24218, n24312, n24219, n24311, n24310, n24240, n762, 
        n24239, n24238, n36_adj_3314, n24308, n28319;
    wire [3:0]csr_read_3__N_1447;
    
    wire n10737, n24307, n41, n43, n24306, n29549, n24305, n31706, 
        n24237, n24304, n5169, n32851, n32850, n24303, clk_c_enable_432, 
        n32842, n24236, n29491, n27888, n24214, n32836, n32835, 
        n32834, n32833, n24259, n17165, n32832, n24302, n24301, 
        n4513, n29884, n45_adj_3315, n32825, clk_c_enable_543, clk_c_enable_154, 
        n29866, n32822, n24300, n24258, n32819, n24257, n24256, 
        n24299, n32818;
    wire [2:0]fsm_state_adj_3463;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(82[15:24])
    
    wire is_writing;
    wire [23:0]addr_adj_3464;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(84[31:35])
    
    wire spi_clk_pos, stop_txn_reg, stop_txn_now_N_2363, n24298, is_writing_N_2331, 
        n24255, n24254, n32874, n24297, n42_adj_3317, n24296, n26811, 
        n32802, n32801, n26691, n32568, clk_c_enable_286, n1072, 
        n63, n32791, clk_c_enable_283, n46;
    wire [12:0]cycle_counter_adj_3482;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(43[25:38])
    wire [3:0]fsm_state_adj_3483;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(47[11:20])
    
    wire next_bit_adj_3332, n38, clk_c_enable_495, n39_adj_3333, n63_adj_3334, 
        n42_adj_3335;
    wire [12:0]cycle_counter_adj_3505;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(39[25:38])
    
    wire next_bit_adj_3349;
    wire [31:0]next_fsm_state_3__N_3046;
    
    wire n28259, n31351, n31350, n1152, n32251, n32771, clk_c_enable_519, 
        clk_c_enable_285, n60_adj_3350, clk_c_enable_354;
    wire [15:0]accum;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(104[22:27])
    wire [19:0]next_accum;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[23:33])
    wire [19:0]d_3__N_1868;
    
    wire n32766, n29357, n24295, n24294, n32763, n28077, n24293, 
        n24292, n29337, n29335, n29333, n32761, n32759, n32756, 
        n32755, n29707, n24290, n16420, n16419, n16417, n12, n29293, 
        n27178, n19, n4, n32745, n14, n14_adj_3351, n29738, n32523, 
        n32737, n32734, n29263, n32522, n32730, n32729, n32728, 
        n26116, n32727, n32725, n32723, n32720, n32520, n32521, 
        n27124, n27120, n32714, n32552, n32710, n32072, n32706, 
        n29741, n32060, n32700, n32695, n32694, n26856, n32693, 
        n32892, n29127, n32685, n32681, n32672, n32660, n27931, 
        n28111, n32656, n32655, n32654, n26466, n11, n32650, n29887, 
        n32642, n32640, n32638;
    
    VHI i2 (.Z(VCC_net));
    INV i30011 (.A(clk_c), .Z(clk_N_45));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    FD1S3AX debug_rd_r_i0 (.D(debug_rd[0]), .CK(clk_c), .Q(debug_rd_r[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(257[12] 259[8])
    defparam debug_rd_r_i0.GSR = "DISABLED";
    FD1S3AX rst_reg_n_53 (.D(rst_n_c), .CK(clk_N_45), .Q(rst_reg_n));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(31[12:46])
    defparam rst_reg_n_53.GSR = "DISABLED";
    FD1S3AX ui_in_sync0_i6 (.D(ui_in_c_6), .CK(clk_c), .Q(ui_in_sync0[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i6.GSR = "DISABLED";
    CCU2C _add_1_5098_add_4_4 (.A0(baud_divider_adj_3410[1]), .B0(cycle_counter_adj_3482[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[2]), .B1(cycle_counter_adj_3482[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24246), .COUT(n24247));
    defparam _add_1_5098_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_5098_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_5098_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_5098_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_7 (.A0(early_branch_addr[7]), .B0(was_early_branch), 
          .C0(pc[7]), .D0(VCC_net), .A1(early_branch_addr[8]), .B1(was_early_branch), 
          .C1(pc[8]), .D1(VCC_net), .CIN(n24282), .COUT(n24283), .S0(instr_addr_23__N_318[6]), 
          .S1(instr_addr_23__N_318[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_7.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_7.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_7.INJECT1_1 = "NO";
    \peripherals_min(CLOCK_MHZ=25)  i_peripherals (.clk_c(clk_c), .clk_c_enable_432(clk_c_enable_432), 
            .\data_to_write[3] (data_to_write[3]), .\peri_data_out[0] (peri_data_out[0]), 
            .data_out_hold(data_out_hold), .n32706(n32706), .\data_to_write[1] (data_to_write[1]), 
            .\peri_data_out[1] (peri_data_out[1]), .n15569(n15569), .\peri_data_out[2] (peri_data_out[2]), 
            .n26116(n26116), .\peri_data_out[3] (peri_data_out[3]), .\peri_data_out[4] (peri_data_out[4]), 
            .clk_c_enable_50(clk_c_enable_50), .\peri_data_out[5] (peri_data_out[5]), 
            .n3(n3), .n32520(n32520), .\addr[7] (addr[7]), .n2(n2), 
            .\peri_data_out[6] (peri_data_out[6]), .n3_adj_47(n3_adj_3303), 
            .n28077(n28077), .\addr[10] (addr[10]), .n32851(n32851), .\addr[6] (addr[6]), 
            .n12(n12), .\gpio_out_func_sel[0] ({\gpio_out_func_sel[0] }), 
            .\data_to_write[4] (data_to_write[4]), .n32835(n32835), .n32836(n32836), 
            .\addr[2] (addr[2]), .n29(n29), .\data_to_write[0] (data_to_write[0]), 
            .\peri_data_out[7] (peri_data_out[7]), .\peri_data_out[8] (peri_data_out[8]), 
            .baud_divider({baud_divider_adj_3410}), .\gpio_out_func_sel[6][2] (\gpio_out_func_sel[6] [2]), 
            .\data_to_write[2] (data_to_write[2]), .\peri_data_out[9] (peri_data_out[9]), 
            .\gpio_out_func_sel[2][4] (\gpio_out_func_sel[2] [4]), .\gpio_out_func_sel[7][4] (\gpio_out_func_sel[7] [4]), 
            .clk_c_enable_154(clk_c_enable_154), .\gpio_out_func_sel[1][4] (\gpio_out_func_sel[1] [4]), 
            .\gpio_out_func_sel[1][2] (\gpio_out_func_sel[1] [2]), .uo_out_c_1(uo_out_c_1), 
            .\gpio_out_func_sel[4] ({Open_0, Open_1, \gpio_out_func_sel[4] [2], 
            Open_2, Open_3}), .n2_adj_48(n2_adj_3304), .n26856(n26856), 
            .\gpio_out_func_sel[7][2] (\gpio_out_func_sel[7] [2]), .\uo_out_from_user_peri[1] ({Open_4, 
            Open_5, Open_6, Open_7, Open_8, Open_9, Open_10, \uo_out_from_user_peri[1] [0]}), 
            .\peri_data_out[10] (peri_data_out[10]), .\gpio_out_func_sel[3][4] (\gpio_out_func_sel[3] [4]), 
            .\gpio_out_func_sel[3][2] (\gpio_out_func_sel[3] [2]), .clk_c_enable_283(clk_c_enable_283), 
            .\gpio_out_func_sel[2][2] (\gpio_out_func_sel[2] [2]), .\peri_data_out[11] (peri_data_out[11]), 
            .\peri_data_out[12] (peri_data_out[12]), .\gpio_out_func_sel[5][4] (\gpio_out_func_sel[5] [4]), 
            .\gpio_out_func_sel[6][4] (\gpio_out_func_sel[6] [4]), .\gpio_out_func_sel[5][2] (\gpio_out_func_sel[5] [2]), 
            .\gpio_out_func_sel[4][4] (\gpio_out_func_sel[4] [4]), .clk_c_enable_354(clk_c_enable_354), 
            .data_ready_r(data_ready_r), .rst_reg_n(rst_reg_n), .data_ready_r_N_2823(data_ready_r_N_2823), 
            .\addr[4] (addr[4]), .\addr[3] (addr[3]), .n32818(n32818), 
            .n10944(n10944), .\uo_out_from_user_peri[1][2] (\uo_out_from_user_peri[1] [2]), 
            .\uo_out_from_user_peri[1][5] (\uo_out_from_user_peri[1] [5]), 
            .\data_to_write[5] (data_to_write[5]), .\uo_out_from_user_peri[1][6] (\uo_out_from_user_peri[1] [6]), 
            .\data_to_write[6] (data_to_write[6]), .\data_to_write[7] (data_to_write[7]), 
            .\gpio_out_sel[7] (gpio_out_sel[7]), .uo_out_c_7(uo_out_c_7), 
            .\ui_in_sync[2] (ui_in_sync[2]), .n31883(n31883), .n26838(n26838), 
            .\data_from_user_peri_1__31__N_2455[2] (data_from_user_peri_1__31__N_2455[2]), 
            .led_state(led_state), .\addr[1] (addr[1]), .n27888(n27888), 
            .n32693(n32693), .n32729(n32729), .n8854(n8854), .n32819(n32819), 
            .\debug_rd_r[0] (debug_rd_r[0]), .debug_register_data(debug_register_data), 
            .uo_out_c_2(uo_out_c_2), .\ui_in_sync[1] (ui_in_sync[1]), .n32761(n32761), 
            .\ui_in_sync[3] (ui_in_sync[3]), .\ui_in_sync[4] (ui_in_sync[4]), 
            .n31794(n31794), .\ui_in_sync[0] (ui_in_sync[0]), .\data_from_user_peri_1__31__N_2455[0] (data_from_user_peri_1__31__N_2455[0]), 
            .n32723(n32723), .n32727(n32727), .n32728(n32728), .n32720(n32720), 
            .n32737(n32737), .\peri_out[3] (peri_out[3]), .\data_from_user_peri_1__31__N_2455[7] (data_from_user_peri_1__31__N_2455[7]), 
            .\peri_out[4] (peri_out[4]), .n32801(n32801), .n8109(n8109), 
            .n32700(n32700), .\peri_out[5] (peri_out[5]), .\peri_out[6] (peri_out[6]), 
            .\data_from_peri_31__N_2415[0] (data_from_peri_31__N_2415[0]), 
            .\data_to_write[12] (data_to_write[12]), .\data_to_write[11] (data_to_write[11]), 
            .\data_to_write[10] (data_to_write[10]), .\data_to_write[9] (data_to_write[9]), 
            .\data_to_write[8] (data_to_write[8]), .\ui_in_sync[7] (ui_in_sync[7]), 
            .n31706(n31706), .\uart_rx_buf_data[2] (uart_rx_buf_data[2]), 
            .\uart_rx_buf_data[3] (uart_rx_buf_data[3]), .\uart_rx_buf_data[4] (uart_rx_buf_data[4]), 
            .\uart_rx_buf_data[5] (uart_rx_buf_data[5]), .\uart_rx_buf_data[6] (uart_rx_buf_data[6]), 
            .\uart_rx_buf_data[7] (uart_rx_buf_data[7]), .\next_fsm_state_3__N_3046[3] (next_fsm_state_3__N_3046[3]), 
            .n31795(n31795), .n31796(n31796), .\addr[5] (addr[5]), .\addr[0] (addr[0]), 
            .n32695(n32695), .n32730(n32730), .n26870(n26870), .n32725(n32725), 
            .qv_data_write_n({qv_data_write_n}), .n32710(n32710), .\imm[6] (imm[6]), 
            .\csr_read_3__N_1447[2] (csr_read_3__N_1447[2]), .n29866(n29866), 
            .n29491(n29491), .cycle_counter({cycle_counter_adj_3482}), .n72({n30, 
            n33, n36_adj_3314, n39, n42_adj_3317, n45_adj_3312, n48, 
            n51_adj_3311, n54_adj_3310, n57_adj_3306, n60_adj_3350, 
            n63_adj_3334, n66}), .n32791(n32791), .fsm_state({fsm_state_adj_3483}), 
            .next_bit(next_bit_adj_3332), .n27757(n27757), .n32763(n32763), 
            .n32251(n32251), .GND_net(GND_net), .VCC_net(VCC_net), .cycle_counter_adj_65({cycle_counter_adj_3505}), 
            .next_bit_adj_62(next_bit_adj_3349), .debug_stop_txn(debug_stop_txn), 
            .instr_active_N_2106(instr_active_N_2106), .stop_txn_reg(stop_txn_reg), 
            .n32755(n32755), .stop_txn_now_N_2363(stop_txn_now_N_2363), 
            .clk_c_enable_208(clk_c_enable_208), .n32714(n32714), .qspi_write_done(qspi_write_done), 
            .n10672(n10672), .spi_clk_pos(spi_clk_pos), .n28259(n28259), 
            .next_bit_adj_63(next_bit), .n32622(n32622), .uart_txd_N_3005(uart_txd_N_3005), 
            .clk_c_enable_495(clk_c_enable_495), .n32832(n32832), .\fsm_state[0]_adj_64 (fsm_state[0]), 
            .clk_c_enable_143(clk_c_enable_143), .n762(n762), .clk_c_enable_519(clk_c_enable_519), 
            .n8177(n8177), .n32524(n32524), .n29357(n29357), .n46(n46), 
            .clk_c_enable_286(clk_c_enable_286), .instr_complete_N_1647(instr_complete_N_1647), 
            .n28957(n28957), .n32771(n32771), .n27178(n27178), .n29549(n29549), 
            .n6142(n6142), .n28319(n28319), .n32681(n32681), .n27931(n27931), 
            .n1072(n1072), .clk_c_enable_543(clk_c_enable_543), .qv_data_read_n({qv_data_read_n}), 
            .n26691(n26691), .\qspi_data_in[1] (qspi_data_in[1]), .\qspi_data_out_3__N_5[1] (qspi_data_out_3__N_5[1]), 
            .n26692(n26692)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(161[46] 180[6])
    CCU2C _add_1_5110_add_4_5 (.A0(early_branch_addr[5]), .B0(was_early_branch), 
          .C0(pc[5]), .D0(VCC_net), .A1(early_branch_addr[6]), .B1(was_early_branch), 
          .C1(pc[6]), .D1(VCC_net), .CIN(n24281), .COUT(n24282), .S0(instr_addr_23__N_318[4]), 
          .S1(instr_addr_23__N_318[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_5.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_5.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_3 (.A0(pc[3]), .B0(was_early_branch), .C0(early_branch_addr[3]), 
          .D0(instr_write_offset[3]), .A1(early_branch_addr[4]), .B1(was_early_branch), 
          .C1(pc[4]), .D1(VCC_net), .CIN(n24280), .COUT(n24281), .S0(instr_addr_23__N_318[2]), 
          .S1(instr_addr_23__N_318[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_5110_add_4_3.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(was_early_branch), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n24280));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5110_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_5110_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_5098_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(baud_divider_adj_3410[0]), .B1(cycle_counter_adj_3482[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n24246));
    defparam _add_1_5098_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_5098_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_5098_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_5098_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_20 (.A0(d_3__N_1868[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_3__N_1868[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24244), .S0(next_accum[18]), .S1(next_accum[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_add_4_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_add_4_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_18 (.A0(d_3__N_1868[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_3__N_1868[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24243), .COUT(n24244), .S0(next_accum[16]), 
          .S1(next_accum[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_add_4_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_add_4_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_16 (.A0(accum[14]), .B0(d_3__N_1868[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[15]), .B1(d_3__N_1868[15]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24242), .COUT(n24243), .S0(next_accum[14]), 
          .S1(next_accum[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_14 (.A0(accum[12]), .B0(d_3__N_1868[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[13]), .B1(d_3__N_1868[13]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24241), .COUT(n24242), .S0(next_accum[12]), 
          .S1(next_accum[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_12 (.A0(accum[10]), .B0(d_3__N_1868[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[11]), .B1(d_3__N_1868[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24240), .COUT(n24241), .S0(next_accum[10]), 
          .S1(next_accum[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_10 (.A0(accum[8]), .B0(d_3__N_1868[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[9]), .B1(d_3__N_1868[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24239), .COUT(n24240), .S0(next_accum[8]), 
          .S1(next_accum[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_21 (.A0(pc[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[23]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24275), .S0(next_pc_for_core[22]), .S1(next_pc_for_core[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_8 (.A0(accum[6]), .B0(d_3__N_1868[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[7]), .B1(d_3__N_1868[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24238), .COUT(n24239), .S0(next_accum[6]), 
          .S1(next_accum[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_19 (.A0(pc[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[21]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24274), .COUT(n24275), .S0(next_pc_for_core[20]), .S1(next_pc_for_core[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_6 (.A0(accum[4]), .B0(d_3__N_1868[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[5]), .B1(d_3__N_1868[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24237), .COUT(n24238), .S0(next_accum[4]), 
          .S1(next_accum[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_4 (.A0(accum[2]), .B0(d_3__N_1868[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[3]), .B1(d_3__N_1868[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24236), .COUT(n24237), .S0(mul_out[2]), 
          .S1(mul_out[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_17 (.A0(pc[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[19]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24273), .COUT(n24274), .S0(next_pc_for_core[18]), .S1(next_pc_for_core[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_2 (.A0(accum[0]), .B0(d_3__N_1868[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[1]), .B1(d_3__N_1868[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n24236), .S1(mul_out[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_add_4_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_15 (.A0(pc[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24272), .COUT(n24273), .S0(next_pc_for_core[16]), .S1(next_pc_for_core[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_13 (.A0(pc[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[15]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24271), .COUT(n24272), .S0(next_pc_for_core[14]), .S1(next_pc_for_core[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_13.INJECT1_1 = "NO";
    LUT4 i14840_2_lut (.A(data_to_write[6]), .B(n762), .Z(gpio_out_sel_7__N_13[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(209[13:93])
    defparam i14840_2_lut.init = 16'h8888;
    CCU2C _add_1_5104_add_4_11 (.A0(pc[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[13]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24270), .COUT(n24271), .S0(next_pc_for_core[12]), .S1(next_pc_for_core[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_9 (.A0(pc[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[11]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24269), .COUT(n24270), .S0(next_pc_for_core[10]), .S1(next_pc_for_core[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_7 (.A0(pc[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[9]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24268), .COUT(n24269), .S0(next_pc_for_core[8]), .S1(next_pc_for_core[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_7.INJECT1_1 = "NO";
    CCU2C time_count_3542_add_4_9 (.A0(time_count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24224), .S0(n38));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542_add_4_9.INIT0 = 16'haaa0;
    defparam time_count_3542_add_4_9.INIT1 = 16'h0000;
    defparam time_count_3542_add_4_9.INJECT1_0 = "NO";
    defparam time_count_3542_add_4_9.INJECT1_1 = "NO";
    CCU2C time_count_3542_add_4_7 (.A0(time_count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24223), .COUT(n24224), .S0(n40), .S1(n39_adj_3333));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542_add_4_7.INIT0 = 16'haaa0;
    defparam time_count_3542_add_4_7.INIT1 = 16'haaa0;
    defparam time_count_3542_add_4_7.INJECT1_0 = "NO";
    defparam time_count_3542_add_4_7.INJECT1_1 = "NO";
    CCU2C time_count_3542_add_4_5 (.A0(time_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24222), .COUT(n24223), .S0(n42_adj_3335), 
          .S1(n41));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542_add_4_5.INIT0 = 16'haaa0;
    defparam time_count_3542_add_4_5.INIT1 = 16'haaa0;
    defparam time_count_3542_add_4_5.INJECT1_0 = "NO";
    defparam time_count_3542_add_4_5.INJECT1_1 = "NO";
    CCU2C time_count_3542_add_4_3 (.A0(time_count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24221), .COUT(n24222), .S0(n44), .S1(n43));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542_add_4_3.INIT0 = 16'haaa0;
    defparam time_count_3542_add_4_3.INIT1 = 16'haaa0;
    defparam time_count_3542_add_4_3.INJECT1_0 = "NO";
    defparam time_count_3542_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5101_add_4_7 (.A0(cycle_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24216), .COUT(n24217), .S0(n51), .S1(n48_adj_3305));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5101_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_5101_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_5101_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5101_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_5101_add_4_13 (.A0(cycle_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24219), .S0(n33_adj_3308), .S1(n30_adj_3309));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5101_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_5101_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_5101_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5101_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_5101_add_4_3 (.A0(cycle_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24214), .COUT(n24215), .S0(n63), .S1(n60));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5101_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_5101_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_5101_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5101_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5101_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycle_counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n24214), .S1(n66_adj_3313));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5101_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5101_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_5101_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5101_add_4_1.INJECT1_1 = "NO";
    CCU2C time_count_3542_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n24221), .S1(n45_adj_3315));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542_add_4_1.INIT0 = 16'h0000;
    defparam time_count_3542_add_4_1.INIT1 = 16'h555f;
    defparam time_count_3542_add_4_1.INJECT1_0 = "NO";
    defparam time_count_3542_add_4_1.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync0_i5 (.D(ui_in_c_5), .CK(clk_c), .Q(ui_in_sync0[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i5.GSR = "DISABLED";
    LUT4 i15156_4_lut (.A(n5169), .B(data_from_read[31]), .C(peri_data_out[0]), 
         .D(n32685), .Z(data_from_read[0])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i15156_4_lut.init = 16'hfcee;
    LUT4 i1_4_lut (.A(peri_data_out[7]), .B(n27124), .C(n7), .D(n32685), 
         .Z(data_from_read[7])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut.init = 16'hfefc;
    LUT4 i1_4_lut_adj_618 (.A(n32685), .B(n19), .C(peri_data_out[3]), 
         .D(n4), .Z(data_from_read[3])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_618.init = 16'heeec;
    GSR GSR_INST (.GSR(n32802));
    LUT4 i1_4_lut_adj_619 (.A(n32685), .B(n19), .C(peri_data_out[2]), 
         .D(n4), .Z(data_from_read[2])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_619.init = 16'heeec;
    LUT4 i1_4_lut_adj_620 (.A(peri_data_out[6]), .B(n27120), .C(n7), .D(n32685), 
         .Z(data_from_read[6])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_620.init = 16'hfefc;
    CCU2C _add_1_5104_add_4_5 (.A0(pc[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[7]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24267), .COUT(n24268), .S0(next_pc_for_core[6]), .S1(next_pc_for_core[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_621 (.A(n32685), .B(n19), .C(peri_data_out[5]), 
         .D(n4), .Z(data_from_read[5])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_621.init = 16'heeec;
    LUT4 i1_4_lut_adj_622 (.A(n32685), .B(n19), .C(peri_data_out[1]), 
         .D(n4), .Z(data_from_read[1])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_622.init = 16'heeec;
    LUT4 i1_4_lut_adj_623 (.A(n32685), .B(n19), .C(peri_data_out[12]), 
         .D(n4), .Z(data_from_read[12])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_623.init = 16'heeec;
    LUT4 i1_4_lut_adj_624 (.A(n32685), .B(n19), .C(peri_data_out[8]), 
         .D(n4), .Z(data_from_read[8])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_624.init = 16'heeec;
    FD1S3IX time_count_3542__i0 (.D(n45_adj_3315), .CK(clk_c), .CD(n765), 
            .Q(time_count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542__i0.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_625 (.A(n32685), .B(n19), .C(peri_data_out[4]), 
         .D(n4), .Z(data_from_read[4])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_625.init = 16'heeec;
    CCU2C _add_1_5104_add_4_3 (.A0(pc[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[5]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24266), .COUT(n24267), .S0(next_pc_for_core[4]), .S1(next_pc_for_core[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5101_add_4_5 (.A0(cycle_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24215), .COUT(n24216), .S0(n57), .S1(n54));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5101_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_5101_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_5101_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5101_add_4_5.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync0_i4 (.D(ui_in_c_4), .CK(clk_c), .Q(ui_in_sync0[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i4.GSR = "DISABLED";
    CCU2C _add_1_5104_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[3]), .B1(n32842), .C1(instr_len[2]), 
          .D1(pc[2]), .COUT(n24266), .S1(next_pc_for_core[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5104_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5104_add_4_1.INIT1 = 16'h566a;
    defparam _add_1_5104_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_1.INJECT1_1 = "NO";
    LUT4 gnd_bdd_2_lut_28651 (.A(n31350), .B(rst_reg_n_adj_3302), .Z(n31351)) /* synthesis lut_function=(A (B)) */ ;
    defparam gnd_bdd_2_lut_28651.init = 16'h8888;
    FD1S3AX ui_in_sync0_i3 (.D(ui_in_c_3), .CK(clk_c), .Q(ui_in_sync0[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i3.GSR = "DISABLED";
    LUT4 rst_reg_n_bdd_4_lut (.A(cycle[0]), .B(n17920), .C(clk_c_enable_285), 
         .D(instr_complete_N_1647), .Z(n31350)) /* synthesis lut_function=(!(A (B (C))+!A (((D)+!C)+!B))) */ ;
    defparam rst_reg_n_bdd_4_lut.init = 16'h2a6a;
    FD1P3AX gpio_out_sel_i7 (.D(gpio_out_sel_7__N_13[1]), .SP(clk_c_enable_519), 
            .CK(clk_c), .Q(gpio_out_sel[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(204[12] 211[8])
    defparam gpio_out_sel_i7.GSR = "DISABLED";
    FD1S3AX ui_in_sync_i7 (.D(ui_in_sync0[7]), .CK(clk_c), .Q(ui_in_sync[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i7.GSR = "DISABLED";
    OB uo_out_pad_3 (.I(uo_out_c_3), .O(uo_out[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    FD1S3AX ui_in_sync_i6 (.D(ui_in_sync0[6]), .CK(clk_c), .Q(ui_in_sync[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i6.GSR = "DISABLED";
    OB uo_out_pad_4 (.I(uo_out_c_4), .O(uo_out[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_5 (.I(uo_out_c_5), .O(uo_out[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_6 (.I(uo_out_c_6), .O(uo_out[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    LUT4 i1530_4_lut (.A(pc[2]), .B(n2191), .C(n34285), .D(pc[1]), .Z(n2150)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i1530_4_lut.init = 16'hcac0;
    FD1S3AX ui_in_sync_i5 (.D(ui_in_sync0[5]), .CK(clk_c), .Q(ui_in_sync[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i5.GSR = "DISABLED";
    tinyQV i_tinyqv (.rst_reg_n_adj_17(rst_reg_n_adj_3302), .clk_c(clk_c), 
           .rst_reg_n(rst_reg_n), .n32771(n32771), .instr_active_N_2106(instr_active_N_2106), 
           .n26692(n26692), .qspi_write_done(qspi_write_done), .\instr_addr_23__N_318[7] (instr_addr_23__N_318[7]), 
           .\instr_addr_23__N_318[6] (instr_addr_23__N_318[6]), .\addr[7] (addr[7]), 
           .\instr_addr_23__N_318[8] (instr_addr_23__N_318[8]), .\instr_addr_23__N_318[20] (instr_addr_23__N_318[20]), 
           .\instr_addr_23__N_318[21] (instr_addr_23__N_318[21]), .\instr_addr_23__N_318[2] (instr_addr_23__N_318[2]), 
           .\addr[3] (addr[3]), .\addr[2] (addr[2]), .\instr_addr[1] (instr_addr[1]), 
           .\addr[1] (addr[1]), .n32522(n32522), .n32755(n32755), .clk_c_enable_432(clk_c_enable_432), 
           .n26691(n26691), .n10672(n10672), .data_stall(data_stall), 
           .n29887(n29887), .n32523(n32523), .data_to_write({Open_11, 
           Open_12, Open_13, Open_14, Open_15, Open_16, Open_17, 
           Open_18, Open_19, Open_20, Open_21, Open_22, Open_23, 
           Open_24, Open_25, Open_26, Open_27, Open_28, Open_29, 
           Open_30, Open_31, Open_32, Open_33, Open_34, Open_35, 
           Open_36, Open_37, Open_38, Open_39, Open_40, Open_41, 
           data_to_write[0]}), .is_writing_N_2331(is_writing_N_2331), .\data_to_write[12] (data_to_write[12]), 
           .\data_to_write[11] (data_to_write[11]), .\data_to_write[10] (data_to_write[10]), 
           .\data_to_write[9] (data_to_write[9]), .\data_to_write[8] (data_to_write[8]), 
           .\data_to_write[7] (data_to_write[7]), .\data_to_write[6] (data_to_write[6]), 
           .\data_to_write[5] (data_to_write[5]), .\data_to_write[4] (data_to_write[4]), 
           .\data_to_write[2] (data_to_write[2]), .\addr[0] (addr[0]), .n32714(n32714), 
           .continue_txn_N_2131(continue_txn_N_2131), .data_stall_N_2158(data_stall_N_2158), 
           .n32801(n32801), .\instr_addr_23__N_318[5] (instr_addr_23__N_318[5]), 
           .\addr[6] (addr[6]), .\instr_addr_23__N_318[11] (instr_addr_23__N_318[11]), 
           .\instr_addr_23__N_318[14] (instr_addr_23__N_318[14]), .\instr_addr_23__N_318[9] (instr_addr_23__N_318[9]), 
           .\addr[10] (addr[10]), .\instr_addr_23__N_318[15] (instr_addr_23__N_318[15]), 
           .\instr_addr_23__N_318[16] (instr_addr_23__N_318[16]), .\instr_addr_23__N_318[17] (instr_addr_23__N_318[17]), 
           .\instr_addr_23__N_318[12] (instr_addr_23__N_318[12]), .\instr_addr_23__N_318[10] (instr_addr_23__N_318[10]), 
           .\instr_addr_23__N_318[13] (instr_addr_23__N_318[13]), .\instr_addr_23__N_318[3] (instr_addr_23__N_318[3]), 
           .\addr[4] (addr[4]), .is_writing(is_writing), .spi_clk_pos(spi_clk_pos), 
           .stop_txn_now_N_2363(stop_txn_now_N_2363), .\instr_addr_23__N_318[22] (instr_addr_23__N_318[22]), 
           .\instr_addr_23__N_318[4] (instr_addr_23__N_318[4]), .\addr[5] (addr[5]), 
           .\instr_addr_23__N_318[19] (instr_addr_23__N_318[19]), .\instr_addr_23__N_318[18] (instr_addr_23__N_318[18]), 
           .fsm_state({Open_42, Open_43, fsm_state_adj_3463[0]}), .clk_c_enable_340(clk_c_enable_340), 
           .n32524(n32524), .clk_c_enable_208(clk_c_enable_208), .clk_c_enable_66(clk_c_enable_66), 
           .n29884(n29884), .n27931(n27931), .n32681(n32681), .n8177(n8177), 
           .qspi_data_out_3__N_5({qspi_data_out_3__N_5}), .\qspi_data_in[3] (qspi_data_in[3]), 
           .\qspi_data_in[2] (qspi_data_in[2]), .qspi_ram_a_select(qspi_ram_a_select), 
           .qspi_ram_b_select(qspi_ram_b_select), .clk_N_45(clk_N_45), .stop_txn_reg(stop_txn_reg), 
           .n32521(n32521), .\qspi_data_oe[1] (qspi_data_oe[1]), .clk_c_enable_341(clk_c_enable_341), 
           .n1072(n1072), .debug_stop_txn(debug_stop_txn), .\writing_N_164[3] (writing_N_164[3]), 
           .n4513(n4513), .n4501(n4501), .n32833(n32833), .n26811(n26811), 
           .n4503(n4503), .\addr[20] (addr_adj_3464[20]), .\addr[22] (addr_adj_3464[22]), 
           .n6218(n6218), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
           .qspi_clk_N_56(qspi_clk_N_56), .n6220(n6220), .clk_c_enable_543(clk_c_enable_543), 
           .n28319(n28319), .n32874(n32874), .n28259(n28259), .\qspi_data_in[0] (qspi_data_in[0]), 
           .n32060(n32060), .n28111(n28111), .n32892(n32892), .\imm[17] (imm[17]), 
           .\instr[31] (instr[31]), .\imm[16] (imm[16]), .\imm[15] (imm[15]), 
           .\imm[14] (imm[14]), .\imm[13] (imm[13]), .\imm[12] (imm[12]), 
           .\imm[11] (imm[11]), .\imm[10] (imm[10]), .\imm[9] (imm[9]), 
           .\imm[8] (imm[8]), .\imm[7] (imm[7]), .\imm[6] (imm[6]), .\imm[5] (imm[5]), 
           .\imm[4] (imm[4]), .\imm[3] (imm[3]), .\imm[2] (imm[2]), .\imm[1] (imm[1]), 
           .was_early_branch(was_early_branch), .\rd[0] (rd[0]), .qv_data_read_n({qv_data_read_n}), 
           .n29738(n29738), .\instr_data[3][0] (\instr_data[3] [0]), .\instr_addr_23__N_318[0] (instr_addr_23__N_318[0]), 
           .n32656(n32656), .n26116(n26116), .debug_instr_valid(debug_instr_valid), 
           .n32851(n32851), .n32835(n32835), .n32723(n32723), .\gpio_out_func_sel[5][2] (\gpio_out_func_sel[5] [2]), 
           .\gpio_out_func_sel[7][2] (\gpio_out_func_sel[7] [2]), .\instr_len[2] (instr_len[2]), 
           .\pc[2] (pc[2]), .\pc[1] (pc[1]), .n2196(n2196), .n32727(n32727), 
           .n2191(n2191), .n32640(n32640), .n32548(n32548), .n32734(n32734), 
           .n32836(n32836), .n27888(n27888), .\gpio_out_func_sel[5][4] (\gpio_out_func_sel[5] [4]), 
           .\gpio_out_func_sel[7][4] (\gpio_out_func_sel[7] [4]), .n29831(n29831), 
           .n32655(n32655), .n32544(n32544), .\instr_write_offset[3] (instr_write_offset[3]), 
           .n2150(n2150), .n2130(n2130), .n4251(n4251), .n32685(n32685), 
           .n19(n19), .n32660(n32660), .\peri_data_out[11] (peri_data_out[11]), 
           .n4(n4), .\peri_data_out[10] (peri_data_out[10]), .n32642(n32642), 
           .\peri_data_out[9] (peri_data_out[9]), .n31796(n31796), .n31795(n31795), 
           .n32520(n32520), .n32654(n32654), .\pc[7] (pc[7]), .\pc[15] (pc[15]), 
           .n32842(n32842), .\next_pc_for_core[6] (next_pc_for_core[6]), 
           .\pc[3] (pc[3]), .\pc[11] (pc[11]), .n32251(n32251), .n31706(n31706), 
           .clk_c_enable_285(clk_c_enable_285), .n28957(n28957), .n34285(n34285), 
           .\pc[6] (pc[6]), .\pc[14] (pc[14]), .\pc[10] (pc[10]), .n3(n3), 
           .n3_adj_18(n3_adj_3303), .n32638(n32638), .n29707(n29707), 
           .qv_data_write_n({qv_data_write_n}), .\addr[27] (addr[27]), .n32850(n32850), 
           .\imm[21] (imm[21]), .\imm[20] (imm[20]), .\next_pc_for_core[9] (next_pc_for_core[9]), 
           .\next_pc_for_core[13] (next_pc_for_core[13]), .\pc[5] (pc[5]), 
           .\pc[13] (pc[13]), .\pc[9] (pc[9]), .\next_pc_for_core[4] (next_pc_for_core[4]), 
           .n12(n12), .data_ready_r_N_2823(data_ready_r_N_2823), .data_ready_r(data_ready_r), 
           .n32706(n32706), .n15569(n15569), .\data_to_write[3] (data_to_write[3]), 
           .\data_to_write[1] (data_to_write[1]), .n2211(n2211), .n17165(n17165), 
           .VCC_net(VCC_net), .n32694(n32694), .n7(n7), .n8854(n8854), 
           .\next_pc_for_core[10] (next_pc_for_core[10]), .\next_pc_for_core[14] (next_pc_for_core[14]), 
           .\instr_data[0][0] (\instr_data[0] [0]), .\instr_data[1][7] (\instr_data[1] [7]), 
           .\instr_data[1][0] (\instr_data[1] [0]), .\instr_data[2][7] (\instr_data[2] [7]), 
           .\next_pc_for_core[8] (next_pc_for_core[8]), .\next_pc_for_core[12] (next_pc_for_core[12]), 
           .\instr_data[2][0] (\instr_data[2] [0]), .\instr_data[3][7] (\instr_data[3] [7]), 
           .n32552(n32552), .n8109(n8109), .n32695(n32695), .n32728(n32728), 
           .n32745(n32745), .\next_pc_for_core[3] (next_pc_for_core[3]), 
           .\next_pc_for_core[5] (next_pc_for_core[5]), .\next_pc_for_core[7] (next_pc_for_core[7]), 
           .\next_pc_for_core[11] (next_pc_for_core[11]), .\pc[21] (pc[21]), 
           .\pc[17] (pc[17]), .\next_pc_for_core[20] (next_pc_for_core[20]), 
           .\next_pc_for_core[16] (next_pc_for_core[16]), .\pc[23] (pc[23]), 
           .\pc[19] (pc[19]), .\pc[22] (pc[22]), .\pc[18] (pc[18]), .\pc[20] (pc[20]), 
           .\pc[16] (pc[16]), .\next_pc_for_core[15] (next_pc_for_core[15]), 
           .\next_pc_for_core[21] (next_pc_for_core[21]), .\next_pc_for_core[17] (next_pc_for_core[17]), 
           .\imm[23] (imm[23]), .\imm[22] (imm[22]), .\imm[19] (imm[19]), 
           .\imm[18] (imm[18]), .\next_pc_for_core[22] (next_pc_for_core[22]), 
           .\next_pc_for_core[18] (next_pc_for_core[18]), .\next_pc_for_core[19] (next_pc_for_core[19]), 
           .n28077(n28077), .\next_pc_for_core[23] (next_pc_for_core[23]), 
           .n32819(n32819), .n32720(n32720), .n29357(n29357), .\uo_out_from_user_peri[1][6] (\uo_out_from_user_peri[1] [6]), 
           .\data_from_user_peri_1__31__N_2455[2] (data_from_user_peri_1__31__N_2455[2]), 
           .\uo_out_from_user_peri[1][2] (\uo_out_from_user_peri[1] [2]), 
           .\uo_out_from_user_peri[1][5] (\uo_out_from_user_peri[1] [5]), 
           .n29491(n29491), .\data_from_read[2] (data_from_read[2]), .\early_branch_addr[7] (early_branch_addr[7]), 
           .\early_branch_addr[3] (early_branch_addr[3]), .\early_branch_addr[6] (early_branch_addr[6]), 
           .\early_branch_addr[2] (early_branch_addr[2]), .\early_branch_addr[4] (early_branch_addr[4]), 
           .n32822(n32822), .\early_branch_addr[8] (early_branch_addr[8]), 
           .\early_branch_addr[5] (early_branch_addr[5]), .\early_branch_addr[9] (early_branch_addr[9]), 
           .\early_branch_addr[10] (early_branch_addr[10]), .\early_branch_addr[11] (early_branch_addr[11]), 
           .\early_branch_addr[12] (early_branch_addr[12]), .\early_branch_addr[13] (early_branch_addr[13]), 
           .\early_branch_addr[14] (early_branch_addr[14]), .\early_branch_addr[15] (early_branch_addr[15]), 
           .\early_branch_addr[17] (early_branch_addr[17]), .\early_branch_addr[18] (early_branch_addr[18]), 
           .\early_branch_addr[19] (early_branch_addr[19]), .\early_branch_addr[20] (early_branch_addr[20]), 
           .\early_branch_addr[21] (early_branch_addr[21]), .\early_branch_addr[22] (early_branch_addr[22]), 
           .\early_branch_addr[23] (early_branch_addr[23]), .\early_branch_addr[16] (early_branch_addr[16]), 
           .n16811(n16811), .n2594(n2594), .n31883(n31883), .\pc_23__N_911[13] (pc_23__N_911[13]), 
           .\pc[12] (pc[12]), .n26838(n26838), .n10944(n10944), .n32725(n32725), 
           .n32761(n32761), .n32729(n32729), .\cycle[0] (cycle[0]), .\pc[8] (pc[8]), 
           .n27178(n27178), .n32766(n32766), .\pc[4] (pc[4]), .n32737(n32737), 
           .\data_from_peri_31__N_2415[0] (data_from_peri_31__N_2415[0]), 
           .n32693(n32693), .clk_c_enable_50(clk_c_enable_50), .n32818(n32818), 
           .clk_c_enable_154(clk_c_enable_154), .clk_c_enable_283(clk_c_enable_283), 
           .clk_c_enable_354(clk_c_enable_354), .\gpio_out_func_sel[0][2] (\gpio_out_func_sel[0] [2]), 
           .\gpio_out_func_sel[1][2] (\gpio_out_func_sel[1] [2]), .\gpio_out_func_sel[2][2] (\gpio_out_func_sel[2] [2]), 
           .\gpio_out_func_sel[3][2] (\gpio_out_func_sel[3] [2]), .n32756(n32756), 
           .n5169(n5169), .n32825(n32825), .n29127(n29127), .\gpio_out_func_sel[4][2] (\gpio_out_func_sel[4] [2]), 
           .\gpio_out_func_sel[6][2] (\gpio_out_func_sel[6] [2]), .\uart_rx_buf_data[4] (uart_rx_buf_data[4]), 
           .\baud_divider[4] (baud_divider_adj_3410[4]), .gpio_out_sel({gpio_out_sel}), 
           .n14(n14), .n14_adj_19(n14_adj_3351), .n29293(n29293), .instr_complete_N_1647(instr_complete_N_1647), 
           .\data_from_read[6] (data_from_read[6]), .n32672(n32672), .n46(n46), 
           .\connect_peripheral[1] (connect_peripheral[1]), .\connect_peripheral[0] (connect_peripheral[0]), 
           .n32568(n32568), .n29741(n29741), .n29(n29), .\uart_rx_buf_data[7] (uart_rx_buf_data[7]), 
           .\baud_divider[7] (baud_divider_adj_3410[7]), .n2(n2_adj_3304), 
           .n32614(n32614), .\next_fsm_state_3__N_3046[3] (next_fsm_state_3__N_3046[3]), 
           .\ui_in_sync[5] (ui_in_sync[5]), .\ui_in_sync[6] (ui_in_sync[6]), 
           .n32072(n32072), .n29549(n29549), .\ui_in_sync[7] (ui_in_sync[7]), 
           .\data_from_user_peri_1__31__N_2455[7] (data_from_user_peri_1__31__N_2455[7]), 
           .\uart_rx_buf_data[6] (uart_rx_buf_data[6]), .n26856(n26856), 
           .\baud_divider[6] (baud_divider_adj_3410[6]), .\uart_rx_buf_data[5] (uart_rx_buf_data[5]), 
           .\baud_divider[5] (baud_divider_adj_3410[5]), .\data_from_read[4] (data_from_read[4]), 
           .\data_from_read[8] (data_from_read[8]), .\data_from_read[12] (data_from_read[12]), 
           .\data_from_read[1] (data_from_read[1]), .\data_from_user_peri_1__31__N_2455[0] (data_from_user_peri_1__31__N_2455[0]), 
           .\uo_out_from_user_peri[1][0] (\uo_out_from_user_peri[1] [0]), 
           .\data_from_read[5] (data_from_read[5]), .data_out_hold(data_out_hold), 
           .\data_from_read[3] (data_from_read[3]), .\data_from_read[7] (data_from_read[7]), 
           .\uart_rx_buf_data[3] (uart_rx_buf_data[3]), .\baud_divider[3] (baud_divider_adj_3410[3]), 
           .n2_adj_20(n2), .\data_from_read[0] (data_from_read[0]), .n32759(n32759), 
           .\uart_rx_buf_data[2] (uart_rx_buf_data[2]), .\baud_divider[2] (baud_divider_adj_3410[2]), 
           .n10737(n10737), .n32650(n32650), .\instr[16] (instr[16]), 
           .n32615(n32615), .n32610(n32610), .clk_c_enable_342(clk_c_enable_342), 
           .\ui_in_sync[1] (ui_in_sync[1]), .\ui_in_sync[0] (ui_in_sync[0]), 
           .debug_rd({debug_rd}), .n29866(n29866), .n17920(n17920), .accum({accum}), 
           .d_3__N_1868({d_3__N_1868}), .fsm_state_adj_24({fsm_state_adj_3483}), 
           .n32791(n32791), .n32763(n32763), .n32730(n32730), .n32834(n32834), 
           .n32710(n32710), .n31351(n31351), .n1152(n1152), .\mul_out[3] (mul_out[3]), 
           .\mul_out[2] (mul_out[2]), .\mul_out[1] (mul_out[1]), .\csr_read_3__N_1447[2] (csr_read_3__N_1447[2]), 
           .\next_accum[5] (next_accum[5]), .GND_net(GND_net), .\next_accum[16] (next_accum[16]), 
           .\next_accum[17] (next_accum[17]), .\next_accum[18] (next_accum[18]), 
           .\next_accum[19] (next_accum[19]), .\next_accum[6] (next_accum[6]), 
           .\next_accum[7] (next_accum[7]), .\next_accum[8] (next_accum[8]), 
           .\next_accum[9] (next_accum[9]), .\next_accum[10] (next_accum[10]), 
           .\next_accum[11] (next_accum[11]), .\next_accum[12] (next_accum[12]), 
           .\next_accum[13] (next_accum[13]), .\next_accum[14] (next_accum[14]), 
           .\next_accum[15] (next_accum[15]), .\next_accum[4] (next_accum[4]), 
           .\return_addr[16] (return_addr[16])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(111[12] 150[6])
    FD1S3AX ui_in_sync_i4 (.D(ui_in_sync0[4]), .CK(clk_c), .Q(ui_in_sync[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i4.GSR = "DISABLED";
    FD1S3AX ui_in_sync0_i2 (.D(ui_in_c_2), .CK(clk_c), .Q(ui_in_sync0[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i2.GSR = "DISABLED";
    FD1P3AX debug_register_data_58 (.D(n8880), .SP(clk_c_enable_286), .CK(clk_c), 
            .Q(debug_register_data));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(250[12] 255[8])
    defparam debug_register_data_58.GSR = "DISABLED";
    FD1S3AX ui_in_sync_i3 (.D(ui_in_sync0[3]), .CK(clk_c), .Q(ui_in_sync[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i3.GSR = "DISABLED";
    CCU2C _add_1_5101_add_4_11 (.A0(cycle_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24218), .COUT(n24219), .S0(n39_adj_3307), 
          .S1(n36));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5101_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_5101_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_5101_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5101_add_4_11.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync0_i1 (.D(ui_in_c_1), .CK(clk_c), .Q(ui_in_sync0[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i1.GSR = "DISABLED";
    FD1S3AX ui_in_sync_i2 (.D(ui_in_sync0[2]), .CK(clk_c), .Q(ui_in_sync[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i2.GSR = "DISABLED";
    CCU2C _add_1_5095_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24316), .S0(next_bit_adj_3349));
    defparam _add_1_5095_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_5095_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_5095_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_5095_add_4_cout.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync0_i0 (.D(ui_in_c_0), .CK(clk_c), .Q(ui_in_sync0[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i0.GSR = "DISABLED";
    IB ui_in_pad_0 (.I(ui_in[0]), .O(ui_in_c_0));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_1 (.I(ui_in[1]), .O(ui_in_c_1));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_2 (.I(ui_in[2]), .O(ui_in_c_2));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_3 (.I(ui_in[3]), .O(ui_in_c_3));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_4 (.I(ui_in[4]), .O(ui_in_c_4));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_5 (.I(ui_in[5]), .O(ui_in_c_5));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_6 (.I(ui_in[6]), .O(ui_in_c_6));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_7 (.I(ui_in[7]), .O(ui_in_c_7));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB rst_n_pad (.I(rst_n), .O(rst_n_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(10[20:25])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    OB uo_out_pad_0 (.I(uo_out_c_0), .O(uo_out[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_1 (.I(uo_out_c_1), .O(uo_out[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    FD1S3AX ui_in_sync_i1 (.D(ui_in_sync0[1]), .CK(clk_c), .Q(ui_in_sync[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i1.GSR = "DISABLED";
    OB uo_out_pad_7 (.I(uo_out_c_7), .O(uo_out[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    LUT4 i28444_3_lut (.A(n32685), .B(n19), .C(n32660), .Z(data_from_read[31])) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i28444_3_lut.init = 16'hcece;
    CCU2C _add_1_5095_add_4_14 (.A0(baud_divider_adj_3410[11]), .B0(cycle_counter_adj_3505[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[12]), 
          .B1(cycle_counter_adj_3505[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24315), .COUT(n24316));
    defparam _add_1_5095_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_5095_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_5095_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_5095_add_4_14.INJECT1_1 = "NO";
    LUT4 i1535_4_lut (.A(pc[2]), .B(n2196), .C(n34285), .D(pc[1]), .Z(n2130)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i1535_4_lut.init = 16'hc5c0;
    LUT4 i24543_4_lut (.A(n32694), .B(n8854), .C(addr[4]), .D(n14), 
         .Z(n27120)) /* synthesis lut_function=(!(A+(B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i24543_4_lut.init = 16'h1511;
    LUT4 i24547_4_lut (.A(n32694), .B(n8854), .C(addr[4]), .D(n14_adj_3351), 
         .Z(n27124)) /* synthesis lut_function=(!(A+(B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i24547_4_lut.init = 16'h1511;
    VLO i1 (.Z(GND_net));
    OB uo_out_pad_2 (.I(uo_out_c_2), .O(uo_out[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    PFUMX i24 (.BLUT(n11), .ALUT(n27757), .C0(\gpio_out_func_sel[0] [1]), 
          .Z(n26466));
    FD1S3AX debug_rd_r_i3 (.D(debug_rd[3]), .CK(clk_c), .Q(debug_rd_r[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(257[12] 259[8])
    defparam debug_rd_r_i3.GSR = "DISABLED";
    FD1S3AX ui_in_sync0_i7 (.D(ui_in_c_7), .CK(clk_c), .Q(ui_in_sync0[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i7.GSR = "DISABLED";
    FD1S3AX debug_rd_r_i2 (.D(debug_rd[2]), .CK(clk_c), .Q(debug_rd_r[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(257[12] 259[8])
    defparam debug_rd_r_i2.GSR = "DISABLED";
    FD1S3AX debug_rd_r_i1 (.D(debug_rd[1]), .CK(clk_c), .Q(debug_rd_r[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(257[12] 259[8])
    defparam debug_rd_r_i1.GSR = "DISABLED";
    CCU2C _add_1_5095_add_4_12 (.A0(baud_divider_adj_3410[9]), .B0(cycle_counter_adj_3505[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[10]), 
          .B1(cycle_counter_adj_3505[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24314), .COUT(n24315));
    defparam _add_1_5095_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_5095_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_5095_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_5095_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_5095_add_4_10 (.A0(baud_divider_adj_3410[7]), .B0(cycle_counter_adj_3505[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[8]), .B1(cycle_counter_adj_3505[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24313), .COUT(n24314));
    defparam _add_1_5095_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_5095_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_5095_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_5095_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_5092_add_4_15 (.A0(addr_adj_3354[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3354[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24259), .S0(addr_24__N_228[13]), .S1(addr_24__N_228[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5092_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_5092_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_5092_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_5092_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_5095_add_4_8 (.A0(baud_divider_adj_3410[5]), .B0(cycle_counter_adj_3505[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[6]), .B1(cycle_counter_adj_3505[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24312), .COUT(n24313));
    defparam _add_1_5095_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_5095_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_5095_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_5095_add_4_8.INJECT1_1 = "NO";
    LUT4 i14152_3_lut (.A(next_pc_for_core[16]), .B(return_addr[16]), .C(n32544), 
         .Z(n16810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(46[23:32])
    defparam i14152_3_lut.init = 16'hcaca;
    LUT4 i14513_3_lut_rep_623 (.A(n2211), .B(n17165), .C(n32734), .Z(n32638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14513_3_lut_rep_623.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut (.A(n2211), .B(n17165), .C(n32734), .D(n32656), 
         .Z(n2594)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h00ca;
    FD1S3IX time_count_3542__i1 (.D(n44), .CK(clk_c), .CD(n765), .Q(time_count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_600_4_lut (.A(n2211), .B(n17165), .C(n32734), .D(n32640), 
         .Z(n32615)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_rep_600_4_lut.init = 16'hffca;
    LUT4 i13753_3_lut (.A(\instr_data[0] [0]), .B(\instr_data[1] [0]), .C(n2130), 
         .Z(n16419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i13753_3_lut.init = 16'hcaca;
    LUT4 i13754_3_lut (.A(\instr_data[2] [0]), .B(\instr_data[3] [0]), .C(n2150), 
         .Z(n16420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i13754_3_lut.init = 16'hcaca;
    CCU2C _add_1_5095_add_4_6 (.A0(baud_divider_adj_3410[3]), .B0(cycle_counter_adj_3505[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[4]), .B1(cycle_counter_adj_3505[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24311), .COUT(n24312));
    defparam _add_1_5095_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_5095_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_5095_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_5095_add_4_6.INJECT1_1 = "NO";
    FD1S3IX time_count_3542__i2 (.D(n43), .CK(clk_c), .CD(n765), .Q(time_count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542__i2.GSR = "DISABLED";
    FD1S3IX time_count_3542__i3 (.D(n42_adj_3335), .CK(clk_c), .CD(n765), 
            .Q(time_count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542__i3.GSR = "DISABLED";
    FD1S3IX time_count_3542__i4 (.D(n41), .CK(clk_c), .CD(n765), .Q(time_count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542__i4.GSR = "DISABLED";
    FD1S3IX time_count_3542__i5 (.D(n40), .CK(clk_c), .CD(n765), .Q(time_count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542__i5.GSR = "DISABLED";
    FD1S3IX time_count_3542__i6 (.D(n39_adj_3333), .CK(clk_c), .CD(n765), 
            .Q(time_count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542__i6.GSR = "DISABLED";
    FD1S3IX time_count_3542__i7 (.D(n38), .CK(clk_c), .CD(n765), .Q(time_count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3542__i7.GSR = "DISABLED";
    CCU2C _add_1_5095_add_4_4 (.A0(baud_divider_adj_3410[1]), .B0(cycle_counter_adj_3505[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[2]), .B1(cycle_counter_adj_3505[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24310), .COUT(n24311));
    defparam _add_1_5095_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_5095_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_5095_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_5095_add_4_4.INJECT1_1 = "NO";
    LUT4 i21743_2_lut_rep_807 (.A(imm[1]), .B(pc[1]), .Z(n32822)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i21743_2_lut_rep_807.init = 16'h6666;
    LUT4 instr_addr_23__I_0_i1_3_lut_4_lut (.A(imm[1]), .B(pc[1]), .C(was_early_branch), 
         .D(instr_addr_23__N_318[0]), .Z(instr_addr[1])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam instr_addr_23__I_0_i1_3_lut_4_lut.init = 16'h6f60;
    CCU2C _add_1_5095_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(baud_divider_adj_3410[0]), .B1(cycle_counter_adj_3505[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n24310));
    defparam _add_1_5095_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_5095_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_5095_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_5095_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_5115_add_4_13 (.A0(cycle_counter_adj_3482[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3482[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n24308), .S0(n33), 
          .S1(n30));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5115_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_5115_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_5115_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5115_add_4_13.INJECT1_1 = "NO";
    LUT4 i3837_4_lut (.A(n32759), .B(n32650), .C(n1152), .D(n32834), 
         .Z(clk_c_enable_342)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B)) */ ;
    defparam i3837_4_lut.init = 16'hccce;
    LUT4 i1_2_lut_rep_810 (.A(addr[3]), .B(addr[4]), .Z(n32825)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_810.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(addr[3]), .B(addr[4]), .C(n32850), .D(addr[27]), 
         .Z(n29263)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_626 (.A(addr_adj_3464[20]), .B(n26811), .C(n4503), 
         .D(fsm_state_adj_3463[0]), .Z(qspi_data_in_3__N_1[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(43[23:51])
    defparam i1_4_lut_adj_626.init = 16'hc088;
    LUT4 i13755_3_lut_rep_639 (.A(n16419), .B(n16420), .C(n32734), .Z(n32654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i13755_3_lut_rep_639.init = 16'hcaca;
    LUT4 \gpio_out_func_sel_0[[4__bdd_3_lut_28904  (.A(\gpio_out_func_sel[2] [4]), 
         .B(addr[2]), .C(\gpio_out_func_sel[3] [4]), .Z(n31791)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam \gpio_out_func_sel_0[[4__bdd_3_lut_28904 .init = 16'he2e2;
    LUT4 i21_1_lut_rep_595_3_lut (.A(n16419), .B(n16420), .C(n32734), 
         .Z(n32610)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam i21_1_lut_rep_595_3_lut.init = 16'h3535;
    LUT4 i2_2_lut_rep_599_4_lut (.A(n16419), .B(n16420), .C(n32734), .D(n32655), 
         .Z(n32614)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;
    defparam i2_2_lut_rep_599_4_lut.init = 16'h3500;
    CCU2C _add_1_5115_add_4_11 (.A0(cycle_counter_adj_3482[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3482[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n24307), .COUT(n24308), 
          .S0(n39), .S1(n36_adj_3314));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5115_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_5115_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_5115_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5115_add_4_11.INJECT1_1 = "NO";
    LUT4 qspi_data_out_3__I_0_i2_3_lut (.A(n4513), .B(qspi_data_oe[1]), 
         .C(n32833), .Z(qspi_data_in_3__N_1[1])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(43[23:51])
    defparam qspi_data_out_3__I_0_i2_3_lut.init = 16'h8c8c;
    CCU2C _add_1_5115_add_4_9 (.A0(cycle_counter_adj_3482[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3482[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n24306), .COUT(n24307), 
          .S0(n45_adj_3312), .S1(n42_adj_3317));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5115_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_5115_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_5115_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5115_add_4_9.INJECT1_1 = "NO";
    LUT4 n29831_bdd_3_lut_29039 (.A(\gpio_out_func_sel[4] [4]), .B(addr[3]), 
         .C(\gpio_out_func_sel[6] [4]), .Z(n31789)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n29831_bdd_3_lut_29039.init = 16'he2e2;
    LUT4 i1_4_lut_adj_627 (.A(addr_adj_3464[22]), .B(n26811), .C(n4501), 
         .D(fsm_state_adj_3463[0]), .Z(qspi_data_in_3__N_1[2])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(43[23:51])
    defparam i1_4_lut_adj_627.init = 16'hc088;
    CCU2C _add_1_5115_add_4_7 (.A0(cycle_counter_adj_3482[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3482[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n24305), .COUT(n24306), 
          .S0(n51_adj_3311), .S1(n48));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5115_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_5115_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_5115_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5115_add_4_7.INJECT1_1 = "NO";
    LUT4 \gpio_out_func_sel_0[[4__bdd_3_lut_29040  (.A(\gpio_out_func_sel[0] [4]), 
         .B(addr[2]), .C(\gpio_out_func_sel[1] [4]), .Z(n31792)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam \gpio_out_func_sel_0[[4__bdd_3_lut_29040 .init = 16'he2e2;
    LUT4 qspi_data_out_3__I_0_i4_3_lut (.A(n32060), .B(qspi_data_oe[1]), 
         .C(n32833), .Z(qspi_data_in_3__N_1[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(43[23:51])
    defparam qspi_data_out_3__I_0_i4_3_lut.init = 16'h8c8c;
    LUT4 i2_3_lut (.A(\gpio_out_func_sel[0] [2]), .B(\gpio_out_func_sel[0] [3]), 
         .C(n26466), .Z(uo_out_c_0)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_3_lut.init = 16'h1010;
    CCU2C _add_1_5115_add_4_5 (.A0(cycle_counter_adj_3482[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3482[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n24304), .COUT(n24305), 
          .S0(n57_adj_3306), .S1(n54_adj_3310));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5115_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_5115_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_5115_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5115_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_5092_add_4_13 (.A0(addr_adj_3354[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3354[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24258), .COUT(n24259), .S0(addr_24__N_228[11]), 
          .S1(addr_24__N_228[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5092_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_5092_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_5092_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5092_add_4_13.INJECT1_1 = "NO";
    FD1P3AX gpio_out_sel_i6 (.D(gpio_out_sel_7__N_13[0]), .SP(clk_c_enable_519), 
            .CK(clk_c), .Q(gpio_out_sel[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(204[12] 211[8])
    defparam gpio_out_sel_i6.GSR = "DISABLED";
    LUT4 i3842_4_lut (.A(n28111), .B(n32524), .C(n6218), .D(n32521), 
         .Z(clk_c_enable_340)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C))) */ ;
    defparam i3842_4_lut.init = 16'hfcdc;
    CCU2C _add_1_5115_add_4_3 (.A0(cycle_counter_adj_3482[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3482[2]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n24303), .COUT(n24304), 
          .S0(n63_adj_3334), .S1(n60_adj_3350));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5115_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_5115_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_5115_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5115_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5115_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycle_counter_adj_3482[0]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .COUT(n24303), .S1(n66));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5115_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5115_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_5115_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5115_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_5092_add_4_11 (.A0(addr_adj_3354[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3354[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24257), .COUT(n24258), .S0(addr_24__N_228[9]), 
          .S1(addr_24__N_228[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5092_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_5092_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_5092_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5092_add_4_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(addr[2]), .B(addr[5]), .Z(n29127)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    CCU2C _add_1_5107_add_4_24 (.A0(imm[23]), .B0(pc[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24302), .S0(early_branch_addr[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_24.INIT1 = 16'h0000;
    defparam _add_1_5107_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_22 (.A0(imm[21]), .B0(pc[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[22]), .B1(pc[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24301), .COUT(n24302), .S0(early_branch_addr[21]), .S1(early_branch_addr[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_20 (.A0(imm[19]), .B0(pc[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[20]), .B1(pc[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24300), .COUT(n24301), .S0(early_branch_addr[19]), .S1(early_branch_addr[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_18 (.A0(imm[17]), .B0(pc[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[18]), .B1(pc[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24299), .COUT(n24300), .S0(early_branch_addr[17]), .S1(early_branch_addr[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_16 (.A0(imm[15]), .B0(pc[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[16]), .B1(pc[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24298), .COUT(n24299), .S0(early_branch_addr[15]), .S1(early_branch_addr[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_5092_add_4_9 (.A0(addr_adj_3354[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3354[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24256), .COUT(n24257), .S0(addr_24__N_228[7]), 
          .S1(addr_24__N_228[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5092_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_5092_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_5092_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5092_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_14 (.A0(imm[13]), .B0(pc[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[14]), .B1(pc[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24297), .COUT(n24298), .S0(early_branch_addr[13]), .S1(early_branch_addr[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_5092_add_4_7 (.A0(addr_adj_3354[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3354[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24255), .COUT(n24256), .S0(addr_24__N_228[5]), 
          .S1(addr_24__N_228[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5092_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_5092_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_5092_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5092_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_5092_add_4_5 (.A0(addr_adj_3354[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3354[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24254), .COUT(n24255), .S0(addr_24__N_228[3]), 
          .S1(addr_24__N_228[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5092_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_5092_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_5092_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5092_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_12 (.A0(imm[11]), .B0(pc[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[12]), .B1(pc[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24296), .COUT(n24297), .S0(early_branch_addr[11]), .S1(early_branch_addr[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_5092_add_4_3 (.A0(addr_adj_3354[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3354[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24253), .COUT(n24254), .S0(addr_24__N_228[1]), 
          .S1(addr_24__N_228[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5092_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_5092_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_5092_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5092_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_10 (.A0(imm[9]), .B0(pc[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[10]), .B1(pc[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24295), .COUT(n24296), .S0(early_branch_addr[9]), .S1(early_branch_addr[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_10.INJECT1_1 = "NO";
    LUT4 i3851_4_lut (.A(n32892), .B(n32524), .C(n32522), .D(n32755), 
         .Z(clk_c_enable_341)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;
    defparam i3851_4_lut.init = 16'heefc;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i3848_4_lut (.A(n32874), .B(n32524), .C(n6220), .D(n1072), 
         .Z(clk_c_enable_66)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C))) */ ;
    defparam i3848_4_lut.init = 16'hfcdc;
    L6MUX21 i28907 (.D0(n31793), .D1(n31790), .SD(addr[4]), .Z(n31794));
    CCU2C _add_1_5107_add_4_8 (.A0(imm[7]), .B0(pc[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[8]), .B1(pc[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24294), .COUT(n24295), .S0(early_branch_addr[7]), .S1(early_branch_addr[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_8.INJECT1_1 = "NO";
    PFUMX i28905 (.BLUT(n31792), .ALUT(n31791), .C0(addr[3]), .Z(n31793));
    CCU2C _add_1_5092_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr_adj_3354[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n24253), .S1(addr_24__N_228[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5092_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5092_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_5092_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5092_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_5098_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24252), .S0(next_bit_adj_3332));
    defparam _add_1_5098_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_5098_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_5098_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_5098_add_4_cout.INJECT1_1 = "NO";
    PFUMX i28902 (.BLUT(n31789), .ALUT(n29831), .C0(addr[2]), .Z(n31790));
    CCU2C _add_1_5107_add_4_6 (.A0(imm[5]), .B0(pc[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[6]), .B1(pc[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24293), .COUT(n24294), .S0(early_branch_addr[5]), .S1(early_branch_addr[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_4 (.A0(imm[3]), .B0(pc[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[4]), .B1(pc[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24292), .COUT(n24293), .S0(early_branch_addr[3]), .S1(early_branch_addr[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_5107_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_4.INJECT1_1 = "NO";
    LUT4 i27175_4_lut (.A(is_writing), .B(is_writing_N_2331), .C(n32523), 
         .D(n8177), .Z(n29884)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i27175_4_lut.init = 16'hcaaa;
    FD1S3AX ui_in_sync_i0 (.D(ui_in_sync0[0]), .CK(clk_c), .Q(ui_in_sync[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i0.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_628 (.A(n29631), .B(n29337), .C(n29333), .D(n29335), 
         .Z(n10737)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_628.init = 16'hfffd;
    LUT4 i26988_2_lut (.A(time_count[3]), .B(time_count[4]), .Z(n29631)) /* synthesis lut_function=(A (B)) */ ;
    defparam i26988_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_629 (.A(time_count[1]), .B(time_count[5]), .Z(n29337)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_629.init = 16'heeee;
    LUT4 i1_2_lut_adj_630 (.A(time_count[2]), .B(time_count[0]), .Z(n29333)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_630.init = 16'heeee;
    LUT4 i1_2_lut_adj_631 (.A(time_count[7]), .B(time_count[6]), .Z(n29335)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_631.init = 16'heeee;
    CCU2C _add_1_5107_add_4_2 (.A0(imm[1]), .B0(pc[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[2]), .B1(pc[2]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n24292), .S1(early_branch_addr[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5107_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_5107_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_5107_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_23 (.A0(early_branch_addr[23]), .B0(was_early_branch), 
          .C0(pc[23]), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24290), .S0(instr_addr_23__N_318[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_23.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_23.INIT1 = 16'h0000;
    defparam _add_1_5110_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_5098_add_4_14 (.A0(baud_divider_adj_3410[11]), .B0(cycle_counter_adj_3482[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[12]), 
          .B1(cycle_counter_adj_3482[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24251), .COUT(n24252));
    defparam _add_1_5098_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_5098_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_5098_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_5098_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_5098_add_4_12 (.A0(baud_divider_adj_3410[9]), .B0(cycle_counter_adj_3482[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[10]), 
          .B1(cycle_counter_adj_3482[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n24250), .COUT(n24251));
    defparam _add_1_5098_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_5098_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_5098_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_5098_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_5098_add_4_10 (.A0(baud_divider_adj_3410[7]), .B0(cycle_counter_adj_3482[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[8]), .B1(cycle_counter_adj_3482[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24249), .COUT(n24250));
    defparam _add_1_5098_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_5098_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_5098_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_5098_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_5098_add_4_8 (.A0(baud_divider_adj_3410[5]), .B0(cycle_counter_adj_3482[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[6]), .B1(cycle_counter_adj_3482[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24248), .COUT(n24249));
    defparam _add_1_5098_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_5098_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_5098_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_5098_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_5098_add_4_6 (.A0(baud_divider_adj_3410[3]), .B0(cycle_counter_adj_3482[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3410[4]), .B1(cycle_counter_adj_3482[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24247), .COUT(n24248));
    defparam _add_1_5098_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_5098_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_5098_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_5098_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_21 (.A0(early_branch_addr[21]), .B0(was_early_branch), 
          .C0(pc[21]), .D0(VCC_net), .A1(early_branch_addr[22]), .B1(was_early_branch), 
          .C1(pc[22]), .D1(VCC_net), .CIN(n24289), .COUT(n24290), .S0(instr_addr_23__N_318[20]), 
          .S1(instr_addr_23__N_318[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_21.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_21.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_19 (.A0(early_branch_addr[19]), .B0(was_early_branch), 
          .C0(pc[19]), .D0(VCC_net), .A1(early_branch_addr[20]), .B1(was_early_branch), 
          .C1(pc[20]), .D1(VCC_net), .CIN(n24288), .COUT(n24289), .S0(instr_addr_23__N_318[18]), 
          .S1(instr_addr_23__N_318[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_19.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_19.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_17 (.A0(early_branch_addr[17]), .B0(was_early_branch), 
          .C0(pc[17]), .D0(VCC_net), .A1(early_branch_addr[18]), .B1(was_early_branch), 
          .C1(pc[18]), .D1(VCC_net), .CIN(n24287), .COUT(n24288), .S0(instr_addr_23__N_318[16]), 
          .S1(instr_addr_23__N_318[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_17.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_17.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_15 (.A0(early_branch_addr[15]), .B0(was_early_branch), 
          .C0(pc[15]), .D0(VCC_net), .A1(early_branch_addr[16]), .B1(was_early_branch), 
          .C1(pc[16]), .D1(VCC_net), .CIN(n24286), .COUT(n24287), .S0(instr_addr_23__N_318[14]), 
          .S1(instr_addr_23__N_318[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_15.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_15.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_5101_add_4_9 (.A0(cycle_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24217), .COUT(n24218), .S0(n45), .S1(n42));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5101_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_5101_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_5101_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5101_add_4_9.INJECT1_1 = "NO";
    LUT4 i27178_3_lut (.A(data_stall), .B(data_stall_N_2158), .C(continue_txn_N_2131), 
         .Z(n29887)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam i27178_3_lut.init = 16'hcece;
    CCU2C _add_1_5110_add_4_13 (.A0(early_branch_addr[13]), .B0(was_early_branch), 
          .C0(pc[13]), .D0(VCC_net), .A1(early_branch_addr[14]), .B1(was_early_branch), 
          .C1(pc[14]), .D1(VCC_net), .CIN(n24285), .COUT(n24286), .S0(instr_addr_23__N_318[12]), 
          .S1(instr_addr_23__N_318[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_13.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_13.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_13.INJECT1_1 = "NO";
    LUT4 i14837_2_lut (.A(qspi_data_in[0]), .B(rst_reg_n), .Z(qspi_data_out_3__N_5[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(127[22:56])
    defparam i14837_2_lut.init = 16'h8888;
    PFUMX i14154 (.BLUT(n16810), .ALUT(n16811), .C0(n32552), .Z(pc_23__N_911[13]));
    LUT4 i6176_2_lut (.A(addr[3]), .B(addr[2]), .Z(n8854)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6176_2_lut.init = 16'h8888;
    CCU2C _add_1_5110_add_4_11 (.A0(early_branch_addr[11]), .B0(was_early_branch), 
          .C0(pc[11]), .D0(VCC_net), .A1(early_branch_addr[12]), .B1(was_early_branch), 
          .C1(pc[12]), .D1(VCC_net), .CIN(n24284), .COUT(n24285), .S0(instr_addr_23__N_318[10]), 
          .S1(instr_addr_23__N_318[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_11.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_11.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_11.INJECT1_1 = "NO";
    LUT4 mux_34_i2_3_lut (.A(ui_in_c_0), .B(data_to_write[7]), .C(n762), 
         .Z(gpio_out_sel_7__N_13[1])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(209[13:93])
    defparam mux_34_i2_3_lut.init = 16'hc5c5;
    LUT4 i28416_2_lut (.A(n10737), .B(rst_reg_n), .Z(n765)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i28416_2_lut.init = 16'h7777;
    CCU2C _add_1_5110_add_4_9 (.A0(early_branch_addr[9]), .B0(was_early_branch), 
          .C0(pc[9]), .D0(VCC_net), .A1(early_branch_addr[10]), .B1(was_early_branch), 
          .C1(pc[10]), .D1(VCC_net), .CIN(n24283), .COUT(n24284), .S0(instr_addr_23__N_318[8]), 
          .S1(instr_addr_23__N_318[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5110_add_4_9.INIT0 = 16'hb8b8;
    defparam _add_1_5110_add_4_9.INIT1 = 16'hb8b8;
    defparam _add_1_5110_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_9.INJECT1_1 = "NO";
    LUT4 i25_4_lut (.A(\uo_out_from_user_peri[1] [0]), .B(led_state), .C(\gpio_out_func_sel[0] [4]), 
         .D(\gpio_out_func_sel[0] [0]), .Z(n11)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    defparam i25_4_lut.init = 16'h0a30;
    LUT4 i1_4_lut_adj_632 (.A(n32685), .B(n32672), .C(n32745), .D(n29263), 
         .Z(debug_uart_tx_start)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_632.init = 16'h0100;
    LUT4 i1_4_lut_adj_633 (.A(connect_peripheral[0]), .B(n46), .C(connect_peripheral[1]), 
         .D(n29293), .Z(n762)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_633.init = 16'h2000;
    LUT4 instr_1__bdd_3_lut (.A(n32548), .B(n32642), .C(rd[0]), .Z(n32072)) /* synthesis lut_function=(!(A (C)+!A !(B))) */ ;
    defparam instr_1__bdd_3_lut.init = 16'h4e4e;
    LUT4 peri_out_3__I_0_3_lut (.A(peri_out[3]), .B(debug_rd_r[1]), .C(debug_register_data), 
         .Z(uo_out_c_3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(155[24:73])
    defparam peri_out_3__I_0_3_lut.init = 16'hcaca;
    LUT4 i14512_3_lut (.A(\instr_data[2] [7]), .B(\instr_data[3] [7]), .C(n2150), 
         .Z(n17165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14512_3_lut.init = 16'hcaca;
    LUT4 i14538_rep_88_3_lut (.A(\instr_data[1] [7]), .B(\instr_data[2] [7]), 
         .C(n2130), .Z(n29707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i14538_rep_88_3_lut.init = 16'hcaca;
    LUT4 i15166_2_lut (.A(qspi_data_in[3]), .B(rst_reg_n), .Z(qspi_data_out_3__N_5[3])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(127[22:56])
    defparam i15166_2_lut.init = 16'h8888;
    LUT4 i15169_2_lut (.A(qspi_data_in[2]), .B(rst_reg_n), .Z(qspi_data_out_3__N_5[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(127[22:56])
    defparam i15169_2_lut.init = 16'h8888;
    LUT4 peri_out_4__I_0_3_lut (.A(peri_out[4]), .B(debug_rd_r[2]), .C(debug_register_data), 
         .Z(uo_out_c_4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(156[24:73])
    defparam peri_out_4__I_0_3_lut.init = 16'hcaca;
    LUT4 peri_out_5__I_0_3_lut (.A(peri_out[5]), .B(debug_rd_r[3]), .C(debug_register_data), 
         .Z(uo_out_c_5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(157[24:73])
    defparam peri_out_5__I_0_3_lut.init = 16'hcaca;
    LUT4 debug_uart_txd_I_0_3_lut (.A(debug_uart_txd), .B(peri_out[6]), 
         .C(gpio_out_sel[6]), .Z(uo_out_c_6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(158[24:70])
    defparam debug_uart_txd_I_0_3_lut.init = 16'hcaca;
    LUT4 i6202_3_lut (.A(ui_in_c_1), .B(data_to_write[0]), .C(rst_reg_n), 
         .Z(n8880)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(250[12] 255[8])
    defparam i6202_3_lut.init = 16'hcaca;
    LUT4 i15555_3_lut_rep_685_4_lut (.A(n32771), .B(n32801), .C(n32727), 
         .D(rst_reg_n), .Z(n32700)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;
    defparam i15555_3_lut_rep_685_4_lut.init = 16'hfddd;
    tqvp_uart_tx_U1 i_debug_uart_tx (.debug_uart_txd(debug_uart_txd), .clk_c(clk_c), 
            .clk_c_enable_432(clk_c_enable_432), .cycle_counter({cycle_counter}), 
            .clk_c_enable_143(clk_c_enable_143), .n6142(n6142), .n72({n30_adj_3309, 
            n33_adj_3308, n36, n39_adj_3307, n42, n45, n48_adj_3305, 
            n51, n54, n57, n60, n63, n66_adj_3313}), .\fsm_state[0] (fsm_state[0]), 
            .next_bit(next_bit), .n32756(n32756), .debug_uart_tx_start(debug_uart_tx_start), 
            .\data_to_write[6] (data_to_write[6]), .\data_to_write[0] (data_to_write[0]), 
            .\data_to_write[5] (data_to_write[5]), .\data_to_write[4] (data_to_write[4]), 
            .\data_to_write[3] (data_to_write[3]), .\data_to_write[2] (data_to_write[2]), 
            .\data_to_write[1] (data_to_write[1]), .clk_c_enable_495(clk_c_enable_495), 
            .n32832(n32832), .uart_txd_N_3005(uart_txd_N_3005), .rst_reg_n(rst_reg_n), 
            .\data_to_write[7] (data_to_write[7]), .n26870(n26870), .n32622(n32622)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[4] 236[3])
    LUT4 i27256_2_lut_rep_553_4_lut (.A(pc[2]), .B(n32766), .C(debug_instr_valid), 
         .D(n4251), .Z(n32568)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i27256_2_lut_rep_553_4_lut.init = 16'h0035;
    LUT4 i13752_rep_119_3_lut (.A(n16417), .B(instr[31]), .C(n4251), .Z(n29738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i13752_rep_119_3_lut.init = 16'hcaca;
    LUT4 i13751_3_lut (.A(\instr_data[3] [0]), .B(\instr_data[0] [0]), .C(n2150), 
         .Z(n16417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i13751_3_lut.init = 16'hcaca;
    LUT4 i13752_3_lut (.A(n29741), .B(n16417), .C(n32734), .Z(instr[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i13752_3_lut.init = 16'hcaca;
    sim_qspi_pmod i_qspi (.qspi_data_in({qspi_data_in}), .qspi_clk_N_56(qspi_clk_N_56), 
            .\addr[14] (addr_adj_3354[14]), .\addr_24__N_228[14] (addr_24__N_228[14]), 
            .\addr[13] (addr_adj_3354[13]), .\addr[12] (addr_adj_3354[12]), 
            .\addr[11] (addr_adj_3354[11]), .\addr[10] (addr_adj_3354[10]), 
            .\addr[9] (addr_adj_3354[9]), .GND_net(GND_net), .VCC_net(VCC_net), 
            .\addr[8] (addr_adj_3354[8]), .\addr[7] (addr_adj_3354[7]), 
            .\addr[6] (addr_adj_3354[6]), .\addr[5] (addr_adj_3354[5]), 
            .\addr[4] (addr_adj_3354[4]), .\addr[3] (addr_adj_3354[3]), 
            .\addr[0] (addr_adj_3354[0]), .\addr[2] (addr_adj_3354[2]), 
            .\addr[1] (addr_adj_3354[1]), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), .\writing_N_164[3] (writing_N_164[3]), 
            .qspi_ram_a_select(qspi_ram_a_select), .qspi_ram_b_select(qspi_ram_b_select), 
            .n32802(n32802), .\addr_24__N_228[0] (addr_24__N_228[0]), .\addr_24__N_228[1] (addr_24__N_228[1]), 
            .\addr_24__N_228[11] (addr_24__N_228[11]), .\addr_24__N_228[13] (addr_24__N_228[13]), 
            .\addr_24__N_228[12] (addr_24__N_228[12]), .\addr_24__N_228[2] (addr_24__N_228[2]), 
            .\addr_24__N_228[3] (addr_24__N_228[3]), .\addr_24__N_228[4] (addr_24__N_228[4]), 
            .\addr_24__N_228[5] (addr_24__N_228[5]), .\addr_24__N_228[6] (addr_24__N_228[6]), 
            .\addr_24__N_228[7] (addr_24__N_228[7]), .\addr_24__N_228[8] (addr_24__N_228[8]), 
            .\addr_24__N_228[9] (addr_24__N_228[9]), .\addr_24__N_228[10] (addr_24__N_228[10])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(42[19] 50[6])
    
endmodule
//
// Verilog Description of module \peripherals_min(CLOCK_MHZ=25) 
//

module \peripherals_min(CLOCK_MHZ=25)  (clk_c, clk_c_enable_432, \data_to_write[3] , 
            \peri_data_out[0] , data_out_hold, n32706, \data_to_write[1] , 
            \peri_data_out[1] , n15569, \peri_data_out[2] , n26116, 
            \peri_data_out[3] , \peri_data_out[4] , clk_c_enable_50, \peri_data_out[5] , 
            n3, n32520, \addr[7] , n2, \peri_data_out[6] , n3_adj_47, 
            n28077, \addr[10] , n32851, \addr[6] , n12, \gpio_out_func_sel[0] , 
            \data_to_write[4] , n32835, n32836, \addr[2] , n29, \data_to_write[0] , 
            \peri_data_out[7] , \peri_data_out[8] , baud_divider, \gpio_out_func_sel[6][2] , 
            \data_to_write[2] , \peri_data_out[9] , \gpio_out_func_sel[2][4] , 
            \gpio_out_func_sel[7][4] , clk_c_enable_154, \gpio_out_func_sel[1][4] , 
            \gpio_out_func_sel[1][2] , uo_out_c_1, \gpio_out_func_sel[4] , 
            n2_adj_48, n26856, \gpio_out_func_sel[7][2] , \uo_out_from_user_peri[1] , 
            \peri_data_out[10] , \gpio_out_func_sel[3][4] , \gpio_out_func_sel[3][2] , 
            clk_c_enable_283, \gpio_out_func_sel[2][2] , \peri_data_out[11] , 
            \peri_data_out[12] , \gpio_out_func_sel[5][4] , \gpio_out_func_sel[6][4] , 
            \gpio_out_func_sel[5][2] , \gpio_out_func_sel[4][4] , clk_c_enable_354, 
            data_ready_r, rst_reg_n, data_ready_r_N_2823, \addr[4] , 
            \addr[3] , n32818, n10944, \uo_out_from_user_peri[1][2] , 
            \uo_out_from_user_peri[1][5] , \data_to_write[5] , \uo_out_from_user_peri[1][6] , 
            \data_to_write[6] , \data_to_write[7] , \gpio_out_sel[7] , 
            uo_out_c_7, \ui_in_sync[2] , n31883, n26838, \data_from_user_peri_1__31__N_2455[2] , 
            led_state, \addr[1] , n27888, n32693, n32729, n8854, 
            n32819, \debug_rd_r[0] , debug_register_data, uo_out_c_2, 
            \ui_in_sync[1] , n32761, \ui_in_sync[3] , \ui_in_sync[4] , 
            n31794, \ui_in_sync[0] , \data_from_user_peri_1__31__N_2455[0] , 
            n32723, n32727, n32728, n32720, n32737, \peri_out[3] , 
            \data_from_user_peri_1__31__N_2455[7] , \peri_out[4] , n32801, 
            n8109, n32700, \peri_out[5] , \peri_out[6] , \data_from_peri_31__N_2415[0] , 
            \data_to_write[12] , \data_to_write[11] , \data_to_write[10] , 
            \data_to_write[9] , \data_to_write[8] , \ui_in_sync[7] , n31706, 
            \uart_rx_buf_data[2] , \uart_rx_buf_data[3] , \uart_rx_buf_data[4] , 
            \uart_rx_buf_data[5] , \uart_rx_buf_data[6] , \uart_rx_buf_data[7] , 
            \next_fsm_state_3__N_3046[3] , n31795, n31796, \addr[5] , 
            \addr[0] , n32695, n32730, n26870, n32725, qv_data_write_n, 
            n32710, \imm[6] , \csr_read_3__N_1447[2] , n29866, n29491, 
            cycle_counter, n72, n32791, fsm_state, next_bit, n27757, 
            n32763, n32251, GND_net, VCC_net, cycle_counter_adj_65, 
            next_bit_adj_62, debug_stop_txn, instr_active_N_2106, stop_txn_reg, 
            n32755, stop_txn_now_N_2363, clk_c_enable_208, n32714, qspi_write_done, 
            n10672, spi_clk_pos, n28259, next_bit_adj_63, n32622, 
            uart_txd_N_3005, clk_c_enable_495, n32832, \fsm_state[0]_adj_64 , 
            clk_c_enable_143, n762, clk_c_enable_519, n8177, n32524, 
            n29357, n46, clk_c_enable_286, instr_complete_N_1647, n28957, 
            n32771, n27178, n29549, n6142, n28319, n32681, n27931, 
            n1072, clk_c_enable_543, qv_data_read_n, n26691, \qspi_data_in[1] , 
            \qspi_data_out_3__N_5[1] , n26692) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output clk_c_enable_432;
    input \data_to_write[3] ;
    output \peri_data_out[0] ;
    output data_out_hold;
    input n32706;
    input \data_to_write[1] ;
    output \peri_data_out[1] ;
    input n15569;
    output \peri_data_out[2] ;
    input n26116;
    output \peri_data_out[3] ;
    output \peri_data_out[4] ;
    input clk_c_enable_50;
    output \peri_data_out[5] ;
    input n3;
    input n32520;
    input \addr[7] ;
    input n2;
    output \peri_data_out[6] ;
    input n3_adj_47;
    input n28077;
    input \addr[10] ;
    input n32851;
    input \addr[6] ;
    output n12;
    output [4:0]\gpio_out_func_sel[0] ;
    input \data_to_write[4] ;
    input n32835;
    output n32836;
    input \addr[2] ;
    output n29;
    input \data_to_write[0] ;
    output \peri_data_out[7] ;
    output \peri_data_out[8] ;
    output [12:0]baud_divider;
    output \gpio_out_func_sel[6][2] ;
    input \data_to_write[2] ;
    output \peri_data_out[9] ;
    output \gpio_out_func_sel[2][4] ;
    output \gpio_out_func_sel[7][4] ;
    input clk_c_enable_154;
    output \gpio_out_func_sel[1][4] ;
    output \gpio_out_func_sel[1][2] ;
    output uo_out_c_1;
    output [4:0]\gpio_out_func_sel[4] ;
    input n2_adj_48;
    output n26856;
    output \gpio_out_func_sel[7][2] ;
    output [7:0]\uo_out_from_user_peri[1] ;
    output \peri_data_out[10] ;
    output \gpio_out_func_sel[3][4] ;
    output \gpio_out_func_sel[3][2] ;
    input clk_c_enable_283;
    output \gpio_out_func_sel[2][2] ;
    output \peri_data_out[11] ;
    output \peri_data_out[12] ;
    output \gpio_out_func_sel[5][4] ;
    output \gpio_out_func_sel[6][4] ;
    output \gpio_out_func_sel[5][2] ;
    output \gpio_out_func_sel[4][4] ;
    input clk_c_enable_354;
    output data_ready_r;
    input rst_reg_n;
    input data_ready_r_N_2823;
    input \addr[4] ;
    input \addr[3] ;
    output n32818;
    output n10944;
    output \uo_out_from_user_peri[1][2] ;
    output \uo_out_from_user_peri[1][5] ;
    input \data_to_write[5] ;
    output \uo_out_from_user_peri[1][6] ;
    input \data_to_write[6] ;
    input \data_to_write[7] ;
    input \gpio_out_sel[7] ;
    output uo_out_c_7;
    input \ui_in_sync[2] ;
    input n31883;
    input n26838;
    output \data_from_user_peri_1__31__N_2455[2] ;
    output led_state;
    input \addr[1] ;
    input n27888;
    input n32693;
    input n32729;
    input n8854;
    input n32819;
    input \debug_rd_r[0] ;
    input debug_register_data;
    output uo_out_c_2;
    input \ui_in_sync[1] ;
    input n32761;
    input \ui_in_sync[3] ;
    input \ui_in_sync[4] ;
    input n31794;
    input \ui_in_sync[0] ;
    output \data_from_user_peri_1__31__N_2455[0] ;
    input n32723;
    input n32727;
    input n32728;
    input n32720;
    input n32737;
    output \peri_out[3] ;
    input \data_from_user_peri_1__31__N_2455[7] ;
    output \peri_out[4] ;
    input n32801;
    input n8109;
    input n32700;
    output \peri_out[5] ;
    output \peri_out[6] ;
    input \data_from_peri_31__N_2415[0] ;
    input \data_to_write[12] ;
    input \data_to_write[11] ;
    input \data_to_write[10] ;
    input \data_to_write[9] ;
    input \data_to_write[8] ;
    input \ui_in_sync[7] ;
    output n31706;
    output \uart_rx_buf_data[2] ;
    output \uart_rx_buf_data[3] ;
    output \uart_rx_buf_data[4] ;
    output \uart_rx_buf_data[5] ;
    output \uart_rx_buf_data[6] ;
    output \uart_rx_buf_data[7] ;
    output \next_fsm_state_3__N_3046[3] ;
    output n31795;
    output n31796;
    input \addr[5] ;
    input \addr[0] ;
    input n32695;
    input n32730;
    input n26870;
    input n32725;
    input [1:0]qv_data_write_n;
    input n32710;
    input \imm[6] ;
    input \csr_read_3__N_1447[2] ;
    output n29866;
    input n29491;
    output [12:0]cycle_counter;
    input [12:0]n72;
    input n32791;
    output [3:0]fsm_state;
    input next_bit;
    output n27757;
    input n32763;
    output n32251;
    input GND_net;
    input VCC_net;
    output [12:0]cycle_counter_adj_65;
    input next_bit_adj_62;
    input debug_stop_txn;
    output instr_active_N_2106;
    input stop_txn_reg;
    input n32755;
    input stop_txn_now_N_2363;
    output clk_c_enable_208;
    input n32714;
    input qspi_write_done;
    output n10672;
    input spi_clk_pos;
    output n28259;
    input next_bit_adj_63;
    input n32622;
    input uart_txd_N_3005;
    output clk_c_enable_495;
    input n32832;
    input \fsm_state[0]_adj_64 ;
    output clk_c_enable_143;
    input n762;
    output clk_c_enable_519;
    output n8177;
    output n32524;
    input n29357;
    input n46;
    output clk_c_enable_286;
    input instr_complete_N_1647;
    input n28957;
    input n32771;
    input n27178;
    input n29549;
    output n6142;
    input n28319;
    input n32681;
    output n27931;
    input n1072;
    output clk_c_enable_543;
    input [1:0]qv_data_read_n;
    output n26691;
    input \qspi_data_in[1] ;
    output \qspi_data_out_3__N_5[1] ;
    output n26692;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [4:0]\gpio_out_func_sel[3] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    
    wire clk_c_enable_278, clk_c_enable_324;
    wire [31:0]data_from_peri;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(47[16:30])
    
    wire clk_c_enable_6;
    wire [4:0]\gpio_out_func_sel[6] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    
    wire clk_c_enable_355, n3_c, n3_adj_3261, n3_adj_3262;
    wire [4:0]\gpio_out_func_sel[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    
    wire n8876, n1, n1_adj_3264, n1_adj_3266;
    wire [4:0]\gpio_out_func_sel[5] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    
    wire clk_c_enable_100, clk_c_enable_356, clk_c_enable_359, n3_adj_3267, 
        n11704;
    wire [4:0]\gpio_out_func_sel[7] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    
    wire clk_c_enable_270;
    wire [4:0]\gpio_out_func_sel[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    
    wire n9031, n3_adj_3268, clk_c_enable_353, n1_adj_3269, clk_c_enable_358;
    wire [4:0]\gpio_out_func_sel[4]_c ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(123[15:32])
    
    wire clk_c_enable_463, clk_c_enable_284, clk_c_enable_366, clk_c_enable_368, 
        clk_c_enable_369, n30269, n30270, n30271, n30276, n30277, 
        n30278, n32719, n30283, n30284, n30285, n30282, n30281;
    wire [7:0]\uo_out_from_user_peri[1]_c ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(59[17:38])
    wire [7:0]\uo_out_from_user_peri[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(59[17:38])
    
    wire n30280, n30279, n30275, n30274, n30273, n30272, n30268, 
        n30267, n30266, n30265, n3_adj_3271, n6;
    wire [7:0]data_from_peri_31__N_2447;
    
    wire n28053, n9;
    wire [31:0]data_from_user_peri_1__31__N_2455;
    
    wire n29531, n3_adj_3272, n3_adj_3273, n32757, n32666, n3_adj_3274, 
        n3_adj_3275, clk_c_enable_64, clk_c_enable_282;
    
    FD1P3IX \gpio_out_func_sel_3[[3__367  (.D(\data_to_write[3] ), .SP(clk_c_enable_278), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[3] [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_3[[3__367 .GSR = "DISABLED";
    FD1P3AX data_out_r_i0_i1 (.D(data_from_peri[0]), .SP(clk_c_enable_324), 
            .CK(clk_c), .Q(\peri_data_out[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i1.GSR = "DISABLED";
    FD1P3IX data_out_hold_347 (.D(n32706), .SP(clk_c_enable_6), .CD(clk_c_enable_432), 
            .CK(clk_c), .Q(data_out_hold)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_hold_347.GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_6[[1__384  (.D(\data_to_write[1] ), .SP(clk_c_enable_355), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[6] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_6[[1__384 .GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i2 (.D(n3_c), .SP(clk_c_enable_324), .CD(n15569), 
            .CK(clk_c), .Q(\peri_data_out[1] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i2.GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i3 (.D(n26116), .SP(clk_c_enable_324), .CD(n15569), 
            .CK(clk_c), .Q(\peri_data_out[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i3.GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i4 (.D(n3_adj_3261), .SP(clk_c_enable_324), .CD(n15569), 
            .CK(clk_c), .Q(\peri_data_out[3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i4.GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i5 (.D(n3_adj_3262), .SP(clk_c_enable_324), .CD(n15569), 
            .CK(clk_c), .Q(\peri_data_out[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i5.GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_2[[0__365  (.D(n8876), .SP(clk_c_enable_50), 
            .CK(clk_c), .Q(\gpio_out_func_sel[2] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_2[[0__365 .GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i6 (.D(n3), .SP(clk_c_enable_324), .CD(n15569), 
            .CK(clk_c), .Q(\peri_data_out[5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i6.GSR = "DISABLED";
    PFUMX addr_in_9__I_0_539_Mux_1_i3 (.BLUT(n1), .ALUT(n32520), .C0(\addr[7] ), 
          .Z(n3_c)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    PFUMX addr_in_9__I_0_539_Mux_3_i3 (.BLUT(n1_adj_3264), .ALUT(n2), .C0(\addr[7] ), 
          .Z(n3_adj_3261)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    FD1P3IX data_out_r_i0_i7 (.D(n3_adj_47), .SP(clk_c_enable_324), .CD(n15569), 
            .CK(clk_c), .Q(\peri_data_out[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i7.GSR = "DISABLED";
    PFUMX addr_in_9__I_0_539_Mux_4_i3 (.BLUT(n1_adj_3266), .ALUT(n28077), 
          .C0(\addr[7] ), .Z(n3_adj_3262)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    LUT4 i1_4_lut (.A(\addr[10] ), .B(\addr[7] ), .C(n32851), .D(\addr[6] ), 
         .Z(n12)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_4_lut.init = 16'hfaea;
    FD1P3AX \gpio_out_func_sel_5[[0__380  (.D(n8876), .SP(clk_c_enable_100), 
            .CK(clk_c), .Q(\gpio_out_func_sel[5] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_5[[0__380 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_0[[4__351  (.D(\data_to_write[4] ), .SP(clk_c_enable_356), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[0] [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_0[[4__351 .GSR = "DISABLED";
    LUT4 i28557_2_lut_4_lut (.A(n32835), .B(n32836), .C(\addr[2] ), .D(\addr[6] ), 
         .Z(n29)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i28557_2_lut_4_lut.init = 16'h0001;
    FD1P3IX \gpio_out_func_sel_0[[0__355  (.D(\data_to_write[0] ), .SP(clk_c_enable_356), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[0] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_0[[0__355 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_2[[3__362  (.D(\data_to_write[3] ), .SP(clk_c_enable_359), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[2] [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_2[[3__362 .GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i8 (.D(n3_adj_3267), .SP(clk_c_enable_324), .CD(n15569), 
            .CK(clk_c), .Q(\peri_data_out[7] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i8.GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i9 (.D(baud_divider[8]), .SP(clk_c_enable_324), 
            .CD(n11704), .CK(clk_c), .Q(\peri_data_out[8] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i9.GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_6[[2__383  (.D(\data_to_write[2] ), .SP(clk_c_enable_355), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[6][2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_6[[2__383 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_3[[1__369  (.D(\data_to_write[1] ), .SP(clk_c_enable_278), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[3] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_3[[1__369 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_7[[1__389  (.D(\data_to_write[1] ), .SP(clk_c_enable_270), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[7] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_7[[1__389 .GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i10 (.D(baud_divider[9]), .SP(clk_c_enable_324), 
            .CD(n11704), .CK(clk_c), .Q(\peri_data_out[9] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i10.GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_2[[4__361  (.D(\data_to_write[4] ), .SP(clk_c_enable_359), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[2][4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_2[[4__361 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_7[[4__386  (.D(\data_to_write[4] ), .SP(clk_c_enable_270), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[7][4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_7[[4__386 .GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_1[[1__359  (.D(n9031), .SP(clk_c_enable_154), 
            .CK(clk_c), .Q(\gpio_out_func_sel[1] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_1[[1__359 .GSR = "DISABLED";
    LUT4 i28547_4_lut (.A(\gpio_out_func_sel[1] [3]), .B(n3_adj_3268), .C(\gpio_out_func_sel[1][4] ), 
         .D(\gpio_out_func_sel[1][2] ), .Z(uo_out_c_1)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam i28547_4_lut.init = 16'h0004;
    FD1P3IX \gpio_out_func_sel_4[[2__373  (.D(\data_to_write[2] ), .SP(clk_c_enable_353), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[4] [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_4[[2__373 .GSR = "DISABLED";
    PFUMX addr_in_9__I_0_539_Mux_7_i3 (.BLUT(n1_adj_3269), .ALUT(n2_adj_48), 
          .C0(\addr[7] ), .Z(n3_adj_3267)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    FD1P3IX \gpio_out_func_sel_1[[4__356  (.D(\data_to_write[4] ), .SP(clk_c_enable_358), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[1][4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_1[[4__356 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_7[[3__387  (.D(\data_to_write[3] ), .SP(clk_c_enable_270), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[7] [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_7[[3__387 .GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(n32835), .B(n32836), .C(\addr[2] ), .D(\addr[7] ), 
         .Z(n26856)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0100;
    FD1P3IX \gpio_out_func_sel_4[[3__372  (.D(\data_to_write[3] ), .SP(clk_c_enable_353), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[4]_c [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_4[[3__372 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_7[[2__388  (.D(\data_to_write[2] ), .SP(clk_c_enable_270), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[7][2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_7[[2__388 .GSR = "DISABLED";
    FD1P3IX gpio_out__i0 (.D(\data_to_write[0] ), .SP(clk_c_enable_463), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\uo_out_from_user_peri[1] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(126[12] 134[8])
    defparam gpio_out__i0.GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i11 (.D(baud_divider[10]), .SP(clk_c_enable_324), 
            .CD(n11704), .CK(clk_c), .Q(\peri_data_out[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i11.GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_3[[4__366  (.D(\data_to_write[4] ), .SP(clk_c_enable_278), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[3][4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_3[[4__366 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_3[[2__368  (.D(\data_to_write[2] ), .SP(clk_c_enable_278), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[3][2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_3[[2__368 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_4[[1__374  (.D(\data_to_write[1] ), .SP(clk_c_enable_353), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[4]_c [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_4[[1__374 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_0[[3__352  (.D(\data_to_write[3] ), .SP(clk_c_enable_356), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[0] [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_0[[3__352 .GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_0[[1__354  (.D(n9031), .SP(clk_c_enable_283), 
            .CK(clk_c), .Q(\gpio_out_func_sel[0] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_0[[1__354 .GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_7[[0__390  (.D(n8876), .SP(clk_c_enable_284), 
            .CK(clk_c), .Q(\gpio_out_func_sel[7] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_7[[0__390 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_5[[1__379  (.D(\data_to_write[1] ), .SP(clk_c_enable_366), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[5] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_5[[1__379 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_2[[2__363  (.D(\data_to_write[2] ), .SP(clk_c_enable_359), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[2][2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_2[[2__363 .GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i12 (.D(baud_divider[11]), .SP(clk_c_enable_324), 
            .CD(n11704), .CK(clk_c), .Q(\peri_data_out[11] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i12.GSR = "DISABLED";
    FD1P3IX data_out_r_i0_i13 (.D(baud_divider[12]), .SP(clk_c_enable_324), 
            .CD(n11704), .CK(clk_c), .Q(\peri_data_out[12] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r_i0_i13.GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_5[[4__376  (.D(\data_to_write[4] ), .SP(clk_c_enable_366), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[5][4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_5[[4__376 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_1[[2__358  (.D(\data_to_write[2] ), .SP(clk_c_enable_358), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[1][2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_1[[2__358 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_6[[4__381  (.D(\data_to_write[4] ), .SP(clk_c_enable_355), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[6][4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_6[[4__381 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_5[[2__378  (.D(\data_to_write[2] ), .SP(clk_c_enable_366), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[5][2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_5[[2__378 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_4[[4__371  (.D(\data_to_write[4] ), .SP(clk_c_enable_353), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[4][4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_4[[4__371 .GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_3[[0__370  (.D(n8876), .SP(clk_c_enable_354), 
            .CK(clk_c), .Q(\gpio_out_func_sel[3] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_3[[0__370 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_6[[3__382  (.D(\data_to_write[3] ), .SP(clk_c_enable_355), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[6] [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_6[[3__382 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_0[[2__353  (.D(\data_to_write[2] ), .SP(clk_c_enable_356), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[0] [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_0[[2__353 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_1[[3__357  (.D(\data_to_write[3] ), .SP(clk_c_enable_358), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[1] [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_1[[3__357 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_1[[0__360  (.D(\data_to_write[0] ), .SP(clk_c_enable_358), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[1] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_1[[0__360 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_2[[1__364  (.D(\data_to_write[1] ), .SP(clk_c_enable_359), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[2] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_2[[1__364 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_5[[3__377  (.D(\data_to_write[3] ), .SP(clk_c_enable_366), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\gpio_out_func_sel[5] [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_5[[3__377 .GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_6[[0__385  (.D(n8876), .SP(clk_c_enable_368), 
            .CK(clk_c), .Q(\gpio_out_func_sel[6] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_6[[0__385 .GSR = "DISABLED";
    FD1P3AX data_ready_r_349 (.D(data_ready_r_N_2823), .SP(rst_reg_n), .CK(clk_c), 
            .Q(data_ready_r)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_ready_r_349.GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_4[[0__375  (.D(n8876), .SP(clk_c_enable_369), 
            .CK(clk_c), .Q(\gpio_out_func_sel[4]_c [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam \gpio_out_func_sel_4[[0__375 .GSR = "DISABLED";
    L6MUX21 i27562 (.D0(n30269), .D1(n30270), .SD(\addr[4] ), .Z(n30271));
    L6MUX21 i27569 (.D0(n30276), .D1(n30277), .SD(\addr[4] ), .Z(n30278));
    LUT4 i1_2_lut_rep_803 (.A(\addr[3] ), .B(\addr[2] ), .Z(n32818)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i1_2_lut_rep_803.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_704_3_lut_4_lut (.A(\addr[3] ), .B(\addr[2] ), .C(n32835), 
         .D(n32836), .Z(n32719)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i1_2_lut_rep_704_3_lut_4_lut.init = 16'hfffb;
    L6MUX21 i27576 (.D0(n30283), .D1(n30284), .SD(\addr[3] ), .Z(n30285));
    LUT4 i27573_3_lut (.A(\gpio_out_func_sel[6] [0]), .B(\gpio_out_func_sel[7] [0]), 
         .C(\addr[2] ), .Z(n30282)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27573_3_lut.init = 16'hcaca;
    LUT4 i27572_3_lut (.A(\gpio_out_func_sel[2] [0]), .B(\gpio_out_func_sel[3] [0]), 
         .C(\addr[2] ), .Z(n30281)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27572_3_lut.init = 16'hcaca;
    LUT4 mux_234_Mux_0_i3_4_lut (.A(\uo_out_from_user_peri[1]_c [1]), .B(\uo_out_from_user_peri[2] [7]), 
         .C(\gpio_out_func_sel[1] [1]), .D(\gpio_out_func_sel[1] [0]), .Z(n3_adj_3268)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(160[62:87])
    defparam mux_234_Mux_0_i3_4_lut.init = 16'h0ac0;
    LUT4 i27571_3_lut (.A(\gpio_out_func_sel[4]_c [0]), .B(\gpio_out_func_sel[5] [0]), 
         .C(\addr[2] ), .Z(n30280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27571_3_lut.init = 16'hcaca;
    LUT4 i27570_3_lut (.A(\gpio_out_func_sel[0] [0]), .B(\gpio_out_func_sel[1] [0]), 
         .C(\addr[2] ), .Z(n30279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27570_3_lut.init = 16'hcaca;
    LUT4 i27566_3_lut (.A(\gpio_out_func_sel[6] [1]), .B(\gpio_out_func_sel[7] [1]), 
         .C(\addr[2] ), .Z(n30275)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27566_3_lut.init = 16'hcaca;
    LUT4 i27565_3_lut (.A(\gpio_out_func_sel[4]_c [1]), .B(\gpio_out_func_sel[5] [1]), 
         .C(\addr[2] ), .Z(n30274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27565_3_lut.init = 16'hcaca;
    LUT4 i27564_3_lut (.A(\gpio_out_func_sel[2] [1]), .B(\gpio_out_func_sel[3] [1]), 
         .C(\addr[2] ), .Z(n30273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27564_3_lut.init = 16'hcaca;
    LUT4 i27563_3_lut (.A(\gpio_out_func_sel[0] [1]), .B(\gpio_out_func_sel[1] [1]), 
         .C(\addr[2] ), .Z(n30272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27563_3_lut.init = 16'hcaca;
    LUT4 i27559_3_lut (.A(\gpio_out_func_sel[6] [3]), .B(\gpio_out_func_sel[7] [3]), 
         .C(\addr[2] ), .Z(n30268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27559_3_lut.init = 16'hcaca;
    LUT4 i27558_3_lut (.A(\gpio_out_func_sel[4]_c [3]), .B(\gpio_out_func_sel[5] [3]), 
         .C(\addr[2] ), .Z(n30267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27558_3_lut.init = 16'hcaca;
    LUT4 i27557_3_lut (.A(\gpio_out_func_sel[2] [3]), .B(\gpio_out_func_sel[3] [3]), 
         .C(\addr[2] ), .Z(n30266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27557_3_lut.init = 16'hcaca;
    LUT4 i27556_3_lut (.A(\gpio_out_func_sel[0] [3]), .B(\gpio_out_func_sel[1] [3]), 
         .C(\addr[2] ), .Z(n30265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27556_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(\addr[2] ), .B(\addr[3] ), .Z(n10944)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i1_2_lut.init = 16'hbbbb;
    FD1P3IX gpio_out__i1 (.D(\data_to_write[1] ), .SP(clk_c_enable_463), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\uo_out_from_user_peri[1]_c [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(126[12] 134[8])
    defparam gpio_out__i1.GSR = "DISABLED";
    FD1P3IX gpio_out__i2 (.D(\data_to_write[2] ), .SP(clk_c_enable_463), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\uo_out_from_user_peri[1][2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(126[12] 134[8])
    defparam gpio_out__i2.GSR = "DISABLED";
    FD1P3IX gpio_out__i3 (.D(\data_to_write[3] ), .SP(clk_c_enable_463), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\uo_out_from_user_peri[1]_c [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(126[12] 134[8])
    defparam gpio_out__i3.GSR = "DISABLED";
    FD1P3IX gpio_out__i4 (.D(\data_to_write[4] ), .SP(clk_c_enable_463), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\uo_out_from_user_peri[1]_c [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(126[12] 134[8])
    defparam gpio_out__i4.GSR = "DISABLED";
    FD1P3IX gpio_out__i5 (.D(\data_to_write[5] ), .SP(clk_c_enable_463), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\uo_out_from_user_peri[1][5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(126[12] 134[8])
    defparam gpio_out__i5.GSR = "DISABLED";
    FD1P3IX gpio_out__i6 (.D(\data_to_write[6] ), .SP(clk_c_enable_463), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\uo_out_from_user_peri[1][6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(126[12] 134[8])
    defparam gpio_out__i6.GSR = "DISABLED";
    FD1P3IX gpio_out__i7 (.D(\data_to_write[7] ), .SP(clk_c_enable_463), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(\uo_out_from_user_peri[1]_c [7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(126[12] 134[8])
    defparam gpio_out__i7.GSR = "DISABLED";
    LUT4 i28550_4_lut (.A(n3_adj_3271), .B(\gpio_out_sel[7] ), .C(\gpio_out_func_sel[7][4] ), 
         .D(n6), .Z(uo_out_c_7)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(146[20] 154[16])
    defparam i28550_4_lut.init = 16'h0008;
    LUT4 mux_240_Mux_0_i3_4_lut (.A(\uo_out_from_user_peri[1]_c [7]), .B(\uo_out_from_user_peri[2] [7]), 
         .C(\gpio_out_func_sel[7] [1]), .D(\gpio_out_func_sel[7] [0]), .Z(n3_adj_3271)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(160[62:87])
    defparam mux_240_Mux_0_i3_4_lut.init = 16'h0ac0;
    LUT4 i1_2_lut_adj_613 (.A(\gpio_out_func_sel[7][2] ), .B(\gpio_out_func_sel[7] [3]), 
         .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_613.init = 16'heeee;
    LUT4 mux_3053_i3_4_lut (.A(\ui_in_sync[2] ), .B(n31883), .C(n32719), 
         .D(n26838), .Z(\data_from_user_peri_1__31__N_2455[2] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(137[45] 139[50])
    defparam mux_3053_i3_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_4_lut (.A(\addr[2] ), .B(led_state), .C(\addr[1] ), 
         .D(n27888), .Z(data_from_peri_31__N_2447[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(137[45:67])
    defparam i1_4_lut_4_lut.init = 16'h0400;
    LUT4 i28459_3_lut_4_lut (.A(n32693), .B(n32729), .C(rst_reg_n), .D(n32818), 
         .Z(clk_c_enable_100)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28459_3_lut_4_lut.init = 16'h0f1f;
    LUT4 i28285_3_lut_4_lut (.A(n32693), .B(n32729), .C(rst_reg_n), .D(n8854), 
         .Z(clk_c_enable_284)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28285_3_lut_4_lut.init = 16'h1f0f;
    LUT4 i28529_3_lut_4_lut (.A(n32693), .B(n32729), .C(rst_reg_n), .D(n10944), 
         .Z(clk_c_enable_368)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28529_3_lut_4_lut.init = 16'h0f1f;
    LUT4 i28524_3_lut_4_lut (.A(n32693), .B(n32729), .C(rst_reg_n), .D(n32819), 
         .Z(clk_c_enable_369)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28524_3_lut_4_lut.init = 16'h0f1f;
    LUT4 i22_3_lut (.A(n28053), .B(\debug_rd_r[0] ), .C(debug_register_data), 
         .Z(uo_out_c_2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(84[9:28])
    defparam i22_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(\gpio_out_func_sel[2] [3]), .B(\gpio_out_func_sel[2][4] ), 
         .C(n9), .D(\gpio_out_func_sel[2][2] ), .Z(n28053)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    LUT4 i23_4_lut (.A(\gpio_out_func_sel[2] [1]), .B(\gpio_out_func_sel[2] [0]), 
         .C(\uo_out_from_user_peri[2] [6]), .D(\uo_out_from_user_peri[1][2] ), 
         .Z(n9)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(84[9:28])
    defparam i23_4_lut.init = 16'h6420;
    LUT4 mux_3053_i2_4_lut (.A(\ui_in_sync[1] ), .B(n30278), .C(n32719), 
         .D(n32761), .Z(data_from_user_peri_1__31__N_2455[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(137[45] 139[50])
    defparam mux_3053_i2_4_lut.init = 16'h0aca;
    LUT4 mux_3053_i4_4_lut (.A(\ui_in_sync[3] ), .B(n30271), .C(n32719), 
         .D(n32761), .Z(data_from_user_peri_1__31__N_2455[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(137[45] 139[50])
    defparam mux_3053_i4_4_lut.init = 16'h0aca;
    LUT4 mux_3053_i5_4_lut (.A(\ui_in_sync[4] ), .B(n31794), .C(n32719), 
         .D(n26838), .Z(data_from_user_peri_1__31__N_2455[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(137[45] 139[50])
    defparam mux_3053_i5_4_lut.init = 16'hca0a;
    PFUMX i27560 (.BLUT(n30265), .ALUT(n30266), .C0(\addr[3] ), .Z(n30269));
    PFUMX i27561 (.BLUT(n30267), .ALUT(n30268), .C0(\addr[3] ), .Z(n30270));
    PFUMX i27567 (.BLUT(n30272), .ALUT(n30273), .C0(\addr[3] ), .Z(n30276));
    PFUMX i27568 (.BLUT(n30274), .ALUT(n30275), .C0(\addr[3] ), .Z(n30277));
    PFUMX i27574 (.BLUT(n30279), .ALUT(n30280), .C0(\addr[4] ), .Z(n30283));
    PFUMX i27575 (.BLUT(n30281), .ALUT(n30282), .C0(\addr[4] ), .Z(n30284));
    LUT4 mux_3053_i1_4_lut (.A(\ui_in_sync[0] ), .B(n32761), .C(n32719), 
         .D(n30285), .Z(\data_from_user_peri_1__31__N_2455[0] )) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(137[45] 139[50])
    defparam mux_3053_i1_4_lut.init = 16'h3a0a;
    LUT4 i8998_4_lut (.A(clk_c_enable_324), .B(n10944), .C(n32723), .D(n29531), 
         .Z(n11704)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam i8998_4_lut.init = 16'haaa8;
    LUT4 i28337_3_lut_4_lut (.A(n32727), .B(n32728), .C(n32720), .D(rst_reg_n), 
         .Z(clk_c_enable_463)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C (D))))) */ ;
    defparam i28337_3_lut_4_lut.init = 16'h01ff;
    LUT4 i1_2_lut_rep_664_4_lut (.A(n12), .B(n32737), .C(data_out_hold), 
         .D(rst_reg_n), .Z(clk_c_enable_324)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_664_4_lut.init = 16'h0200;
    LUT4 i3_4_lut_adj_614 (.A(n3_adj_3272), .B(\gpio_out_func_sel[3][4] ), 
         .C(\gpio_out_func_sel[3][2] ), .D(\gpio_out_func_sel[3] [3]), .Z(\peri_out[3] )) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut_adj_614.init = 16'h0002;
    LUT4 mux_236_Mux_0_i3_4_lut (.A(\uo_out_from_user_peri[1]_c [3]), .B(\uo_out_from_user_peri[2] [7]), 
         .C(\gpio_out_func_sel[3] [1]), .D(\gpio_out_func_sel[3] [0]), .Z(n3_adj_3272)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(160[62:87])
    defparam mux_236_Mux_0_i3_4_lut.init = 16'h0ac0;
    LUT4 i15187_4_lut (.A(\uo_out_from_user_peri[1]_c [7]), .B(\addr[6] ), 
         .C(\data_from_user_peri_1__31__N_2455[7] ), .D(n32720), .Z(n1_adj_3269)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(111[50:62])
    defparam i15187_4_lut.init = 16'hc088;
    LUT4 i3_4_lut_adj_615 (.A(n3_adj_3273), .B(\gpio_out_func_sel[4]_c [3]), 
         .C(\gpio_out_func_sel[4] [2]), .D(\gpio_out_func_sel[4][4] ), .Z(\peri_out[4] )) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut_adj_615.init = 16'h0002;
    LUT4 mux_237_Mux_0_i3_4_lut (.A(\uo_out_from_user_peri[1]_c [4]), .B(\uo_out_from_user_peri[2] [6]), 
         .C(\gpio_out_func_sel[4]_c [1]), .D(\gpio_out_func_sel[4]_c [0]), 
         .Z(n3_adj_3273)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(160[62:87])
    defparam mux_237_Mux_0_i3_4_lut.init = 16'h0ac0;
    LUT4 i15024_2_lut_rep_651_3_lut_4_lut (.A(n32819), .B(n32757), .C(n32801), 
         .D(n8109), .Z(n32666)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(137[45:67])
    defparam i15024_2_lut_rep_651_3_lut_4_lut.init = 16'hfeff;
    LUT4 i28503_2_lut_3_lut_4_lut (.A(n32761), .B(\addr[4] ), .C(n32819), 
         .D(n32700), .Z(clk_c_enable_356)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28503_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i28500_2_lut_3_lut_4_lut (.A(n32761), .B(\addr[4] ), .C(n8854), 
         .D(n32700), .Z(clk_c_enable_278)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28500_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i28509_2_lut_3_lut_4_lut (.A(n32761), .B(\addr[4] ), .C(n10944), 
         .D(n32700), .Z(clk_c_enable_359)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28509_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i28498_2_lut_3_lut_4_lut (.A(n32761), .B(\addr[4] ), .C(n32818), 
         .D(n32700), .Z(clk_c_enable_358)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28498_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i3_4_lut_adj_616 (.A(n3_adj_3274), .B(\gpio_out_func_sel[5][4] ), 
         .C(\gpio_out_func_sel[5][2] ), .D(\gpio_out_func_sel[5] [3]), .Z(\peri_out[5] )) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut_adj_616.init = 16'h0002;
    LUT4 mux_238_Mux_0_i3_4_lut (.A(\uo_out_from_user_peri[1][5] ), .B(\uo_out_from_user_peri[2] [7]), 
         .C(\gpio_out_func_sel[5] [1]), .D(\gpio_out_func_sel[5] [0]), .Z(n3_adj_3274)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(160[62:87])
    defparam mux_238_Mux_0_i3_4_lut.init = 16'h0ac0;
    LUT4 i3_4_lut_adj_617 (.A(n3_adj_3275), .B(\gpio_out_func_sel[6][2] ), 
         .C(\gpio_out_func_sel[6][4] ), .D(\gpio_out_func_sel[6] [3]), .Z(\peri_out[6] )) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut_adj_617.init = 16'h0002;
    LUT4 mux_239_Mux_0_i3_4_lut (.A(\uo_out_from_user_peri[1][6] ), .B(\uo_out_from_user_peri[2] [6]), 
         .C(\gpio_out_func_sel[6] [1]), .D(\gpio_out_func_sel[6] [0]), .Z(n3_adj_3275)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(160[62:87])
    defparam mux_239_Mux_0_i3_4_lut.init = 16'h0ac0;
    LUT4 i28331_2_lut_rep_658_3_lut_4_lut (.A(n10944), .B(n32757), .C(n32801), 
         .D(n8109), .Z(clk_c_enable_64)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(136[45:67])
    defparam i28331_2_lut_rep_658_3_lut_4_lut.init = 16'h0100;
    LUT4 i28512_2_lut_3_lut_4_lut (.A(n32761), .B(\addr[4] ), .C(n10944), 
         .D(n32700), .Z(clk_c_enable_355)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28512_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i28514_2_lut_3_lut_4_lut (.A(n32761), .B(\addr[4] ), .C(n8854), 
         .D(n32700), .Z(clk_c_enable_270)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28514_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i28517_2_lut_3_lut_4_lut (.A(n32761), .B(\addr[4] ), .C(n32819), 
         .D(n32700), .Z(clk_c_enable_353)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28517_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i28506_2_lut_3_lut_4_lut (.A(n32761), .B(\addr[4] ), .C(n32818), 
         .D(n32700), .Z(clk_c_enable_366)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(138[45:83])
    defparam i28506_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i15191_4_lut (.A(\uo_out_from_user_peri[1]_c [4]), .B(\addr[6] ), 
         .C(data_from_user_peri_1__31__N_2455[4]), .D(n32720), .Z(n1_adj_3266)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(111[50:62])
    defparam i15191_4_lut.init = 16'hc088;
    LUT4 i15192_4_lut (.A(\uo_out_from_user_peri[1]_c [3]), .B(\addr[6] ), 
         .C(data_from_user_peri_1__31__N_2455[3]), .D(n32720), .Z(n1_adj_3264)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(111[50:62])
    defparam i15192_4_lut.init = 16'hc088;
    LUT4 i15197_4_lut (.A(\uo_out_from_user_peri[1]_c [1]), .B(\addr[6] ), 
         .C(data_from_user_peri_1__31__N_2455[1]), .D(n32720), .Z(n1)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(111[50:62])
    defparam i15197_4_lut.init = 16'hc088;
    PFUMX mux_5202_i1 (.BLUT(\data_from_peri_31__N_2415[0] ), .ALUT(data_from_peri_31__N_2447[0]), 
          .C0(\addr[10] ), .Z(data_from_peri[0]));
    \tqvp_uart_wrapper(CLOCK_MHZ=25)  i_uart (.baud_divider({baud_divider}), 
            .clk_c(clk_c), .clk_c_enable_432(clk_c_enable_432), .\data_to_write[4] (\data_to_write[4] ), 
            .\data_to_write[6] (\data_to_write[6] ), .\data_to_write[7] (\data_to_write[7] ), 
            .\data_to_write[12] (\data_to_write[12] ), .\data_to_write[11] (\data_to_write[11] ), 
            .\data_to_write[10] (\data_to_write[10] ), .\data_to_write[9] (\data_to_write[9] ), 
            .\data_to_write[8] (\data_to_write[8] ), .clk_c_enable_64(clk_c_enable_64), 
            .\data_to_write[5] (\data_to_write[5] ), .\data_to_write[2] (\data_to_write[2] ), 
            .\data_to_write[1] (\data_to_write[1] ), .\data_to_write[0] (\data_to_write[0] ), 
            .\ui_in_sync[7] (\ui_in_sync[7] ), .\ui_in_sync[3] (\ui_in_sync[3] ), 
            .\addr[2] (\addr[2] ), .n31706(n31706), .\uart_rx_buf_data[2] (\uart_rx_buf_data[2] ), 
            .\uart_rx_buf_data[3] (\uart_rx_buf_data[3] ), .\uart_rx_buf_data[4] (\uart_rx_buf_data[4] ), 
            .\uart_rx_buf_data[5] (\uart_rx_buf_data[5] ), .\uart_rx_buf_data[6] (\uart_rx_buf_data[6] ), 
            .\uart_rx_buf_data[7] (\uart_rx_buf_data[7] ), .\addr[3] (\addr[3] ), 
            .\next_fsm_state_3__N_3046[3] (\next_fsm_state_3__N_3046[3] ), 
            .n31795(n31795), .n31796(n31796), .\addr[4] (\addr[4] ), .\addr[5] (\addr[5] ), 
            .n32836(n32836), .\addr[7] (\addr[7] ), .n29531(n29531), .\addr[0] (\addr[0] ), 
            .\addr[1] (\addr[1] ), .n32757(n32757), .n32720(n32720), .n32695(n32695), 
            .rst_reg_n(rst_reg_n), .n32730(n32730), .n26870(n26870), .\data_to_write[3] (\data_to_write[3] ), 
            .n8109(n8109), .n32725(n32725), .qv_data_write_n({qv_data_write_n}), 
            .n32710(n32710), .\imm[6] (\imm[6] ), .\csr_read_3__N_1447[2] (\csr_read_3__N_1447[2] ), 
            .n29866(n29866), .n32801(n32801), .n29491(n29491), .n8854(n8854), 
            .cycle_counter({cycle_counter}), .n72({n72}), .n32791(n32791), 
            .fsm_state({fsm_state}), .next_bit(next_bit), .\uo_out_from_user_peri[2][6] (\uo_out_from_user_peri[2] [6]), 
            .n32666(n32666), .\gpio_out_func_sel[0][0] (\gpio_out_func_sel[0] [0]), 
            .\gpio_out_func_sel[0][4] (\gpio_out_func_sel[0] [4]), .n27757(n27757), 
            .n32763(n32763), .n32251(n32251), .GND_net(GND_net), .VCC_net(VCC_net), 
            .cycle_counter_adj_46({cycle_counter_adj_65}), .next_bit_adj_43(next_bit_adj_62), 
            .\uo_out_from_user_peri[2][7] (\uo_out_from_user_peri[2] [7]), 
            .debug_stop_txn(debug_stop_txn), .instr_active_N_2106(instr_active_N_2106), 
            .stop_txn_reg(stop_txn_reg), .n32755(n32755), .stop_txn_now_N_2363(stop_txn_now_N_2363), 
            .clk_c_enable_208(clk_c_enable_208), .n32714(n32714), .qspi_write_done(qspi_write_done), 
            .n10672(n10672), .spi_clk_pos(spi_clk_pos), .n28259(n28259), 
            .next_bit_adj_44(next_bit_adj_63), .n32622(n32622), .uart_txd_N_3005(uart_txd_N_3005), 
            .clk_c_enable_495(clk_c_enable_495), .n32832(n32832), .\fsm_state[0]_adj_45 (\fsm_state[0]_adj_64 ), 
            .clk_c_enable_143(clk_c_enable_143), .n9031(n9031), .n762(n762), 
            .clk_c_enable_519(clk_c_enable_519), .n8177(n8177), .n32524(n32524), 
            .n29357(n29357), .n46(n46), .n32728(n32728), .clk_c_enable_286(clk_c_enable_286), 
            .instr_complete_N_1647(instr_complete_N_1647), .n28957(n28957), 
            .n32706(n32706), .clk_c_enable_6(clk_c_enable_6), .n8876(n8876), 
            .n32771(n32771), .n27178(n27178), .n29549(n29549), .clk_c_enable_282(clk_c_enable_282), 
            .n6142(n6142), .n28319(n28319), .n32681(n32681), .n27931(n27931), 
            .n1072(n1072), .clk_c_enable_543(clk_c_enable_543), .qv_data_read_n({qv_data_read_n}), 
            .n26691(n26691), .\qspi_data_in[1] (\qspi_data_in[1] ), .\qspi_data_out_3__N_5[1] (\qspi_data_out_3__N_5[1] ), 
            .n26692(n26692)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(194[45] 206[3])
    tqvp_led_byte i_led_byte (.led_state(led_state), .clk_c(clk_c), .clk_c_enable_282(clk_c_enable_282), 
            .clk_c_enable_432(clk_c_enable_432), .\data_to_write[0] (\data_to_write[0] )) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(250[16] 264[3])
    
endmodule
//
// Verilog Description of module \tqvp_uart_wrapper(CLOCK_MHZ=25) 
//

module \tqvp_uart_wrapper(CLOCK_MHZ=25)  (baud_divider, clk_c, clk_c_enable_432, 
            \data_to_write[4] , \data_to_write[6] , \data_to_write[7] , 
            \data_to_write[12] , \data_to_write[11] , \data_to_write[10] , 
            \data_to_write[9] , \data_to_write[8] , clk_c_enable_64, \data_to_write[5] , 
            \data_to_write[2] , \data_to_write[1] , \data_to_write[0] , 
            \ui_in_sync[7] , \ui_in_sync[3] , \addr[2] , n31706, \uart_rx_buf_data[2] , 
            \uart_rx_buf_data[3] , \uart_rx_buf_data[4] , \uart_rx_buf_data[5] , 
            \uart_rx_buf_data[6] , \uart_rx_buf_data[7] , \addr[3] , \next_fsm_state_3__N_3046[3] , 
            n31795, n31796, \addr[4] , \addr[5] , n32836, \addr[7] , 
            n29531, \addr[0] , \addr[1] , n32757, n32720, n32695, 
            rst_reg_n, n32730, n26870, \data_to_write[3] , n8109, 
            n32725, qv_data_write_n, n32710, \imm[6] , \csr_read_3__N_1447[2] , 
            n29866, n32801, n29491, n8854, cycle_counter, n72, n32791, 
            fsm_state, next_bit, \uo_out_from_user_peri[2][6] , n32666, 
            \gpio_out_func_sel[0][0] , \gpio_out_func_sel[0][4] , n27757, 
            n32763, n32251, GND_net, VCC_net, cycle_counter_adj_46, 
            next_bit_adj_43, \uo_out_from_user_peri[2][7] , debug_stop_txn, 
            instr_active_N_2106, stop_txn_reg, n32755, stop_txn_now_N_2363, 
            clk_c_enable_208, n32714, qspi_write_done, n10672, spi_clk_pos, 
            n28259, next_bit_adj_44, n32622, uart_txd_N_3005, clk_c_enable_495, 
            n32832, \fsm_state[0]_adj_45 , clk_c_enable_143, n9031, 
            n762, clk_c_enable_519, n8177, n32524, n29357, n46, 
            n32728, clk_c_enable_286, instr_complete_N_1647, n28957, 
            n32706, clk_c_enable_6, n8876, n32771, n27178, n29549, 
            clk_c_enable_282, n6142, n28319, n32681, n27931, n1072, 
            clk_c_enable_543, qv_data_read_n, n26691, \qspi_data_in[1] , 
            \qspi_data_out_3__N_5[1] , n26692) /* synthesis syn_module_defined=1 */ ;
    output [12:0]baud_divider;
    input clk_c;
    output clk_c_enable_432;
    input \data_to_write[4] ;
    input \data_to_write[6] ;
    input \data_to_write[7] ;
    input \data_to_write[12] ;
    input \data_to_write[11] ;
    input \data_to_write[10] ;
    input \data_to_write[9] ;
    input \data_to_write[8] ;
    input clk_c_enable_64;
    input \data_to_write[5] ;
    input \data_to_write[2] ;
    input \data_to_write[1] ;
    input \data_to_write[0] ;
    input \ui_in_sync[7] ;
    input \ui_in_sync[3] ;
    input \addr[2] ;
    output n31706;
    output \uart_rx_buf_data[2] ;
    output \uart_rx_buf_data[3] ;
    output \uart_rx_buf_data[4] ;
    output \uart_rx_buf_data[5] ;
    output \uart_rx_buf_data[6] ;
    output \uart_rx_buf_data[7] ;
    input \addr[3] ;
    output \next_fsm_state_3__N_3046[3] ;
    output n31795;
    output n31796;
    input \addr[4] ;
    input \addr[5] ;
    output n32836;
    input \addr[7] ;
    output n29531;
    input \addr[0] ;
    input \addr[1] ;
    output n32757;
    input n32720;
    input n32695;
    input rst_reg_n;
    input n32730;
    input n26870;
    input \data_to_write[3] ;
    input n8109;
    input n32725;
    input [1:0]qv_data_write_n;
    input n32710;
    input \imm[6] ;
    input \csr_read_3__N_1447[2] ;
    output n29866;
    input n32801;
    input n29491;
    input n8854;
    output [12:0]cycle_counter;
    input [12:0]n72;
    input n32791;
    output [3:0]fsm_state;
    input next_bit;
    output \uo_out_from_user_peri[2][6] ;
    input n32666;
    input \gpio_out_func_sel[0][0] ;
    input \gpio_out_func_sel[0][4] ;
    output n27757;
    input n32763;
    output n32251;
    input GND_net;
    input VCC_net;
    output [12:0]cycle_counter_adj_46;
    input next_bit_adj_43;
    output \uo_out_from_user_peri[2][7] ;
    input debug_stop_txn;
    output instr_active_N_2106;
    input stop_txn_reg;
    input n32755;
    input stop_txn_now_N_2363;
    output clk_c_enable_208;
    input n32714;
    input qspi_write_done;
    output n10672;
    input spi_clk_pos;
    output n28259;
    input next_bit_adj_44;
    input n32622;
    input uart_txd_N_3005;
    output clk_c_enable_495;
    input n32832;
    input \fsm_state[0]_adj_45 ;
    output clk_c_enable_143;
    output n9031;
    input n762;
    output clk_c_enable_519;
    output n8177;
    output n32524;
    input n29357;
    input n46;
    input n32728;
    output clk_c_enable_286;
    input instr_complete_N_1647;
    input n28957;
    input n32706;
    output clk_c_enable_6;
    output n8876;
    input n32771;
    input n27178;
    input n29549;
    output clk_c_enable_282;
    output n6142;
    input n28319;
    input n32681;
    output n27931;
    input n1072;
    output clk_c_enable_543;
    input [1:0]qv_data_read_n;
    output n26691;
    input \qspi_data_in[1] ;
    output \qspi_data_out_3__N_5[1] ;
    output n26692;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire clk_c_enable_544, clk_c_enable_61;
    wire [7:0]uart_rx_buf_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(98[15:31])
    
    wire clk_c_enable_451;
    wire [7:0]uart_rx_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(81[16:28])
    
    wire rxd_select, clk_c_enable_327, n32803, mid_bit;
    wire [3:0]next_fsm_state_3__N_3042;
    
    wire n17837, n26872, clk_c_enable_526, n27992, n32636, n29569;
    wire [3:0]fsm_state_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(47[11:20])
    
    wire clk_c_enable_269, n6162, clk_c_enable_515, uart_txd_N_3005_c;
    
    FD1P3JX baud_divider_i4 (.D(\data_to_write[4] ), .SP(clk_c_enable_544), 
            .PD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[4])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i4.GSR = "DISABLED";
    FD1P3JX baud_divider_i6 (.D(\data_to_write[6] ), .SP(clk_c_enable_544), 
            .PD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[6])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i6.GSR = "DISABLED";
    FD1P3JX baud_divider_i7 (.D(\data_to_write[7] ), .SP(clk_c_enable_544), 
            .PD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[7])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i7.GSR = "DISABLED";
    FD1P3IX baud_divider_i12 (.D(\data_to_write[12] ), .SP(clk_c_enable_61), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[12])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i12.GSR = "DISABLED";
    FD1P3IX baud_divider_i11 (.D(\data_to_write[11] ), .SP(clk_c_enable_61), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[11])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i11.GSR = "DISABLED";
    FD1P3IX baud_divider_i10 (.D(\data_to_write[10] ), .SP(clk_c_enable_61), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[10])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i10.GSR = "DISABLED";
    FD1P3IX baud_divider_i9 (.D(\data_to_write[9] ), .SP(clk_c_enable_61), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[9])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i9.GSR = "DISABLED";
    FD1P3IX baud_divider_i8 (.D(\data_to_write[8] ), .SP(clk_c_enable_61), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[8])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i8.GSR = "DISABLED";
    FD1P3IX baud_divider_i5 (.D(\data_to_write[5] ), .SP(clk_c_enable_64), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[5])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i5.GSR = "DISABLED";
    FD1P3IX baud_divider_i2 (.D(\data_to_write[2] ), .SP(clk_c_enable_64), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[2])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i2.GSR = "DISABLED";
    FD1P3IX baud_divider_i1 (.D(\data_to_write[1] ), .SP(clk_c_enable_64), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[1])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i1.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i0 (.D(uart_rx_data[0]), .SP(clk_c_enable_451), 
            .CK(clk_c), .Q(uart_rx_buf_data[0])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i0.GSR = "DISABLED";
    FD1P3IX rxd_select_58 (.D(\data_to_write[0] ), .SP(clk_c_enable_327), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(rxd_select)) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(50[12] 58[8])
    defparam rxd_select_58.GSR = "DISABLED";
    LUT4 ui_in_7__I_0_3_lut_rep_788 (.A(\ui_in_sync[7] ), .B(\ui_in_sync[3] ), 
         .C(rxd_select), .Z(n32803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(82[21:53])
    defparam ui_in_7__I_0_3_lut_rep_788.init = 16'hcaca;
    LUT4 i15452_2_lut_4_lut (.A(\ui_in_sync[7] ), .B(\ui_in_sync[3] ), .C(rxd_select), 
         .D(mid_bit), .Z(next_fsm_state_3__N_3042[1])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(82[21:53])
    defparam i15452_2_lut_4_lut.init = 16'hcaff;
    LUT4 uart_tx_busy_bdd_3_lut_28845 (.A(baud_divider[0]), .B(rxd_select), 
         .C(\addr[2] ), .Z(n31706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam uart_tx_busy_bdd_3_lut_28845.init = 16'hcaca;
    FD1P3AX uart_rx_buf_data_i0_i1 (.D(uart_rx_data[1]), .SP(clk_c_enable_451), 
            .CK(clk_c), .Q(uart_rx_buf_data[1])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i1.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i2 (.D(uart_rx_data[2]), .SP(clk_c_enable_451), 
            .CK(clk_c), .Q(\uart_rx_buf_data[2] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i2.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i3 (.D(uart_rx_data[3]), .SP(clk_c_enable_451), 
            .CK(clk_c), .Q(\uart_rx_buf_data[3] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i3.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i4 (.D(uart_rx_data[4]), .SP(clk_c_enable_451), 
            .CK(clk_c), .Q(\uart_rx_buf_data[4] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i4.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i5 (.D(uart_rx_data[5]), .SP(clk_c_enable_451), 
            .CK(clk_c), .Q(\uart_rx_buf_data[5] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i5.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i6 (.D(uart_rx_data[6]), .SP(clk_c_enable_451), 
            .CK(clk_c), .Q(\uart_rx_buf_data[6] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i6.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i7 (.D(uart_rx_data[7]), .SP(clk_c_enable_451), 
            .CK(clk_c), .Q(\uart_rx_buf_data[7] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i7.GSR = "DISABLED";
    LUT4 addr_2__bdd_2_lut (.A(\addr[3] ), .B(\next_fsm_state_3__N_3046[3] ), 
         .Z(n31795)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam addr_2__bdd_2_lut.init = 16'h4444;
    LUT4 addr_2__bdd_3_lut (.A(uart_rx_buf_data[1]), .B(\addr[3] ), .C(baud_divider[1]), 
         .Z(n31796)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam addr_2__bdd_3_lut.init = 16'he2e2;
    LUT4 i15559_2_lut_rep_821 (.A(\addr[4] ), .B(\addr[5] ), .Z(n32836)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15559_2_lut_rep_821.init = 16'heeee;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\addr[4] ), .B(\addr[5] ), .C(\addr[7] ), 
         .Z(n29531)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_742_3_lut_4_lut (.A(\addr[4] ), .B(\addr[5] ), .C(\addr[0] ), 
         .D(\addr[1] ), .Z(n32757)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_742_3_lut_4_lut.init = 16'hfffe;
    LUT4 i28359_3_lut_4_lut (.A(n32720), .B(n32695), .C(rst_reg_n), .D(n32730), 
         .Z(n17837)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B (C)))) */ ;
    defparam i28359_3_lut_4_lut.init = 16'h0fef;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32720), .B(n32695), .C(n26870), .D(n32730), 
         .Z(n26872)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    FD1P3AX uart_rx_buffered_59 (.D(n27992), .SP(clk_c_enable_526), .CK(clk_c), 
            .Q(\next_fsm_state_3__N_3046[3] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buffered_59.GSR = "DISABLED";
    FD1P3JX baud_divider_i0 (.D(\data_to_write[0] ), .SP(clk_c_enable_544), 
            .PD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[0])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i0.GSR = "DISABLED";
    FD1P3JX baud_divider_i3 (.D(\data_to_write[3] ), .SP(clk_c_enable_544), 
            .PD(clk_c_enable_432), .CK(clk_c), .Q(baud_divider[3])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=194, LSE_RLINE=206 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i3.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n8109), .B(n32725), .C(qv_data_write_n[1]), .D(qv_data_write_n[0]), 
         .Z(clk_c_enable_61)) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(41[13] 44[16])
    defparam i1_4_lut.init = 16'h0220;
    LUT4 i27948_3_lut_4_lut (.A(\next_fsm_state_3__N_3046[3] ), .B(n32710), 
         .C(\imm[6] ), .D(\csr_read_3__N_1447[2] ), .Z(n29866)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam i27948_3_lut_4_lut.init = 16'h8f80;
    LUT4 i15026_2_lut_rep_621_3_lut_4_lut (.A(n8109), .B(n32801), .C(n32730), 
         .D(n32720), .Z(n32636)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i15026_2_lut_rep_621_3_lut_4_lut.init = 16'hfffd;
    LUT4 i28461_2_lut_3_lut_4_lut (.A(n8109), .B(n32801), .C(rst_reg_n), 
         .D(n32725), .Z(clk_c_enable_544)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C))) */ ;
    defparam i28461_2_lut_3_lut_4_lut.init = 16'h0f2f;
    LUT4 i572_2_lut (.A(\next_fsm_state_3__N_3046[3] ), .B(rst_reg_n), .Z(clk_c_enable_451)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(103[18] 112[12])
    defparam i572_2_lut.init = 16'h4444;
    LUT4 i28391_4_lut (.A(rst_reg_n), .B(n29491), .C(\next_fsm_state_3__N_3046[3] ), 
         .D(n32720), .Z(clk_c_enable_526)) /* synthesis lut_function=(!(A (B (C)+!B (C (D))))) */ ;
    defparam i28391_4_lut.init = 16'h5f7f;
    LUT4 i1_4_lut_adj_612 (.A(\next_fsm_state_3__N_3046[3] ), .B(rst_reg_n), 
         .C(n29569), .D(fsm_state_c[2]), .Z(n27992)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_612.init = 16'h0040;
    LUT4 i1_3_lut (.A(fsm_state_c[0]), .B(fsm_state_c[3]), .C(fsm_state_c[1]), 
         .Z(n29569)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i28299_4_lut (.A(n32695), .B(rst_reg_n), .C(n8854), .D(n32757), 
         .Z(clk_c_enable_327)) /* synthesis lut_function=(!(A+(B ((D)+!C)))) */ ;
    defparam i28299_4_lut.init = 16'h1151;
    tqvp_uart_tx i_uart_tx (.cycle_counter({cycle_counter}), .clk_c(clk_c), 
            .clk_c_enable_269(clk_c_enable_269), .n6162(n6162), .n72({n72}), 
            .n32791(n32791), .fsm_state({fsm_state}), .rst_reg_n(rst_reg_n), 
            .next_bit(next_bit), .n17837(n17837), .\uo_out_from_user_peri[2][6] (\uo_out_from_user_peri[2][6] ), 
            .clk_c_enable_432(clk_c_enable_432), .n32730(n32730), .n32666(n32666), 
            .\data_to_write[0] (\data_to_write[0] ), .\data_to_write[6] (\data_to_write[6] ), 
            .\data_to_write[5] (\data_to_write[5] ), .\data_to_write[4] (\data_to_write[4] ), 
            .\data_to_write[3] (\data_to_write[3] ), .\data_to_write[2] (\data_to_write[2] ), 
            .\data_to_write[1] (\data_to_write[1] ), .clk_c_enable_515(clk_c_enable_515), 
            .n26872(n26872), .\gpio_out_func_sel[0][0] (\gpio_out_func_sel[0][0] ), 
            .\gpio_out_func_sel[0][4] (\gpio_out_func_sel[0][4] ), .n27757(n27757), 
            .uart_txd_N_3005(uart_txd_N_3005_c), .n32763(n32763), .\addr[2] (\addr[2] ), 
            .\uart_rx_buf_data[0] (uart_rx_buf_data[0]), .n32251(n32251)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(65[18] 73[6])
    tqvp_uart_rx i_uart_rx (.GND_net(GND_net), .VCC_net(VCC_net), .cycle_counter({cycle_counter_adj_46}), 
            .\baud_divider[8] (baud_divider[8]), .\baud_divider[7] (baud_divider[7]), 
            .\baud_divider[6] (baud_divider[6]), .\baud_divider[5] (baud_divider[5]), 
            .mid_bit(mid_bit), .\baud_divider[4] (baud_divider[4]), .\baud_divider[3] (baud_divider[3]), 
            .\baud_divider[2] (baud_divider[2]), .\baud_divider[1] (baud_divider[1]), 
            .\baud_divider[12] (baud_divider[12]), .\baud_divider[11] (baud_divider[11]), 
            .\baud_divider[10] (baud_divider[10]), .\baud_divider[9] (baud_divider[9]), 
            .\next_fsm_state_3__N_3046[3] (\next_fsm_state_3__N_3046[3] ), 
            .fsm_state({fsm_state_c}), .next_bit(next_bit_adj_43), .n32803(n32803), 
            .clk_c(clk_c), .clk_c_enable_432(clk_c_enable_432), .uart_rx_data({uart_rx_data}), 
            .\uo_out_from_user_peri[2][7] (\uo_out_from_user_peri[2][7] ), 
            .rst_reg_n(rst_reg_n), .debug_stop_txn(debug_stop_txn), .instr_active_N_2106(instr_active_N_2106), 
            .next_bit_adj_25(next_bit), .n32763(n32763), .\fsm_state[0]_adj_26 (fsm_state[0]), 
            .clk_c_enable_269(clk_c_enable_269), .stop_txn_reg(stop_txn_reg), 
            .n32755(n32755), .stop_txn_now_N_2363(stop_txn_now_N_2363), 
            .clk_c_enable_208(clk_c_enable_208), .n6162(n6162), .n32714(n32714), 
            .qspi_write_done(qspi_write_done), .n10672(n10672), .spi_clk_pos(spi_clk_pos), 
            .n28259(n28259), .next_bit_adj_27(next_bit_adj_44), .n32622(n32622), 
            .uart_txd_N_3005(uart_txd_N_3005), .clk_c_enable_495(clk_c_enable_495), 
            .n32832(n32832), .\fsm_state[0]_adj_28 (\fsm_state[0]_adj_45 ), 
            .clk_c_enable_143(clk_c_enable_143), .\data_to_write[1] (\data_to_write[1] ), 
            .n9031(n9031), .n762(n762), .clk_c_enable_519(clk_c_enable_519), 
            .n8177(n8177), .n32524(n32524), .n29357(n29357), .n46(n46), 
            .n32728(n32728), .clk_c_enable_286(clk_c_enable_286), .instr_complete_N_1647(instr_complete_N_1647), 
            .n28957(n28957), .n32706(n32706), .clk_c_enable_6(clk_c_enable_6), 
            .\data_to_write[0] (\data_to_write[0] ), .n8876(n8876), .n32771(n32771), 
            .n27178(n27178), .n29549(n29549), .clk_c_enable_282(clk_c_enable_282), 
            .n32636(n32636), .uart_txd_N_3005_adj_29(uart_txd_N_3005_c), 
            .clk_c_enable_515(clk_c_enable_515), .n6142(n6142), .n28319(n28319), 
            .n32681(n32681), .n27931(n27931), .n1072(n1072), .clk_c_enable_543(clk_c_enable_543), 
            .qv_data_read_n({qv_data_read_n}), .qv_data_write_n({qv_data_write_n}), 
            .n26691(n26691), .\qspi_data_in[1] (\qspi_data_in[1] ), .\qspi_data_out_3__N_5[1] (\qspi_data_out_3__N_5[1] ), 
            .n26692(n26692), .\next_fsm_state_3__N_3042[1] (next_fsm_state_3__N_3042[1])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(85[18] 94[6])
    
endmodule
//
// Verilog Description of module tqvp_uart_tx
//

module tqvp_uart_tx (cycle_counter, clk_c, clk_c_enable_269, n6162, 
            n72, n32791, fsm_state, rst_reg_n, next_bit, n17837, 
            \uo_out_from_user_peri[2][6] , clk_c_enable_432, n32730, n32666, 
            \data_to_write[0] , \data_to_write[6] , \data_to_write[5] , 
            \data_to_write[4] , \data_to_write[3] , \data_to_write[2] , 
            \data_to_write[1] , clk_c_enable_515, n26872, \gpio_out_func_sel[0][0] , 
            \gpio_out_func_sel[0][4] , n27757, uart_txd_N_3005, n32763, 
            \addr[2] , \uart_rx_buf_data[0] , n32251) /* synthesis syn_module_defined=1 */ ;
    output [12:0]cycle_counter;
    input clk_c;
    input clk_c_enable_269;
    input n6162;
    input [12:0]n72;
    input n32791;
    output [3:0]fsm_state;
    input rst_reg_n;
    input next_bit;
    input n17837;
    output \uo_out_from_user_peri[2][6] ;
    input clk_c_enable_432;
    input n32730;
    input n32666;
    input \data_to_write[0] ;
    input \data_to_write[6] ;
    input \data_to_write[5] ;
    input \data_to_write[4] ;
    input \data_to_write[3] ;
    input \data_to_write[2] ;
    input \data_to_write[1] ;
    input clk_c_enable_515;
    input n26872;
    input \gpio_out_func_sel[0][0] ;
    input \gpio_out_func_sel[0][4] ;
    output n27757;
    output uart_txd_N_3005;
    input n32763;
    input \addr[2] ;
    input \uart_rx_buf_data[0] ;
    output n32251;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n32684, n31502, clk_c_enable_271, n32865, n31493;
    wire [3:0]n162;
    
    wire uart_txd_N_3003;
    wire [7:0]data_to_send;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(39[24:36])
    wire [7:0]data_to_send_7__N_2975;
    
    FD1P3IX cycle_counter__i0 (.D(n72[0]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i0.GSR = "DISABLED";
    LUT4 i28493_2_lut_rep_669_3_lut_4_lut (.A(n32791), .B(fsm_state[2]), 
         .C(rst_reg_n), .D(fsm_state[0]), .Z(n32684)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(72[17:37])
    defparam i28493_2_lut_rep_669_3_lut_4_lut.init = 16'h0f1f;
    FD1P3IX cycle_counter__i12 (.D(n72[12]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[12])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i12.GSR = "DISABLED";
    FD1P3IX cycle_counter__i11 (.D(n72[11]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[11])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i11.GSR = "DISABLED";
    FD1P3IX cycle_counter__i10 (.D(n72[10]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[10])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i10.GSR = "DISABLED";
    FD1P3IX cycle_counter__i9 (.D(n72[9]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[9])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i9.GSR = "DISABLED";
    FD1P3IX cycle_counter__i8 (.D(n72[8]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[8])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i8.GSR = "DISABLED";
    FD1P3IX cycle_counter__i7 (.D(n72[7]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[7])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i7.GSR = "DISABLED";
    FD1P3IX cycle_counter__i6 (.D(n72[6]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[6])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i6.GSR = "DISABLED";
    FD1P3IX cycle_counter__i5 (.D(n72[5]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[5])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i5.GSR = "DISABLED";
    FD1P3IX cycle_counter__i4 (.D(n72[4]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[4])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i4.GSR = "DISABLED";
    FD1P3IX cycle_counter__i3 (.D(n72[3]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i3.GSR = "DISABLED";
    FD1P3IX cycle_counter__i2 (.D(n72[2]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i2.GSR = "DISABLED";
    FD1P3IX cycle_counter__i1 (.D(n72[1]), .SP(clk_c_enable_269), .CD(n6162), 
            .CK(clk_c), .Q(cycle_counter[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i1.GSR = "DISABLED";
    FD1P3IX fsm_state__i3 (.D(n31502), .SP(next_bit), .CD(n32684), .CK(clk_c), 
            .Q(fsm_state[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i3.GSR = "DISABLED";
    FD1P3IX fsm_state__i0 (.D(n32865), .SP(clk_c_enable_271), .CD(n17837), 
            .CK(clk_c), .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i0.GSR = "DISABLED";
    FD1P3IX fsm_state__i2 (.D(n31493), .SP(next_bit), .CD(n32684), .CK(clk_c), 
            .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1P3IX fsm_state__i1 (.D(n162[1]), .SP(next_bit), .CD(n32684), .CK(clk_c), 
            .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i1.GSR = "DISABLED";
    LUT4 i15474_3_lut_3_lut_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(fsm_state[0]), .Z(n162[1])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(72[17:37])
    defparam i15474_3_lut_3_lut_4_lut.init = 16'h33c4;
    FD1S3JX txd_reg_46 (.D(uart_txd_N_3003), .CK(clk_c), .PD(clk_c_enable_432), 
            .Q(\uo_out_from_user_peri[2][6] )) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(123[8] 133[4])
    defparam txd_reg_46.GSR = "DISABLED";
    LUT4 mux_13_i1_3_lut_4_lut (.A(n32730), .B(n32666), .C(\data_to_write[0] ), 
         .D(data_to_send[1]), .Z(data_to_send_7__N_2975[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_13_i1_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_13_i7_3_lut_4_lut (.A(n32730), .B(n32666), .C(\data_to_write[6] ), 
         .D(data_to_send[7]), .Z(data_to_send_7__N_2975[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_13_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_13_i6_3_lut_4_lut (.A(n32730), .B(n32666), .C(\data_to_write[5] ), 
         .D(data_to_send[6]), .Z(data_to_send_7__N_2975[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_13_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_13_i5_3_lut_4_lut (.A(n32730), .B(n32666), .C(\data_to_write[4] ), 
         .D(data_to_send[5]), .Z(data_to_send_7__N_2975[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_13_i5_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_13_i4_3_lut_4_lut (.A(n32730), .B(n32666), .C(\data_to_write[3] ), 
         .D(data_to_send[4]), .Z(data_to_send_7__N_2975[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_13_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_13_i3_3_lut_4_lut (.A(n32730), .B(n32666), .C(\data_to_write[2] ), 
         .D(data_to_send[3]), .Z(data_to_send_7__N_2975[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_13_i3_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_13_i2_3_lut_4_lut (.A(n32730), .B(n32666), .C(\data_to_write[1] ), 
         .D(data_to_send[2]), .Z(data_to_send_7__N_2975[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_13_i2_3_lut_4_lut.init = 16'hfe10;
    FD1P3IX data_to_send__i0 (.D(data_to_send_7__N_2975[0]), .SP(clk_c_enable_515), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i0.GSR = "DISABLED";
    FD1P3IX data_to_send__i6 (.D(data_to_send_7__N_2975[6]), .SP(clk_c_enable_515), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[6])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i6.GSR = "DISABLED";
    FD1P3IX data_to_send__i5 (.D(data_to_send_7__N_2975[5]), .SP(clk_c_enable_515), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[5])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i5.GSR = "DISABLED";
    FD1P3IX data_to_send__i4 (.D(data_to_send_7__N_2975[4]), .SP(clk_c_enable_515), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[4])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i4.GSR = "DISABLED";
    LUT4 fsm_state_0__bdd_4_lut (.A(fsm_state[0]), .B(fsm_state[2]), .C(fsm_state[1]), 
         .D(fsm_state[3]), .Z(n32865)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;
    defparam fsm_state_0__bdd_4_lut.init = 16'h4555;
    FD1P3IX data_to_send__i3 (.D(data_to_send_7__N_2975[3]), .SP(clk_c_enable_515), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i3.GSR = "DISABLED";
    FD1P3IX data_to_send__i2 (.D(data_to_send_7__N_2975[2]), .SP(clk_c_enable_515), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i2.GSR = "DISABLED";
    FD1P3IX data_to_send__i1 (.D(data_to_send_7__N_2975[1]), .SP(clk_c_enable_515), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i1.GSR = "DISABLED";
    FD1P3AX data_to_send__i7 (.D(n26872), .SP(clk_c_enable_515), .CK(clk_c), 
            .Q(data_to_send[7])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i7.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(\gpio_out_func_sel[0][0] ), .B(\gpio_out_func_sel[0][4] ), 
         .C(\uo_out_from_user_peri[2][6] ), .Z(n27757)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(123[8] 133[4])
    defparam i2_3_lut.init = 16'h1010;
    LUT4 fsm_state_1__bdd_3_lut (.A(fsm_state[1]), .B(fsm_state[3]), .C(fsm_state[2]), 
         .Z(uart_txd_N_3005)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;
    defparam fsm_state_1__bdd_3_lut.init = 16'h3636;
    LUT4 fsm_state_3__bdd_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(fsm_state[0]), .Z(n31502)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B (C (D))))) */ ;
    defparam fsm_state_3__bdd_4_lut.init = 16'h6aa2;
    LUT4 fsm_state_2__bdd_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(fsm_state[0]), 
         .Z(n31493)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam fsm_state_2__bdd_3_lut.init = 16'h6a6a;
    LUT4 i15248_4_lut (.A(data_to_send[0]), .B(fsm_state[0]), .C(uart_txd_N_3005), 
         .D(n32763), .Z(uart_txd_N_3003)) /* synthesis lut_function=(A ((D)+!B)+!A !(B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(128[14] 132[8])
    defparam i15248_4_lut.init = 16'haf23;
    LUT4 uart_tx_busy_bdd_3_lut_4_lut (.A(fsm_state[0]), .B(n32763), .C(\addr[2] ), 
         .D(\uart_rx_buf_data[0] ), .Z(n32251)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam uart_tx_busy_bdd_3_lut_4_lut.init = 16'hefe0;
    LUT4 i28568_2_lut_3_lut_4_lut (.A(fsm_state[0]), .B(n32763), .C(next_bit), 
         .D(rst_reg_n), .Z(clk_c_enable_271)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i28568_2_lut_3_lut_4_lut.init = 16'hf1ff;
    
endmodule
//
// Verilog Description of module tqvp_uart_rx
//

module tqvp_uart_rx (GND_net, VCC_net, cycle_counter, \baud_divider[8] , 
            \baud_divider[7] , \baud_divider[6] , \baud_divider[5] , mid_bit, 
            \baud_divider[4] , \baud_divider[3] , \baud_divider[2] , \baud_divider[1] , 
            \baud_divider[12] , \baud_divider[11] , \baud_divider[10] , 
            \baud_divider[9] , \next_fsm_state_3__N_3046[3] , fsm_state, 
            next_bit, n32803, clk_c, clk_c_enable_432, uart_rx_data, 
            \uo_out_from_user_peri[2][7] , rst_reg_n, debug_stop_txn, 
            instr_active_N_2106, next_bit_adj_25, n32763, \fsm_state[0]_adj_26 , 
            clk_c_enable_269, stop_txn_reg, n32755, stop_txn_now_N_2363, 
            clk_c_enable_208, n6162, n32714, qspi_write_done, n10672, 
            spi_clk_pos, n28259, next_bit_adj_27, n32622, uart_txd_N_3005, 
            clk_c_enable_495, n32832, \fsm_state[0]_adj_28 , clk_c_enable_143, 
            \data_to_write[1] , n9031, n762, clk_c_enable_519, n8177, 
            n32524, n29357, n46, n32728, clk_c_enable_286, instr_complete_N_1647, 
            n28957, n32706, clk_c_enable_6, \data_to_write[0] , n8876, 
            n32771, n27178, n29549, clk_c_enable_282, n32636, uart_txd_N_3005_adj_29, 
            clk_c_enable_515, n6142, n28319, n32681, n27931, n1072, 
            clk_c_enable_543, qv_data_read_n, qv_data_write_n, n26691, 
            \qspi_data_in[1] , \qspi_data_out_3__N_5[1] , n26692, \next_fsm_state_3__N_3042[1] ) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input VCC_net;
    output [12:0]cycle_counter;
    input \baud_divider[8] ;
    input \baud_divider[7] ;
    input \baud_divider[6] ;
    input \baud_divider[5] ;
    output mid_bit;
    input \baud_divider[4] ;
    input \baud_divider[3] ;
    input \baud_divider[2] ;
    input \baud_divider[1] ;
    input \baud_divider[12] ;
    input \baud_divider[11] ;
    input \baud_divider[10] ;
    input \baud_divider[9] ;
    input \next_fsm_state_3__N_3046[3] ;
    output [3:0]fsm_state;
    input next_bit;
    input n32803;
    input clk_c;
    output clk_c_enable_432;
    output [7:0]uart_rx_data;
    output \uo_out_from_user_peri[2][7] ;
    input rst_reg_n;
    input debug_stop_txn;
    output instr_active_N_2106;
    input next_bit_adj_25;
    input n32763;
    input \fsm_state[0]_adj_26 ;
    output clk_c_enable_269;
    input stop_txn_reg;
    input n32755;
    input stop_txn_now_N_2363;
    output clk_c_enable_208;
    output n6162;
    input n32714;
    input qspi_write_done;
    output n10672;
    input spi_clk_pos;
    output n28259;
    input next_bit_adj_27;
    input n32622;
    input uart_txd_N_3005;
    output clk_c_enable_495;
    input n32832;
    input \fsm_state[0]_adj_28 ;
    output clk_c_enable_143;
    input \data_to_write[1] ;
    output n9031;
    input n762;
    output clk_c_enable_519;
    output n8177;
    output n32524;
    input n29357;
    input n46;
    input n32728;
    output clk_c_enable_286;
    input instr_complete_N_1647;
    input n28957;
    input n32706;
    output clk_c_enable_6;
    input \data_to_write[0] ;
    output n8876;
    input n32771;
    input n27178;
    input n29549;
    output clk_c_enable_282;
    input n32636;
    input uart_txd_N_3005_adj_29;
    output clk_c_enable_515;
    output n6142;
    input n28319;
    input n32681;
    output n27931;
    input n1072;
    output clk_c_enable_543;
    input [1:0]qv_data_read_n;
    input [1:0]qv_data_write_n;
    output n26691;
    input \qspi_data_in[1] ;
    output \qspi_data_out_3__N_5[1] ;
    output n26692;
    input \next_fsm_state_3__N_3042[1] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n24131, n24132, n24133, n24134, n24233;
    wire [12:0]n57;
    
    wire n32799;
    wire [2:0]n5273;
    wire [2:0]n5255;
    
    wire n32879, n32878, n24228, bit_sample, clk_c_enable_106, n24232, 
        n1105, uart_rx_data_7__N_3090, n24231;
    wire [3:0]next_fsm_state;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(71[11:25])
    
    wire uart_rts_N_3110, n30077, n9, n24230, n24229, n32572, n9529;
    wire [31:0]next_fsm_state_3__N_3058;
    
    CCU2C cycle_counter_12__I_0_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n24131));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(67[21:55])
    defparam cycle_counter_12__I_0_0.INIT0 = 16'h000F;
    defparam cycle_counter_12__I_0_0.INIT1 = 16'h5555;
    defparam cycle_counter_12__I_0_0.INJECT1_0 = "NO";
    defparam cycle_counter_12__I_0_0.INJECT1_1 = "YES";
    CCU2C cycle_counter_12__I_0_11 (.A0(\baud_divider[8] ), .B0(cycle_counter[7]), 
          .C0(\baud_divider[7] ), .D0(cycle_counter[6]), .A1(\baud_divider[6] ), 
          .B1(cycle_counter[5]), .C1(\baud_divider[5] ), .D1(cycle_counter[4]), 
          .CIN(n24132), .COUT(n24133));
    defparam cycle_counter_12__I_0_11.INIT0 = 16'h9009;
    defparam cycle_counter_12__I_0_11.INIT1 = 16'h9009;
    defparam cycle_counter_12__I_0_11.INJECT1_0 = "YES";
    defparam cycle_counter_12__I_0_11.INJECT1_1 = "YES";
    CCU2C cycle_counter_12__I_0_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24134), .S0(mid_bit));
    defparam cycle_counter_12__I_0_13.INIT0 = 16'h0000;
    defparam cycle_counter_12__I_0_13.INIT1 = 16'h0000;
    defparam cycle_counter_12__I_0_13.INJECT1_0 = "NO";
    defparam cycle_counter_12__I_0_13.INJECT1_1 = "NO";
    CCU2C cycle_counter_12__I_0_13_21660 (.A0(\baud_divider[4] ), .B0(cycle_counter[3]), 
          .C0(\baud_divider[3] ), .D0(cycle_counter[2]), .A1(\baud_divider[2] ), 
          .B1(cycle_counter[1]), .C1(\baud_divider[1] ), .D1(cycle_counter[0]), 
          .CIN(n24133), .COUT(n24134));
    defparam cycle_counter_12__I_0_13_21660.INIT0 = 16'h9009;
    defparam cycle_counter_12__I_0_13_21660.INIT1 = 16'h9009;
    defparam cycle_counter_12__I_0_13_21660.INJECT1_0 = "YES";
    defparam cycle_counter_12__I_0_13_21660.INJECT1_1 = "YES";
    CCU2C cycle_counter_12__I_0_9 (.A0(\baud_divider[12] ), .B0(cycle_counter[11]), 
          .C0(\baud_divider[11] ), .D0(cycle_counter[10]), .A1(\baud_divider[10] ), 
          .B1(cycle_counter[9]), .C1(\baud_divider[9] ), .D1(cycle_counter[8]), 
          .CIN(n24131), .COUT(n24132));
    defparam cycle_counter_12__I_0_9.INIT0 = 16'h9009;
    defparam cycle_counter_12__I_0_9.INIT1 = 16'h9009;
    defparam cycle_counter_12__I_0_9.INJECT1_0 = "YES";
    defparam cycle_counter_12__I_0_9.INJECT1_1 = "YES";
    CCU2C cycle_counter_3546_add_4_13 (.A0(cycle_counter[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24233), .S0(n57[11]), .S1(n57[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546_add_4_13.INIT0 = 16'haaa0;
    defparam cycle_counter_3546_add_4_13.INIT1 = 16'haaa0;
    defparam cycle_counter_3546_add_4_13.INJECT1_0 = "NO";
    defparam cycle_counter_3546_add_4_13.INJECT1_1 = "NO";
    LUT4 mux_3161_i1_4_lut (.A(\next_fsm_state_3__N_3046[3] ), .B(fsm_state[0]), 
         .C(n32799), .D(next_bit), .Z(n5273[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A !(B (C+(D))+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3161_i1_4_lut.init = 16'ha3ac;
    LUT4 mux_3159_i1_3_lut (.A(n32803), .B(mid_bit), .C(fsm_state[1]), 
         .Z(n5255[0])) /* synthesis lut_function=(A (B (C))+!A !(C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3159_i1_3_lut.init = 16'h8585;
    LUT4 mux_3020_i4_4_lut_then_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), 
         .C(next_bit), .D(fsm_state[0]), .Z(n32879)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3020_i4_4_lut_then_4_lut.init = 16'h6aaa;
    LUT4 mux_3020_i4_4_lut_else_4_lut (.A(fsm_state[3]), .B(n5273[1]), .C(fsm_state[1]), 
         .D(fsm_state[0]), .Z(n32878)) /* synthesis lut_function=(A (B+!(C))+!A !((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3020_i4_4_lut_else_4_lut.init = 16'h8a8e;
    CCU2C cycle_counter_3546_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycle_counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n24228), .S1(n57[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546_add_4_1.INIT0 = 16'h0000;
    defparam cycle_counter_3546_add_4_1.INIT1 = 16'h555f;
    defparam cycle_counter_3546_add_4_1.INJECT1_0 = "NO";
    defparam cycle_counter_3546_add_4_1.INJECT1_1 = "NO";
    FD1P3IX bit_sample_47 (.D(n32803), .SP(clk_c_enable_106), .CD(clk_c_enable_432), 
            .CK(clk_c), .Q(bit_sample)) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(112[8] 118[4])
    defparam bit_sample_47.GSR = "DISABLED";
    CCU2C cycle_counter_3546_add_4_11 (.A0(cycle_counter[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24232), .COUT(n24233), .S0(n57[9]), 
          .S1(n57[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546_add_4_11.INIT0 = 16'haaa0;
    defparam cycle_counter_3546_add_4_11.INIT1 = 16'haaa0;
    defparam cycle_counter_3546_add_4_11.INJECT1_0 = "NO";
    defparam cycle_counter_3546_add_4_11.INJECT1_1 = "NO";
    FD1S3IX cycle_counter_3546__i0 (.D(n57[0]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i0.GSR = "DISABLED";
    LUT4 next_bit_bdd_4_lut (.A(next_bit), .B(fsm_state[1]), .C(fsm_state[3]), 
         .D(fsm_state[2]), .Z(uart_rx_data_7__N_3090)) /* synthesis lut_function=(!((B (C)+!B (C (D)+!C !(D)))+!A)) */ ;
    defparam next_bit_bdd_4_lut.init = 16'h0a28;
    CCU2C cycle_counter_3546_add_4_9 (.A0(cycle_counter[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24231), .COUT(n24232), .S0(n57[7]), 
          .S1(n57[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546_add_4_9.INIT0 = 16'haaa0;
    defparam cycle_counter_3546_add_4_9.INIT1 = 16'haaa0;
    defparam cycle_counter_3546_add_4_9.INJECT1_0 = "NO";
    defparam cycle_counter_3546_add_4_9.INJECT1_1 = "NO";
    FD1P3AX recieved_data_i0_i0 (.D(uart_rx_data[1]), .SP(uart_rx_data_7__N_3090), 
            .CK(clk_c), .Q(uart_rx_data[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i0.GSR = "DISABLED";
    FD1S3IX fsm_state__i0 (.D(next_fsm_state[0]), .CK(clk_c), .CD(clk_c_enable_432), 
            .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(136[8] 142[4])
    defparam fsm_state__i0.GSR = "DISABLED";
    FD1S3JX uart_rts_50 (.D(uart_rts_N_3110), .CK(clk_c), .PD(clk_c_enable_432), 
            .Q(\uo_out_from_user_peri[2][7] )) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(145[8] 152[4])
    defparam uart_rts_50.GSR = "DISABLED";
    LUT4 i1_4_lut_rep_784 (.A(fsm_state[2]), .B(fsm_state[0]), .C(fsm_state[1]), 
         .D(fsm_state[3]), .Z(n32799)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_rep_784.init = 16'h5001;
    LUT4 i28593_2_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(fsm_state[1]), 
         .D(fsm_state[3]), .Z(n30077)) /* synthesis lut_function=(A+(B+!(C (D)+!C !(D)))) */ ;
    defparam i28593_2_lut_4_lut.init = 16'heffe;
    LUT4 uart_rts_I_274_2_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[1]), 
         .C(fsm_state[3]), .D(\next_fsm_state_3__N_3046[3] ), .Z(uart_rts_N_3110)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam uart_rts_I_274_2_lut_4_lut.init = 16'hfe00;
    LUT4 i22_4_lut_3_lut (.A(fsm_state[1]), .B(fsm_state[3]), .C(fsm_state[0]), 
         .Z(n9)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;
    defparam i22_4_lut_3_lut.init = 16'h8181;
    CCU2C cycle_counter_3546_add_4_7 (.A0(cycle_counter[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24230), .COUT(n24231), .S0(n57[5]), 
          .S1(n57[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546_add_4_7.INIT0 = 16'haaa0;
    defparam cycle_counter_3546_add_4_7.INIT1 = 16'haaa0;
    defparam cycle_counter_3546_add_4_7.INJECT1_0 = "NO";
    defparam cycle_counter_3546_add_4_7.INJECT1_1 = "NO";
    CCU2C cycle_counter_3546_add_4_5 (.A0(cycle_counter[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24229), .COUT(n24230), .S0(n57[3]), 
          .S1(n57[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546_add_4_5.INIT0 = 16'haaa0;
    defparam cycle_counter_3546_add_4_5.INIT1 = 16'haaa0;
    defparam cycle_counter_3546_add_4_5.INJECT1_0 = "NO";
    defparam cycle_counter_3546_add_4_5.INJECT1_1 = "NO";
    FD1S3IX cycle_counter_3546__i1 (.D(n57[1]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i1.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i2 (.D(n57[2]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i2.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i3 (.D(n57[3]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i3.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i4 (.D(n57[4]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i4.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i5 (.D(n57[5]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i5.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i6 (.D(n57[6]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i6.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i7 (.D(n57[7]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i7.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i8 (.D(n57[8]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i8.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i9 (.D(n57[9]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i9.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i10 (.D(n57[10]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i10.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i11 (.D(n57[11]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i11.GSR = "DISABLED";
    FD1S3IX cycle_counter_3546__i12 (.D(n57[12]), .CK(clk_c), .CD(n1105), 
            .Q(cycle_counter[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546__i12.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i1 (.D(uart_rx_data[2]), .SP(uart_rx_data_7__N_3090), 
            .CK(clk_c), .Q(uart_rx_data[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i1.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i2 (.D(uart_rx_data[3]), .SP(uart_rx_data_7__N_3090), 
            .CK(clk_c), .Q(uart_rx_data[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i2.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i3 (.D(uart_rx_data[4]), .SP(uart_rx_data_7__N_3090), 
            .CK(clk_c), .Q(uart_rx_data[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i3.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i4 (.D(uart_rx_data[5]), .SP(uart_rx_data_7__N_3090), 
            .CK(clk_c), .Q(uart_rx_data[4])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i4.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i5 (.D(uart_rx_data[6]), .SP(uart_rx_data_7__N_3090), 
            .CK(clk_c), .Q(uart_rx_data[5])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i5.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i6 (.D(uart_rx_data[7]), .SP(uart_rx_data_7__N_3090), 
            .CK(clk_c), .Q(uart_rx_data[6])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i6.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i7 (.D(bit_sample), .SP(uart_rx_data_7__N_3090), 
            .CK(clk_c), .Q(uart_rx_data[7])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i7.GSR = "DISABLED";
    FD1S3IX fsm_state__i1 (.D(next_fsm_state[1]), .CK(clk_c), .CD(clk_c_enable_432), 
            .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(136[8] 142[4])
    defparam fsm_state__i1.GSR = "DISABLED";
    LUT4 i4650_2_lut_rep_557 (.A(fsm_state[0]), .B(next_bit), .Z(n32572)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(93[33:48])
    defparam i4650_2_lut_rep_557.init = 16'h8888;
    FD1S3IX fsm_state__i2 (.D(next_fsm_state_3__N_3058[2]), .CK(clk_c), 
            .CD(n9529), .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(136[8] 142[4])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1S3IX fsm_state__i3 (.D(next_fsm_state[3]), .CK(clk_c), .CD(clk_c_enable_432), 
            .Q(fsm_state[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(136[8] 142[4])
    defparam fsm_state__i3.GSR = "DISABLED";
    LUT4 i4663_2_lut_3_lut_4_lut (.A(fsm_state[0]), .B(next_bit), .C(fsm_state[2]), 
         .D(fsm_state[1]), .Z(next_fsm_state_3__N_3058[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(93[33:48])
    defparam i4663_2_lut_3_lut_4_lut.init = 16'h78f0;
    CCU2C cycle_counter_3546_add_4_3 (.A0(cycle_counter[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n24228), .COUT(n24229), .S0(n57[1]), 
          .S1(n57[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3546_add_4_3.INIT0 = 16'haaa0;
    defparam cycle_counter_3546_add_4_3.INIT1 = 16'haaa0;
    defparam cycle_counter_3546_add_4_3.INJECT1_0 = "NO";
    defparam cycle_counter_3546_add_4_3.INJECT1_1 = "NO";
    LUT4 rst_reg_n_I_0_1_lut_rep_829 (.A(rst_reg_n), .Z(clk_c_enable_432)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam rst_reg_n_I_0_1_lut_rep_829.init = 16'h5555;
    LUT4 rstn_N_2029_I_0_2_lut_2_lut (.A(rst_reg_n), .B(debug_stop_txn), 
         .Z(instr_active_N_2106)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam rstn_N_2029_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(next_bit_adj_25), .C(n32763), 
         .D(\fsm_state[0]_adj_26 ), .Z(clk_c_enable_269)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut (.A(rst_reg_n), .B(stop_txn_reg), .C(n32755), 
         .D(stop_txn_now_N_2363), .Z(clk_c_enable_208)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut.init = 16'hfffd;
    LUT4 i735_2_lut_2_lut (.A(rst_reg_n), .B(next_bit_adj_25), .Z(n6162)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i735_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(n32714), .C(qspi_write_done), 
         .D(n32755), .Z(n10672)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 i1_3_lut_3_lut (.A(rst_reg_n), .B(stop_txn_reg), .C(spi_clk_pos), 
         .Z(n28259)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i1_4_lut_4_lut_adj_601 (.A(rst_reg_n), .B(next_bit_adj_27), .C(n32622), 
         .D(uart_txd_N_3005), .Z(clk_c_enable_495)) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_601.init = 16'hfdf5;
    LUT4 i1_3_lut_4_lut_4_lut_adj_602 (.A(rst_reg_n), .B(next_bit_adj_27), 
         .C(n32832), .D(\fsm_state[0]_adj_28 ), .Z(clk_c_enable_143)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_602.init = 16'hfffd;
    LUT4 i14935_2_lut_2_lut (.A(rst_reg_n), .B(\data_to_write[1] ), .Z(n9031)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i14935_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_2_lut (.A(rst_reg_n), .B(n762), .Z(clk_c_enable_519)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_603 (.A(rst_reg_n), .B(stop_txn_now_N_2363), 
         .C(n32755), .D(stop_txn_reg), .Z(n8177)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_603.init = 16'hffdf;
    LUT4 i1_4_lut_4_lut_adj_604 (.A(rst_reg_n), .B(n9), .C(next_bit), 
         .D(fsm_state[2]), .Z(n1105)) /* synthesis lut_function=((B (C+!(D))+!B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_604.init = 16'hf5fd;
    LUT4 i1_2_lut_rep_509_3_lut_3_lut (.A(rst_reg_n), .B(stop_txn_now_N_2363), 
         .C(stop_txn_reg), .Z(n32524)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_2_lut_rep_509_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i1_4_lut_4_lut_adj_605 (.A(rst_reg_n), .B(n29357), .C(n46), .D(n32728), 
         .Z(clk_c_enable_286)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_605.init = 16'h55d5;
    LUT4 i1_4_lut_4_lut_adj_606 (.A(rst_reg_n), .B(instr_complete_N_1647), 
         .C(n28957), .D(n32706), .Z(clk_c_enable_6)) /* synthesis lut_function=((B (C+(D))+!B (D))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_606.init = 16'hffd5;
    LUT4 i15001_2_lut_2_lut (.A(rst_reg_n), .B(\data_to_write[0] ), .Z(n8876)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i15001_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut_adj_607 (.A(rst_reg_n), .B(n32771), .C(n27178), 
         .D(n29549), .Z(clk_c_enable_282)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_607.init = 16'h5d55;
    LUT4 i1_4_lut_4_lut_adj_608 (.A(rst_reg_n), .B(next_bit_adj_25), .C(n32636), 
         .D(uart_txd_N_3005_adj_29), .Z(clk_c_enable_515)) /* synthesis lut_function=((B ((D)+!C)+!B !(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_608.init = 16'hdf5f;
    LUT4 i444_2_lut_2_lut (.A(rst_reg_n), .B(next_bit_adj_27), .Z(n6142)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i444_2_lut_2_lut.init = 16'hdddd;
    LUT4 i3868_2_lut_2_lut (.A(rst_reg_n), .B(mid_bit), .Z(clk_c_enable_106)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i3868_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut_adj_609 (.A(rst_reg_n), .B(n28319), .C(stop_txn_now_N_2363), 
         .D(n32681), .Z(n27931)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_609.init = 16'hfffd;
    LUT4 i6847_2_lut_2_lut (.A(rst_reg_n), .B(n32799), .Z(n9529)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i6847_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_610 (.A(rst_reg_n), .B(stop_txn_now_N_2363), 
         .C(n1072), .D(stop_txn_reg), .Z(clk_c_enable_543)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_610.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_611 (.A(rst_reg_n), .B(qv_data_read_n[1]), .C(qv_data_write_n[1]), 
         .D(n32771), .Z(n26691)) /* synthesis lut_function=((B (C+(D))+!B (D))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_611.init = 16'hffd5;
    LUT4 i15175_2_lut_2_lut (.A(rst_reg_n), .B(\qspi_data_in[1] ), .Z(\qspi_data_out_3__N_5[1] )) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i15175_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut (.A(qv_data_write_n[0]), .B(n26691), .C(qv_data_read_n[0]), 
         .Z(n26692)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 mux_3020_i2_4_lut (.A(fsm_state[1]), .B(n5273[1]), .C(n32799), 
         .D(n32572), .Z(next_fsm_state[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3020_i2_4_lut.init = 16'hc5ca;
    LUT4 mux_3161_i2_4_lut (.A(\next_fsm_state_3__N_3042[1] ), .B(\next_fsm_state_3__N_3046[3] ), 
         .C(fsm_state[0]), .D(fsm_state[1]), .Z(n5273[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3161_i2_4_lut.init = 16'hcac0;
    PFUMX i29318 (.BLUT(n32878), .ALUT(n32879), .C0(fsm_state[2]), .Z(next_fsm_state[3]));
    PFUMX mux_3020_i1 (.BLUT(n5255[0]), .ALUT(n5273[0]), .C0(n30077), 
          .Z(next_fsm_state[0]));
    
endmodule
//
// Verilog Description of module tqvp_led_byte
//

module tqvp_led_byte (led_state, clk_c, clk_c_enable_282, clk_c_enable_432, 
            \data_to_write[0] ) /* synthesis syn_module_defined=1 */ ;
    output led_state;
    input clk_c;
    input clk_c_enable_282;
    input clk_c_enable_432;
    input \data_to_write[0] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    FD1P3IX led_state_15 (.D(\data_to_write[0] ), .SP(clk_c_enable_282), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(led_state)) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=16, LSE_RCOL=3, LSE_LLINE=250, LSE_RLINE=264 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/led.v(22[12] 28[8])
    defparam led_state_15.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module tinyQV
//

module tinyQV (rst_reg_n_adj_17, clk_c, rst_reg_n, n32771, instr_active_N_2106, 
            n26692, qspi_write_done, \instr_addr_23__N_318[7] , \instr_addr_23__N_318[6] , 
            \addr[7] , \instr_addr_23__N_318[8] , \instr_addr_23__N_318[20] , 
            \instr_addr_23__N_318[21] , \instr_addr_23__N_318[2] , \addr[3] , 
            \addr[2] , \instr_addr[1] , \addr[1] , n32522, n32755, 
            clk_c_enable_432, n26691, n10672, data_stall, n29887, 
            n32523, data_to_write, is_writing_N_2331, \data_to_write[12] , 
            \data_to_write[11] , \data_to_write[10] , \data_to_write[9] , 
            \data_to_write[8] , \data_to_write[7] , \data_to_write[6] , 
            \data_to_write[5] , \data_to_write[4] , \data_to_write[2] , 
            \addr[0] , n32714, continue_txn_N_2131, data_stall_N_2158, 
            n32801, \instr_addr_23__N_318[5] , \addr[6] , \instr_addr_23__N_318[11] , 
            \instr_addr_23__N_318[14] , \instr_addr_23__N_318[9] , \addr[10] , 
            \instr_addr_23__N_318[15] , \instr_addr_23__N_318[16] , \instr_addr_23__N_318[17] , 
            \instr_addr_23__N_318[12] , \instr_addr_23__N_318[10] , \instr_addr_23__N_318[13] , 
            \instr_addr_23__N_318[3] , \addr[4] , is_writing, spi_clk_pos, 
            stop_txn_now_N_2363, \instr_addr_23__N_318[22] , \instr_addr_23__N_318[4] , 
            \addr[5] , \instr_addr_23__N_318[19] , \instr_addr_23__N_318[18] , 
            fsm_state, clk_c_enable_340, n32524, clk_c_enable_208, clk_c_enable_66, 
            n29884, n27931, n32681, n8177, qspi_data_out_3__N_5, \qspi_data_in[3] , 
            \qspi_data_in[2] , qspi_ram_a_select, qspi_ram_b_select, clk_N_45, 
            stop_txn_reg, n32521, \qspi_data_oe[1] , clk_c_enable_341, 
            n1072, debug_stop_txn, \writing_N_164[3] , n4513, n4501, 
            n32833, n26811, n4503, \addr[20] , \addr[22] , n6218, 
            spi_clk_pos_derived_59, qspi_clk_N_56, n6220, clk_c_enable_543, 
            n28319, n32874, n28259, \qspi_data_in[0] , n32060, n28111, 
            n32892, \imm[17] , \instr[31] , \imm[16] , \imm[15] , 
            \imm[14] , \imm[13] , \imm[12] , \imm[11] , \imm[10] , 
            \imm[9] , \imm[8] , \imm[7] , \imm[6] , \imm[5] , \imm[4] , 
            \imm[3] , \imm[2] , \imm[1] , was_early_branch, \rd[0] , 
            qv_data_read_n, n29738, \instr_data[3][0] , \instr_addr_23__N_318[0] , 
            n32656, n26116, debug_instr_valid, n32851, n32835, n32723, 
            \gpio_out_func_sel[5][2] , \gpio_out_func_sel[7][2] , \instr_len[2] , 
            \pc[2] , \pc[1] , n2196, n32727, n2191, n32640, n32548, 
            n32734, n32836, n27888, \gpio_out_func_sel[5][4] , \gpio_out_func_sel[7][4] , 
            n29831, n32655, n32544, \instr_write_offset[3] , n2150, 
            n2130, n4251, n32685, n19, n32660, \peri_data_out[11] , 
            n4, \peri_data_out[10] , n32642, \peri_data_out[9] , n31796, 
            n31795, n32520, n32654, \pc[7] , \pc[15] , n32842, \next_pc_for_core[6] , 
            \pc[3] , \pc[11] , n32251, n31706, clk_c_enable_285, n28957, 
            n34285, \pc[6] , \pc[14] , \pc[10] , n3, n3_adj_18, 
            n32638, n29707, qv_data_write_n, \addr[27] , n32850, \imm[21] , 
            \imm[20] , \next_pc_for_core[9] , \next_pc_for_core[13] , 
            \pc[5] , \pc[13] , \pc[9] , \next_pc_for_core[4] , n12, 
            data_ready_r_N_2823, data_ready_r, n32706, n15569, \data_to_write[3] , 
            \data_to_write[1] , n2211, n17165, VCC_net, n32694, n7, 
            n8854, \next_pc_for_core[10] , \next_pc_for_core[14] , \instr_data[0][0] , 
            \instr_data[1][7] , \instr_data[1][0] , \instr_data[2][7] , 
            \next_pc_for_core[8] , \next_pc_for_core[12] , \instr_data[2][0] , 
            \instr_data[3][7] , n32552, n8109, n32695, n32728, n32745, 
            \next_pc_for_core[3] , \next_pc_for_core[5] , \next_pc_for_core[7] , 
            \next_pc_for_core[11] , \pc[21] , \pc[17] , \next_pc_for_core[20] , 
            \next_pc_for_core[16] , \pc[23] , \pc[19] , \pc[22] , \pc[18] , 
            \pc[20] , \pc[16] , \next_pc_for_core[15] , \next_pc_for_core[21] , 
            \next_pc_for_core[17] , \imm[23] , \imm[22] , \imm[19] , 
            \imm[18] , \next_pc_for_core[22] , \next_pc_for_core[18] , 
            \next_pc_for_core[19] , n28077, \next_pc_for_core[23] , n32819, 
            n32720, n29357, \uo_out_from_user_peri[1][6] , \data_from_user_peri_1__31__N_2455[2] , 
            \uo_out_from_user_peri[1][2] , \uo_out_from_user_peri[1][5] , 
            n29491, \data_from_read[2] , \early_branch_addr[7] , \early_branch_addr[3] , 
            \early_branch_addr[6] , \early_branch_addr[2] , \early_branch_addr[4] , 
            n32822, \early_branch_addr[8] , \early_branch_addr[5] , \early_branch_addr[9] , 
            \early_branch_addr[10] , \early_branch_addr[11] , \early_branch_addr[12] , 
            \early_branch_addr[13] , \early_branch_addr[14] , \early_branch_addr[15] , 
            \early_branch_addr[17] , \early_branch_addr[18] , \early_branch_addr[19] , 
            \early_branch_addr[20] , \early_branch_addr[21] , \early_branch_addr[22] , 
            \early_branch_addr[23] , \early_branch_addr[16] , n16811, 
            n2594, n31883, \pc_23__N_911[13] , \pc[12] , n26838, n10944, 
            n32725, n32761, n32729, \cycle[0] , \pc[8] , n27178, 
            n32766, \pc[4] , n32737, \data_from_peri_31__N_2415[0] , 
            n32693, clk_c_enable_50, n32818, clk_c_enable_154, clk_c_enable_283, 
            clk_c_enable_354, \gpio_out_func_sel[0][2] , \gpio_out_func_sel[1][2] , 
            \gpio_out_func_sel[2][2] , \gpio_out_func_sel[3][2] , n32756, 
            n5169, n32825, n29127, \gpio_out_func_sel[4][2] , \gpio_out_func_sel[6][2] , 
            \uart_rx_buf_data[4] , \baud_divider[4] , gpio_out_sel, n14, 
            n14_adj_19, n29293, instr_complete_N_1647, \data_from_read[6] , 
            n32672, n46, \connect_peripheral[1] , \connect_peripheral[0] , 
            n32568, n29741, n29, \uart_rx_buf_data[7] , \baud_divider[7] , 
            n2, n32614, \next_fsm_state_3__N_3046[3] , \ui_in_sync[5] , 
            \ui_in_sync[6] , n32072, n29549, \ui_in_sync[7] , \data_from_user_peri_1__31__N_2455[7] , 
            \uart_rx_buf_data[6] , n26856, \baud_divider[6] , \uart_rx_buf_data[5] , 
            \baud_divider[5] , \data_from_read[4] , \data_from_read[8] , 
            \data_from_read[12] , \data_from_read[1] , \data_from_user_peri_1__31__N_2455[0] , 
            \uo_out_from_user_peri[1][0] , \data_from_read[5] , data_out_hold, 
            \data_from_read[3] , \data_from_read[7] , \uart_rx_buf_data[3] , 
            \baud_divider[3] , n2_adj_20, \data_from_read[0] , n32759, 
            \uart_rx_buf_data[2] , \baud_divider[2] , n10737, n32650, 
            \instr[16] , n32615, n32610, clk_c_enable_342, \ui_in_sync[1] , 
            \ui_in_sync[0] , debug_rd, n29866, n17920, accum, d_3__N_1868, 
            fsm_state_adj_24, n32791, n32763, n32730, n32834, n32710, 
            n31351, n1152, \mul_out[3] , \mul_out[2] , \mul_out[1] , 
            \csr_read_3__N_1447[2] , \next_accum[5] , GND_net, \next_accum[16] , 
            \next_accum[17] , \next_accum[18] , \next_accum[19] , \next_accum[6] , 
            \next_accum[7] , \next_accum[8] , \next_accum[9] , \next_accum[10] , 
            \next_accum[11] , \next_accum[12] , \next_accum[13] , \next_accum[14] , 
            \next_accum[15] , \next_accum[4] , \return_addr[16] ) /* synthesis syn_module_defined=1 */ ;
    output rst_reg_n_adj_17;
    input clk_c;
    input rst_reg_n;
    output n32771;
    input instr_active_N_2106;
    input n26692;
    output qspi_write_done;
    input \instr_addr_23__N_318[7] ;
    input \instr_addr_23__N_318[6] ;
    output \addr[7] ;
    input \instr_addr_23__N_318[8] ;
    input \instr_addr_23__N_318[20] ;
    input \instr_addr_23__N_318[21] ;
    input \instr_addr_23__N_318[2] ;
    output \addr[3] ;
    output \addr[2] ;
    input \instr_addr[1] ;
    output \addr[1] ;
    output n32522;
    output n32755;
    input clk_c_enable_432;
    input n26691;
    input n10672;
    output data_stall;
    input n29887;
    output n32523;
    output [31:0]data_to_write;
    output is_writing_N_2331;
    output \data_to_write[12] ;
    output \data_to_write[11] ;
    output \data_to_write[10] ;
    output \data_to_write[9] ;
    output \data_to_write[8] ;
    output \data_to_write[7] ;
    output \data_to_write[6] ;
    output \data_to_write[5] ;
    output \data_to_write[4] ;
    output \data_to_write[2] ;
    output \addr[0] ;
    output n32714;
    output continue_txn_N_2131;
    output data_stall_N_2158;
    output n32801;
    input \instr_addr_23__N_318[5] ;
    output \addr[6] ;
    input \instr_addr_23__N_318[11] ;
    input \instr_addr_23__N_318[14] ;
    input \instr_addr_23__N_318[9] ;
    output \addr[10] ;
    input \instr_addr_23__N_318[15] ;
    input \instr_addr_23__N_318[16] ;
    input \instr_addr_23__N_318[17] ;
    input \instr_addr_23__N_318[12] ;
    input \instr_addr_23__N_318[10] ;
    input \instr_addr_23__N_318[13] ;
    input \instr_addr_23__N_318[3] ;
    output \addr[4] ;
    output is_writing;
    output spi_clk_pos;
    output stop_txn_now_N_2363;
    input \instr_addr_23__N_318[22] ;
    input \instr_addr_23__N_318[4] ;
    output \addr[5] ;
    input \instr_addr_23__N_318[19] ;
    input \instr_addr_23__N_318[18] ;
    output [2:0]fsm_state;
    input clk_c_enable_340;
    input n32524;
    input clk_c_enable_208;
    input clk_c_enable_66;
    input n29884;
    input n27931;
    output n32681;
    input n8177;
    input [3:0]qspi_data_out_3__N_5;
    input \qspi_data_in[3] ;
    input \qspi_data_in[2] ;
    output qspi_ram_a_select;
    output qspi_ram_b_select;
    input clk_N_45;
    output stop_txn_reg;
    output n32521;
    output \qspi_data_oe[1] ;
    input clk_c_enable_341;
    output n1072;
    output debug_stop_txn;
    output \writing_N_164[3] ;
    output n4513;
    output n4501;
    output n32833;
    output n26811;
    output n4503;
    output \addr[20] ;
    output \addr[22] ;
    output n6218;
    output spi_clk_pos_derived_59;
    output qspi_clk_N_56;
    output n6220;
    input clk_c_enable_543;
    output n28319;
    output n32874;
    input n28259;
    input \qspi_data_in[0] ;
    output n32060;
    output n28111;
    output n32892;
    output \imm[17] ;
    output \instr[31] ;
    output \imm[16] ;
    output \imm[15] ;
    output \imm[14] ;
    output \imm[13] ;
    output \imm[12] ;
    output \imm[11] ;
    output \imm[10] ;
    output \imm[9] ;
    output \imm[8] ;
    output \imm[7] ;
    output \imm[6] ;
    output \imm[5] ;
    output \imm[4] ;
    output \imm[3] ;
    output \imm[2] ;
    output \imm[1] ;
    output was_early_branch;
    output \rd[0] ;
    output [1:0]qv_data_read_n;
    input n29738;
    output \instr_data[3][0] ;
    output \instr_addr_23__N_318[0] ;
    output n32656;
    output n26116;
    output debug_instr_valid;
    output n32851;
    output n32835;
    output n32723;
    input \gpio_out_func_sel[5][2] ;
    input \gpio_out_func_sel[7][2] ;
    output \instr_len[2] ;
    output \pc[2] ;
    output \pc[1] ;
    output n2196;
    output n32727;
    output n2191;
    output n32640;
    output n32548;
    output n32734;
    input n32836;
    output n27888;
    input \gpio_out_func_sel[5][4] ;
    input \gpio_out_func_sel[7][4] ;
    output n29831;
    output n32655;
    output n32544;
    output \instr_write_offset[3] ;
    input n2150;
    input n2130;
    output n4251;
    output n32685;
    output n19;
    output n32660;
    input \peri_data_out[11] ;
    output n4;
    input \peri_data_out[10] ;
    output n32642;
    input \peri_data_out[9] ;
    input n31796;
    input n31795;
    output n32520;
    input n32654;
    output \pc[7] ;
    output \pc[15] ;
    output n32842;
    input \next_pc_for_core[6] ;
    output \pc[3] ;
    output \pc[11] ;
    input n32251;
    input n31706;
    output clk_c_enable_285;
    output n28957;
    output n34285;
    output \pc[6] ;
    output \pc[14] ;
    output \pc[10] ;
    output n3;
    output n3_adj_18;
    input n32638;
    input n29707;
    output [1:0]qv_data_write_n;
    output \addr[27] ;
    output n32850;
    output \imm[21] ;
    output \imm[20] ;
    input \next_pc_for_core[9] ;
    input \next_pc_for_core[13] ;
    output \pc[5] ;
    output \pc[13] ;
    output \pc[9] ;
    input \next_pc_for_core[4] ;
    input n12;
    output data_ready_r_N_2823;
    input data_ready_r;
    output n32706;
    output n15569;
    output \data_to_write[3] ;
    output \data_to_write[1] ;
    output n2211;
    input n17165;
    input VCC_net;
    output n32694;
    output n7;
    input n8854;
    input \next_pc_for_core[10] ;
    input \next_pc_for_core[14] ;
    output \instr_data[0][0] ;
    output \instr_data[1][7] ;
    output \instr_data[1][0] ;
    output \instr_data[2][7] ;
    input \next_pc_for_core[8] ;
    input \next_pc_for_core[12] ;
    output \instr_data[2][0] ;
    output \instr_data[3][7] ;
    output n32552;
    output n8109;
    output n32695;
    output n32728;
    output n32745;
    input \next_pc_for_core[3] ;
    input \next_pc_for_core[5] ;
    input \next_pc_for_core[7] ;
    input \next_pc_for_core[11] ;
    output \pc[21] ;
    output \pc[17] ;
    input \next_pc_for_core[20] ;
    input \next_pc_for_core[16] ;
    output \pc[23] ;
    output \pc[19] ;
    output \pc[22] ;
    output \pc[18] ;
    output \pc[20] ;
    output \pc[16] ;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[21] ;
    input \next_pc_for_core[17] ;
    output \imm[23] ;
    output \imm[22] ;
    output \imm[19] ;
    output \imm[18] ;
    input \next_pc_for_core[22] ;
    input \next_pc_for_core[18] ;
    input \next_pc_for_core[19] ;
    output n28077;
    input \next_pc_for_core[23] ;
    output n32819;
    output n32720;
    output n29357;
    input \uo_out_from_user_peri[1][6] ;
    input \data_from_user_peri_1__31__N_2455[2] ;
    input \uo_out_from_user_peri[1][2] ;
    input \uo_out_from_user_peri[1][5] ;
    output n29491;
    input \data_from_read[2] ;
    input \early_branch_addr[7] ;
    input \early_branch_addr[3] ;
    input \early_branch_addr[6] ;
    input \early_branch_addr[2] ;
    input \early_branch_addr[4] ;
    input n32822;
    input \early_branch_addr[8] ;
    input \early_branch_addr[5] ;
    input \early_branch_addr[9] ;
    input \early_branch_addr[10] ;
    input \early_branch_addr[11] ;
    input \early_branch_addr[12] ;
    input \early_branch_addr[13] ;
    input \early_branch_addr[14] ;
    input \early_branch_addr[15] ;
    input \early_branch_addr[17] ;
    input \early_branch_addr[18] ;
    input \early_branch_addr[19] ;
    input \early_branch_addr[20] ;
    input \early_branch_addr[21] ;
    input \early_branch_addr[22] ;
    input \early_branch_addr[23] ;
    input \early_branch_addr[16] ;
    output n16811;
    input n2594;
    output n31883;
    input \pc_23__N_911[13] ;
    output \pc[12] ;
    output n26838;
    input n10944;
    output n32725;
    output n32761;
    output n32729;
    output \cycle[0] ;
    output \pc[8] ;
    output n27178;
    output n32766;
    output \pc[4] ;
    output n32737;
    output \data_from_peri_31__N_2415[0] ;
    output n32693;
    output clk_c_enable_50;
    input n32818;
    output clk_c_enable_154;
    output clk_c_enable_283;
    output clk_c_enable_354;
    input \gpio_out_func_sel[0][2] ;
    input \gpio_out_func_sel[1][2] ;
    input \gpio_out_func_sel[2][2] ;
    input \gpio_out_func_sel[3][2] ;
    input n32756;
    output n5169;
    input n32825;
    input n29127;
    input \gpio_out_func_sel[4][2] ;
    input \gpio_out_func_sel[6][2] ;
    input \uart_rx_buf_data[4] ;
    input \baud_divider[4] ;
    input [7:6]gpio_out_sel;
    output n14;
    output n14_adj_19;
    output n29293;
    output instr_complete_N_1647;
    input \data_from_read[6] ;
    output n32672;
    output n46;
    output \connect_peripheral[1] ;
    output \connect_peripheral[0] ;
    input n32568;
    output n29741;
    input n29;
    input \uart_rx_buf_data[7] ;
    input \baud_divider[7] ;
    output n2;
    input n32614;
    input \next_fsm_state_3__N_3046[3] ;
    input \ui_in_sync[5] ;
    input \ui_in_sync[6] ;
    input n32072;
    output n29549;
    input \ui_in_sync[7] ;
    output \data_from_user_peri_1__31__N_2455[7] ;
    input \uart_rx_buf_data[6] ;
    input n26856;
    input \baud_divider[6] ;
    input \uart_rx_buf_data[5] ;
    input \baud_divider[5] ;
    input \data_from_read[4] ;
    input \data_from_read[8] ;
    input \data_from_read[12] ;
    input \data_from_read[1] ;
    input \data_from_user_peri_1__31__N_2455[0] ;
    input \uo_out_from_user_peri[1][0] ;
    input \data_from_read[5] ;
    input data_out_hold;
    input \data_from_read[3] ;
    input \data_from_read[7] ;
    input \uart_rx_buf_data[3] ;
    input \baud_divider[3] ;
    output n2_adj_20;
    input \data_from_read[0] ;
    output n32759;
    input \uart_rx_buf_data[2] ;
    input \baud_divider[2] ;
    input n10737;
    output n32650;
    input \instr[16] ;
    input n32615;
    input n32610;
    input clk_c_enable_342;
    input \ui_in_sync[1] ;
    input \ui_in_sync[0] ;
    output [3:0]debug_rd;
    input n29866;
    output n17920;
    output [15:0]accum;
    output [19:0]d_3__N_1868;
    input [3:0]fsm_state_adj_24;
    output n32791;
    output n32763;
    output n32730;
    output n32834;
    output n32710;
    input n31351;
    output n1152;
    input \mul_out[3] ;
    input \mul_out[2] ;
    input \mul_out[1] ;
    output \csr_read_3__N_1447[2] ;
    input \next_accum[5] ;
    input GND_net;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[4] ;
    output \return_addr[16] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    
    wire n34287, mem_data_ready, n29059, n18458, debug_data_ready, 
        instr_active, start_instr;
    wire [1:0]qspi_data_byte_idx;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(59[15:33])
    wire [1:0]data_txn_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(49[15:27])
    wire [15:0]instr_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(61[15:25])
    wire [27:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    wire [23:1]instr_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(56[15:25])
    wire [31:0]mem_data_from_read;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(74[15:33])
    wire [31:0]qspi_data_buf;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(58[16:29])
    
    wire clk_c_enable_91;
    wire [31:0]instr_data_7__N_1969;
    
    wire debug_data_continue;
    wire [1:0]n174;
    
    wire instr_fetch_running_N_945, n32537, n11193, qspi_data_ready, 
        n32826, n32712, n32598, instr_fetch_stopped, n32531, debug_stop_txn_N_2142;
    wire [31:0]data_to_write_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(56[17:30])
    
    wire n32545, n8, n28687, n16, n32787, n32711, n32788, n1, 
        n21414, n32689, instr_fetch_running, n29618, n32578;
    wire [2:0]fsm_state_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(82[15:24])
    
    wire n32740;
    wire [1:0]read_cycles_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(105[15:32])
    
    wire n32778, data_req_N_2334, n19867, n32542, data_ready_N_2347, 
        n31866;
    wire [2:0]n329;
    
    wire n32789;
    
    FD1S3AX rst_reg_n_16 (.D(rst_reg_n), .CK(clk_c), .Q(rst_reg_n_adj_17)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=111, LSE_RLINE=150 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(92[10:43])
    defparam rst_reg_n_16.GSR = "DISABLED";
    FD1S3AX rst_reg_n_16_rep_850 (.D(rst_reg_n), .CK(clk_c), .Q(n34287)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=111, LSE_RLINE=150 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(92[10:43])
    defparam rst_reg_n_16_rep_850.GSR = "DISABLED";
    LUT4 data_ready_I_0_4_lut (.A(mem_data_ready), .B(n29059), .C(n32771), 
         .D(n18458), .Z(debug_data_ready)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(77[26:62])
    defparam data_ready_I_0_4_lut.init = 16'hcafa;
    tinyqv_mem_ctrl mem (.instr_active(instr_active), .clk_c(clk_c), .instr_active_N_2106(instr_active_N_2106), 
            .start_instr(start_instr), .qspi_data_byte_idx({qspi_data_byte_idx}), 
            .data_txn_len({data_txn_len}), .n26692(n26692), .qspi_write_done(qspi_write_done), 
            .instr_data({instr_data}), .\instr_addr_23__N_318[7] (\instr_addr_23__N_318[7] ), 
            .\addr[8] (addr[8]), .\instr_addr_23__N_318[6] (\instr_addr_23__N_318[6] ), 
            .\addr[7] (\addr[7] ), .\instr_addr_23__N_318[8] (\instr_addr_23__N_318[8] ), 
            .\addr[9] (addr[9]), .\instr_addr_23__N_318[20] (\instr_addr_23__N_318[20] ), 
            .\addr[21] (addr[21]), .\instr_addr_23__N_318[21] (\instr_addr_23__N_318[21] ), 
            .\addr[22] (addr[22]), .\instr_addr_23__N_318[2] (\instr_addr_23__N_318[2] ), 
            .\addr[3] (\addr[3] ), .\instr_addr[2] (instr_addr[2]), .\addr[2] (\addr[2] ), 
            .\mem_data_from_read[23] (mem_data_from_read[23]), .\mem_data_from_read[22] (mem_data_from_read[22]), 
            .\mem_data_from_read[21] (mem_data_from_read[21]), .\mem_data_from_read[20] (mem_data_from_read[20]), 
            .\mem_data_from_read[19] (mem_data_from_read[19]), .\mem_data_from_read[18] (mem_data_from_read[18]), 
            .\mem_data_from_read[17] (mem_data_from_read[17]), .\mem_data_from_read[16] (mem_data_from_read[16]), 
            .\qspi_data_buf[15] (qspi_data_buf[15]), .clk_c_enable_91(clk_c_enable_91), 
            .\qspi_data_buf[14] (qspi_data_buf[14]), .\qspi_data_buf[13] (qspi_data_buf[13]), 
            .\qspi_data_buf[11] (qspi_data_buf[11]), .\qspi_data_buf[10] (qspi_data_buf[10]), 
            .\qspi_data_buf[9] (qspi_data_buf[9]), .\instr_data_7__N_1969[3] (instr_data_7__N_1969[3]), 
            .\instr_data_7__N_1969[1] (instr_data_7__N_1969[1]), .\instr_addr[1] (\instr_addr[1] ), 
            .\addr[1] (\addr[1] ), .mem_data_ready(mem_data_ready), .\mem_data_from_read[29] (mem_data_from_read[29]), 
            .\mem_data_from_read[25] (mem_data_from_read[25]), .n32522(n32522), 
            .\mem_data_from_read[31] (mem_data_from_read[31]), .\mem_data_from_read[27] (mem_data_from_read[27]), 
            .\mem_data_from_read[28] (mem_data_from_read[28]), .\mem_data_from_read[24] (mem_data_from_read[24]), 
            .\mem_data_from_read[30] (mem_data_from_read[30]), .\mem_data_from_read[26] (mem_data_from_read[26]), 
            .n32755(n32755), .clk_c_enable_432(clk_c_enable_432), .debug_data_continue(debug_data_continue), 
            .n175(n174[1]), .n26691(n26691), .instr_fetch_running_N_945(instr_fetch_running_N_945), 
            .n10672(n10672), .n32537(n32537), .n11193(n11193), .qspi_data_ready(qspi_data_ready), 
            .data_stall(data_stall), .rst_reg_n(rst_reg_n), .n29887(n29887), 
            .n32523(n32523), .n32826(n32826), .n32712(n32712), .\addr[24] (addr[24]), 
            .n32598(n32598), .\mem_data_from_read[0] (mem_data_from_read[0]), 
            .\mem_data_from_read[7] (mem_data_from_read[7]), .\mem_data_from_read[3] (mem_data_from_read[3]), 
            .\data_to_write[0] (data_to_write[0]), .\mem_data_from_read[5] (mem_data_from_read[5]), 
            .\mem_data_from_read[1] (mem_data_from_read[1]), .\mem_data_from_read[4] (mem_data_from_read[4]), 
            .instr_fetch_stopped(instr_fetch_stopped), .n32531(n32531), 
            .is_writing_N_2331(is_writing_N_2331), .\mem_data_from_read[12] (mem_data_from_read[12]), 
            .\mem_data_from_read[8] (mem_data_from_read[8]), .debug_stop_txn_N_2142(debug_stop_txn_N_2142), 
            .\data_to_write[31] (data_to_write_c[31]), .n32545(n32545), 
            .n8(n8), .n28687(n28687), .n16(n16), .\data_to_write[30] (data_to_write_c[30]), 
            .\data_to_write[29] (data_to_write_c[29]), .\data_to_write[28] (data_to_write_c[28]), 
            .\data_to_write[27] (data_to_write_c[27]), .\data_to_write[26] (data_to_write_c[26]), 
            .\data_to_write[25] (data_to_write_c[25]), .\data_to_write[24] (data_to_write_c[24]), 
            .\data_to_write[23] (data_to_write_c[23]), .\data_to_write[22] (data_to_write_c[22]), 
            .\data_to_write[21] (data_to_write_c[21]), .\data_to_write[20] (data_to_write_c[20]), 
            .\data_to_write[19] (data_to_write_c[19]), .\data_to_write[18] (data_to_write_c[18]), 
            .\data_to_write[17] (data_to_write_c[17]), .\data_to_write[16] (data_to_write_c[16]), 
            .\data_to_write[15] (data_to_write_c[15]), .\data_to_write[14] (data_to_write_c[14]), 
            .\data_to_write[13] (data_to_write_c[13]), .\data_to_write[12] (\data_to_write[12] ), 
            .\data_to_write[11] (\data_to_write[11] ), .\data_to_write[10] (\data_to_write[10] ), 
            .n32787(n32787), .\data_to_write[9] (\data_to_write[9] ), .\data_to_write[8] (\data_to_write[8] ), 
            .\data_to_write[7] (\data_to_write[7] ), .\data_to_write[6] (\data_to_write[6] ), 
            .\data_to_write[5] (\data_to_write[5] ), .\data_to_write[4] (\data_to_write[4] ), 
            .\data_to_write[2] (\data_to_write[2] ), .\addr[0] (\addr[0] ), 
            .n32711(n32711), .n32714(n32714), .continue_txn_N_2131(continue_txn_N_2131), 
            .data_stall_N_2158(data_stall_N_2158), .n32788(n32788), .n1(n1), 
            .n32771(n32771), .n32801(n32801), .n21414(n21414), .n32689(n32689), 
            .\addr[23] (addr[23]), .instr_fetch_running(instr_fetch_running), 
            .n29618(n29618), .\instr_addr_23__N_318[5] (\instr_addr_23__N_318[5] ), 
            .\addr[6] (\addr[6] ), .\instr_addr_23__N_318[11] (\instr_addr_23__N_318[11] ), 
            .\addr[12] (addr[12]), .\instr_addr_23__N_318[14] (\instr_addr_23__N_318[14] ), 
            .\addr[15] (addr[15]), .\instr_addr_23__N_318[9] (\instr_addr_23__N_318[9] ), 
            .\addr[10] (\addr[10] ), .\instr_addr_23__N_318[15] (\instr_addr_23__N_318[15] ), 
            .\addr[16] (addr[16]), .\instr_addr_23__N_318[16] (\instr_addr_23__N_318[16] ), 
            .\addr[17] (addr[17]), .\instr_addr_23__N_318[17] (\instr_addr_23__N_318[17] ), 
            .\addr[18] (addr[18]), .\instr_addr_23__N_318[12] (\instr_addr_23__N_318[12] ), 
            .\addr[13] (addr[13]), .n32578(n32578), .\instr_addr_23__N_318[10] (\instr_addr_23__N_318[10] ), 
            .\addr[11] (addr[11]), .\instr_addr_23__N_318[13] (\instr_addr_23__N_318[13] ), 
            .\addr[14] (addr[14]), .\instr_addr_23__N_318[3] (\instr_addr_23__N_318[3] ), 
            .\addr[4] (\addr[4] ), .is_writing(is_writing), .spi_clk_pos(spi_clk_pos), 
            .stop_txn_now_N_2363(stop_txn_now_N_2363), .\instr_addr_23__N_318[22] (\instr_addr_23__N_318[22] ), 
            .\instr_addr_23__N_318[4] (\instr_addr_23__N_318[4] ), .\addr[5] (\addr[5] ), 
            .\instr_addr_23__N_318[19] (\instr_addr_23__N_318[19] ), .\addr[20] (addr[20]), 
            .\instr_addr_23__N_318[18] (\instr_addr_23__N_318[18] ), .\addr[19] (addr[19]), 
            .fsm_state({fsm_state_c[2:1], fsm_state[0]}), .clk_c_enable_340(clk_c_enable_340), 
            .n32524(n32524), .clk_c_enable_208(clk_c_enable_208), .clk_c_enable_66(clk_c_enable_66), 
            .n29884(n29884), .n27931(n27931), .n32681(n32681), .n32740(n32740), 
            .n8177(n8177), .qspi_data_out_3__N_5({qspi_data_out_3__N_5}), 
            .\qspi_data_in[3] (\qspi_data_in[3] ), .\qspi_data_in[2] (\qspi_data_in[2] ), 
            .\read_cycles_count[1] (read_cycles_count[1]), .n32778(n32778), 
            .data_req_N_2334(data_req_N_2334), .qspi_ram_a_select(qspi_ram_a_select), 
            .qspi_ram_b_select(qspi_ram_b_select), .clk_N_45(clk_N_45), 
            .stop_txn_reg(stop_txn_reg), .n32521(n32521), .\qspi_data_oe[1] (\qspi_data_oe[1] ), 
            .clk_c_enable_341(clk_c_enable_341), .n1072(n1072), .n19867(n19867), 
            .debug_stop_txn(debug_stop_txn), .\writing_N_164[3] (\writing_N_164[3] ), 
            .n32542(n32542), .data_ready_N_2347(data_ready_N_2347), .n4513(n4513), 
            .n4501(n4501), .n32833(n32833), .n26811(n26811), .n4503(n4503), 
            .\addr[20]_adj_15 (\addr[20] ), .\addr[22]_adj_16 (\addr[22] ), 
            .n6218(n6218), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .qspi_clk_N_56(qspi_clk_N_56), .n6220(n6220), .n31866(n31866), 
            .clk_c_enable_543(clk_c_enable_543), .n28319(n28319), .n32874(n32874), 
            .n28259(n28259), .\qspi_data_in[0] (\qspi_data_in[0] ), .n332(n329[0]), 
            .n32060(n32060), .n28111(n28111), .n32789(n32789), .n32892(n32892)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(132[19] 164[6])
    tinyqv_cpu cpu (.imm({Open_44, Open_45, Open_46, Open_47, Open_48, 
            Open_49, Open_50, Open_51, Open_52, Open_53, Open_54, 
            Open_55, Open_56, Open_57, \imm[17] , \imm[16] , \imm[15] , 
            \imm[14] , Open_58, Open_59, Open_60, Open_61, Open_62, 
            Open_63, Open_64, Open_65, Open_66, Open_67, Open_68, 
            Open_69, Open_70, Open_71}), .clk_c(clk_c), .\instr[31] (\instr[31] ), 
            .\imm[13] (\imm[13] ), .n32578(n32578), .\imm[12] (\imm[12] ), 
            .\imm[11] (\imm[11] ), .\imm[10] (\imm[10] ), .\imm[9] (\imm[9] ), 
            .\imm[8] (\imm[8] ), .\imm[7] (\imm[7] ), .\imm[6] (\imm[6] ), 
            .\imm[5] (\imm[5] ), .\imm[4] (\imm[4] ), .\imm[3] (\imm[3] ), 
            .\imm[2] (\imm[2] ), .\imm[1] (\imm[1] ), .was_early_branch(was_early_branch), 
            .data_to_write({data_to_write_c[31:13], \data_to_write[12] , 
            \data_to_write[11] , \data_to_write[10] , \data_to_write[9] , 
            \data_to_write[8] , \data_to_write[7] , \data_to_write[6] , 
            \data_to_write[5] , \data_to_write[4] , \data_to_write[3] , 
            \data_to_write[2] , \data_to_write[1] , data_to_write[0]}), 
            .addr({\addr[27] , Open_72, Open_73, Open_74, Open_75, 
            Open_76, Open_77, Open_78, Open_79, Open_80, Open_81, 
            Open_82, Open_83, Open_84, Open_85, Open_86, Open_87, 
            \addr[10] , Open_88, Open_89, \addr[7] , \addr[6] , Open_90, 
            Open_91, \addr[3] , \addr[2] , Open_92, \addr[0] }), .rd({Open_93, 
            Open_94, Open_95, \rd[0] }), .qv_data_read_n({qv_data_read_n}), 
            .n29738(n29738), .\instr_data[3]_adj_13 ({Open_96, Open_97, 
            Open_98, Open_99, Open_100, Open_101, Open_102, Open_103, 
            Open_104, Open_105, Open_106, Open_107, Open_108, Open_109, 
            Open_110, \instr_data[3][0] }), .\instr_addr_23__N_318[0] (\instr_addr_23__N_318[0] ), 
            .n32656(n32656), .n26116(n26116), .debug_data_continue(debug_data_continue), 
            .debug_instr_valid(debug_instr_valid), .n32851(n32851), .n32835(n32835), 
            .n32723(n32723), .\gpio_out_func_sel[5][2] (\gpio_out_func_sel[5][2] ), 
            .\gpio_out_func_sel[7][2] (\gpio_out_func_sel[7][2] ), .\instr_len[2] (\instr_len[2] ), 
            .\pc[2] (\pc[2] ), .\pc[1] (\pc[1] ), .n2196(n2196), .n32727(n32727), 
            .n2191(n2191), .n32640(n32640), .instr_data({instr_data}), 
            .n32548(n32548), .n32734(n32734), .\qspi_data_buf[10] (qspi_data_buf[10]), 
            .\qspi_data_buf[14] (qspi_data_buf[14]), .n32836(n32836), .n27888(n27888), 
            .\gpio_out_func_sel[5][4] (\gpio_out_func_sel[5][4] ), .\gpio_out_func_sel[7][4] (\gpio_out_func_sel[7][4] ), 
            .n29831(n29831), .n32655(n32655), .n34287(n34287), .instr_fetch_running(instr_fetch_running), 
            .n32544(n32544), .n32537(n32537), .instr_fetch_running_N_945(instr_fetch_running_N_945), 
            .n19867(n19867), .\instr_write_offset[3] (\instr_write_offset[3] ), 
            .qspi_data_byte_idx({qspi_data_byte_idx}), .qspi_data_ready(qspi_data_ready), 
            .n2150(n2150), .n2130(n2130), .n4251(n4251), .n32685(n32685), 
            .n19(n19), .n32660(n32660), .\qspi_data_buf[11] (qspi_data_buf[11]), 
            .\qspi_data_buf[15] (qspi_data_buf[15]), .\peri_data_out[11] (\peri_data_out[11] ), 
            .n4(n4), .\peri_data_out[10] (\peri_data_out[10] ), .n32642(n32642), 
            .\mem_data_from_read[20] (mem_data_from_read[20]), .\mem_data_from_read[16] (mem_data_from_read[16]), 
            .n32771(n32771), .\peri_data_out[9] (\peri_data_out[9] ), .rst_reg_n_adj_6(rst_reg_n_adj_17), 
            .n31796(n31796), .n31795(n31795), .n32520(n32520), .n21414(n21414), 
            .n32654(n32654), .\pc[7] (\pc[7] ), .\pc[15] (\pc[15] ), .n32842(n32842), 
            .\next_pc_for_core[6] (\next_pc_for_core[6] ), .\pc[3] (\pc[3] ), 
            .\pc[11] (\pc[11] ), .n32251(n32251), .n31706(n31706), .clk_c_enable_285(clk_c_enable_285), 
            .n28957(n28957), .n34285(n34285), .\pc[6] (\pc[6] ), .\pc[14] (\pc[14] ), 
            .\pc[10] (\pc[10] ), .n3(n3), .n3_adj_7(n3_adj_18), .n32638(n32638), 
            .n29707(n29707), .qv_data_write_n({qv_data_write_n}), .n32850(n32850), 
            .\addr[24] (addr[24]), .\addr[23] (addr[23]), .\addr[22] (addr[22]), 
            .\addr[21] (addr[21]), .\imm[21] (\imm[21] ), .\imm[20] (\imm[20] ), 
            .\next_pc_for_core[9] (\next_pc_for_core[9] ), .\next_pc_for_core[13] (\next_pc_for_core[13] ), 
            .\addr[20] (addr[20]), .\addr[19] (addr[19]), .\addr[18] (addr[18]), 
            .\addr[17] (addr[17]), .\addr[16] (addr[16]), .\pc[5] (\pc[5] ), 
            .\pc[13] (\pc[13] ), .\addr[15] (addr[15]), .\pc[9] (\pc[9] ), 
            .\addr[14] (addr[14]), .\addr[13] (addr[13]), .\addr[12] (addr[12]), 
            .\addr[11] (addr[11]), .\addr[9] (addr[9]), .\addr[8] (addr[8]), 
            .\addr[5] (\addr[5] ), .\addr[4] (\addr[4] ), .\addr[1] (\addr[1] ), 
            .\next_pc_for_core[4] (\next_pc_for_core[4] ), .n12(n12), .data_ready_r_N_2823(data_ready_r_N_2823), 
            .data_ready_r(data_ready_r), .n32801(n32801), .n29059(n29059), 
            .n32598(n32598), .data_txn_len({data_txn_len}), .n32714(n32714), 
            .n32689(n32689), .n32531(n32531), .rst_reg_n(rst_reg_n), .n32706(n32706), 
            .n15569(n15569), .n2211(n2211), .n17165(n17165), .VCC_net(VCC_net), 
            .n32694(n32694), .n7(n7), .n8854(n8854), .\next_pc_for_core[10] (\next_pc_for_core[10] ), 
            .\next_pc_for_core[14] (\next_pc_for_core[14] ), .debug_stop_txn_N_2142(debug_stop_txn_N_2142), 
            .\instr_data[0][0] (\instr_data[0][0] ), .\instr_data[1][7] (\instr_data[1][7] ), 
            .\instr_data[1][0] (\instr_data[1][0] ), .\instr_data[2][7] (\instr_data[2][7] ), 
            .data_stall(data_stall), .n32542(n32542), .\next_pc_for_core[8] (\next_pc_for_core[8] ), 
            .\next_pc_for_core[12] (\next_pc_for_core[12] ), .n32787(n32787), 
            .n32740(n32740), .data_req_N_2334(data_req_N_2334), .n332(n329[0]), 
            .instr_active(instr_active), .n11193(n11193), .clk_c_enable_91(clk_c_enable_91), 
            .\mem_data_from_read[19] (mem_data_from_read[19]), .\mem_data_from_read[23] (mem_data_from_read[23]), 
            .n32788(n32788), .n1(n1), .n175(n174[1]), .\read_cycles_count[1] (read_cycles_count[1]), 
            .n32789(n32789), .data_ready_N_2347(data_ready_N_2347), .\instr_data[2][0] (\instr_data[2][0] ), 
            .\instr_data[3][7] (\instr_data[3][7] ), .n32545(n32545), .n32552(n32552), 
            .n8109(n8109), .n32695(n32695), .n32728(n32728), .n32712(n32712), 
            .n32745(n32745), .\next_pc_for_core[3] (\next_pc_for_core[3] ), 
            .\next_pc_for_core[5] (\next_pc_for_core[5] ), .\next_pc_for_core[7] (\next_pc_for_core[7] ), 
            .\next_pc_for_core[11] (\next_pc_for_core[11] ), .\pc[21] (\pc[21] ), 
            .\pc[17] (\pc[17] ), .\next_pc_for_core[20] (\next_pc_for_core[20] ), 
            .\next_pc_for_core[16] (\next_pc_for_core[16] ), .\pc[23] (\pc[23] ), 
            .\pc[19] (\pc[19] ), .\pc[22] (\pc[22] ), .\pc[18] (\pc[18] ), 
            .\pc[20] (\pc[20] ), .\pc[16] (\pc[16] ), .\next_pc_for_core[15] (\next_pc_for_core[15] ), 
            .\next_pc_for_core[21] (\next_pc_for_core[21] ), .\next_pc_for_core[17] (\next_pc_for_core[17] ), 
            .\imm[23] (\imm[23] ), .\imm[22] (\imm[22] ), .\imm[19] (\imm[19] ), 
            .\imm[18] (\imm[18] ), .\next_pc_for_core[22] (\next_pc_for_core[22] ), 
            .\next_pc_for_core[18] (\next_pc_for_core[18] ), .\next_pc_for_core[19] (\next_pc_for_core[19] ), 
            .n28077(n28077), .\next_pc_for_core[23] (\next_pc_for_core[23] ), 
            .n32819(n32819), .n32720(n32720), .n29357(n29357), .\uo_out_from_user_peri[1][6] (\uo_out_from_user_peri[1][6] ), 
            .\data_from_user_peri_1__31__N_2455[2] (\data_from_user_peri_1__31__N_2455[2] ), 
            .\uo_out_from_user_peri[1][2] (\uo_out_from_user_peri[1][2] ), 
            .\uo_out_from_user_peri[1][5] (\uo_out_from_user_peri[1][5] ), 
            .n29491(n29491), .\data_from_read[2] (\data_from_read[2] ), 
            .\early_branch_addr[7] (\early_branch_addr[7] ), .\early_branch_addr[3] (\early_branch_addr[3] ), 
            .\early_branch_addr[6] (\early_branch_addr[6] ), .\early_branch_addr[2] (\early_branch_addr[2] ), 
            .\early_branch_addr[4] (\early_branch_addr[4] ), .n32822(n32822), 
            .\early_branch_addr[8] (\early_branch_addr[8] ), .\early_branch_addr[5] (\early_branch_addr[5] ), 
            .\early_branch_addr[9] (\early_branch_addr[9] ), .\early_branch_addr[10] (\early_branch_addr[10] ), 
            .\early_branch_addr[11] (\early_branch_addr[11] ), .\early_branch_addr[12] (\early_branch_addr[12] ), 
            .\early_branch_addr[13] (\early_branch_addr[13] ), .\early_branch_addr[14] (\early_branch_addr[14] ), 
            .\early_branch_addr[15] (\early_branch_addr[15] ), .\early_branch_addr[17] (\early_branch_addr[17] ), 
            .\early_branch_addr[18] (\early_branch_addr[18] ), .\early_branch_addr[19] (\early_branch_addr[19] ), 
            .\early_branch_addr[20] (\early_branch_addr[20] ), .\early_branch_addr[21] (\early_branch_addr[21] ), 
            .\early_branch_addr[22] (\early_branch_addr[22] ), .\early_branch_addr[23] (\early_branch_addr[23] ), 
            .\early_branch_addr[16] (\early_branch_addr[16] ), .n16811(n16811), 
            .n2594(n2594), .n31883(n31883), .\pc_23__N_911[13] (\pc_23__N_911[13] ), 
            .\pc[12] (\pc[12] ), .n26838(n26838), .n10944(n10944), .n32725(n32725), 
            .n32761(n32761), .n32729(n32729), .\cycle[0] (\cycle[0] ), 
            .debug_data_ready(debug_data_ready), .\pc[8] (\pc[8] ), .n27178(n27178), 
            .n32766(n32766), .\pc[4] (\pc[4] ), .n32711(n32711), .n32737(n32737), 
            .\data_from_peri_31__N_2415[0] (\data_from_peri_31__N_2415[0] ), 
            .fsm_state({fsm_state_c[2:1], fsm_state[0]}), .n32778(n32778), 
            .n31866(n31866), .n32693(n32693), .clk_c_enable_50(clk_c_enable_50), 
            .n32818(n32818), .clk_c_enable_154(clk_c_enable_154), .clk_c_enable_283(clk_c_enable_283), 
            .clk_c_enable_354(clk_c_enable_354), .\gpio_out_func_sel[0][2] (\gpio_out_func_sel[0][2] ), 
            .\gpio_out_func_sel[1][2] (\gpio_out_func_sel[1][2] ), .\gpio_out_func_sel[2][2] (\gpio_out_func_sel[2][2] ), 
            .\gpio_out_func_sel[3][2] (\gpio_out_func_sel[3][2] ), .n32756(n32756), 
            .n5169(n5169), .n29618(n29618), .start_instr(start_instr), 
            .n32825(n32825), .n29127(n29127), .n18458(n18458), .\gpio_out_func_sel[4][2] (\gpio_out_func_sel[4][2] ), 
            .\gpio_out_func_sel[6][2] (\gpio_out_func_sel[6][2] ), .n8(n8), 
            .\uart_rx_buf_data[4] (\uart_rx_buf_data[4] ), .\baud_divider[4] (\baud_divider[4] ), 
            .instr_fetch_stopped(instr_fetch_stopped), .n16(n16), .n32826(n32826), 
            .\instr_data_7__N_1969[3] (instr_data_7__N_1969[3]), .\instr_data_7__N_1969[1] (instr_data_7__N_1969[1]), 
            .gpio_out_sel({gpio_out_sel}), .n14(n14), .n14_adj_8(n14_adj_19), 
            .n29293(n29293), .instr_complete_N_1647(instr_complete_N_1647), 
            .\data_from_read[6] (\data_from_read[6] ), .n32672(n32672), 
            .n46(n46), .\connect_peripheral[1] (\connect_peripheral[1] ), 
            .\connect_peripheral[0] (\connect_peripheral[0] ), .\qspi_data_buf[9] (qspi_data_buf[9]), 
            .\qspi_data_buf[13] (qspi_data_buf[13]), .\instr_addr[2] (instr_addr[2]), 
            .n32568(n32568), .n29741(n29741), .n29(n29), .\uart_rx_buf_data[7] (\uart_rx_buf_data[7] ), 
            .\baud_divider[7] (\baud_divider[7] ), .n2(n2), .n32614(n32614), 
            .\next_fsm_state_3__N_3046[3] (\next_fsm_state_3__N_3046[3] ), 
            .\ui_in_sync[5] (\ui_in_sync[5] ), .\ui_in_sync[6] (\ui_in_sync[6] ), 
            .n32072(n32072), .n29549(n29549), .\ui_in_sync[7] (\ui_in_sync[7] ), 
            .\data_from_user_peri_1__31__N_2455[7] (\data_from_user_peri_1__31__N_2455[7] ), 
            .\uart_rx_buf_data[6] (\uart_rx_buf_data[6] ), .n26856(n26856), 
            .\baud_divider[6] (\baud_divider[6] ), .\uart_rx_buf_data[5] (\uart_rx_buf_data[5] ), 
            .\baud_divider[5] (\baud_divider[5] ), .\mem_data_from_read[4] (mem_data_from_read[4]), 
            .\data_from_read[4] (\data_from_read[4] ), .\mem_data_from_read[8] (mem_data_from_read[8]), 
            .\data_from_read[8] (\data_from_read[8] ), .\mem_data_from_read[12] (mem_data_from_read[12]), 
            .\data_from_read[12] (\data_from_read[12] ), .\mem_data_from_read[1] (mem_data_from_read[1]), 
            .\data_from_read[1] (\data_from_read[1] ), .\data_from_user_peri_1__31__N_2455[0] (\data_from_user_peri_1__31__N_2455[0] ), 
            .\uo_out_from_user_peri[1][0] (\uo_out_from_user_peri[1][0] ), 
            .\mem_data_from_read[5] (mem_data_from_read[5]), .\data_from_read[5] (\data_from_read[5] ), 
            .data_out_hold(data_out_hold), .\mem_data_from_read[3] (mem_data_from_read[3]), 
            .\data_from_read[3] (\data_from_read[3] ), .\mem_data_from_read[7] (mem_data_from_read[7]), 
            .\data_from_read[7] (\data_from_read[7] ), .\uart_rx_buf_data[3] (\uart_rx_buf_data[3] ), 
            .\baud_divider[3] (\baud_divider[3] ), .n2_adj_9(n2_adj_20), 
            .\mem_data_from_read[0] (mem_data_from_read[0]), .\data_from_read[0] (\data_from_read[0] ), 
            .n32759(n32759), .\mem_data_from_read[18] (mem_data_from_read[18]), 
            .\mem_data_from_read[22] (mem_data_from_read[22]), .\mem_data_from_read[26] (mem_data_from_read[26]), 
            .\mem_data_from_read[30] (mem_data_from_read[30]), .\mem_data_from_read[24] (mem_data_from_read[24]), 
            .\mem_data_from_read[28] (mem_data_from_read[28]), .\uart_rx_buf_data[2] (\uart_rx_buf_data[2] ), 
            .\baud_divider[2] (\baud_divider[2] ), .\mem_data_from_read[27] (mem_data_from_read[27]), 
            .\mem_data_from_read[31] (mem_data_from_read[31]), .\mem_data_from_read[25] (mem_data_from_read[25]), 
            .\mem_data_from_read[29] (mem_data_from_read[29]), .n10737(n10737), 
            .n32650(n32650), .\instr[16] (\instr[16] ), .n32615(n32615), 
            .n32610(n32610), .clk_c_enable_342(clk_c_enable_342), .\ui_in_sync[1] (\ui_in_sync[1] ), 
            .\ui_in_sync[0] (\ui_in_sync[0] ), .debug_rd({debug_rd}), .n29866(n29866), 
            .n17920(n17920), .n28687(n28687), .accum({accum}), .d_3__N_1868({d_3__N_1868}), 
            .fsm_state_adj_14({fsm_state_adj_24}), .n32791(n32791), .n32763(n32763), 
            .n32730(n32730), .n32834(n32834), .n32710(n32710), .n31351(n31351), 
            .n1152(n1152), .\mem_data_from_read[17] (mem_data_from_read[17]), 
            .\mem_data_from_read[21] (mem_data_from_read[21]), .\mul_out[3] (\mul_out[3] ), 
            .\mul_out[2] (\mul_out[2] ), .\mul_out[1] (\mul_out[1] ), .\csr_read_3__N_1447[2] (\csr_read_3__N_1447[2] ), 
            .\next_accum[5] (\next_accum[5] ), .GND_net(GND_net), .\next_accum[16] (\next_accum[16] ), 
            .\next_accum[17] (\next_accum[17] ), .\next_accum[18] (\next_accum[18] ), 
            .\next_accum[19] (\next_accum[19] ), .\next_accum[6] (\next_accum[6] ), 
            .\next_accum[7] (\next_accum[7] ), .\next_accum[8] (\next_accum[8] ), 
            .\next_accum[9] (\next_accum[9] ), .\next_accum[10] (\next_accum[10] ), 
            .\next_accum[11] (\next_accum[11] ), .\next_accum[12] (\next_accum[12] ), 
            .\next_accum[13] (\next_accum[13] ), .\next_accum[14] (\next_accum[14] ), 
            .\next_accum[15] (\next_accum[15] ), .\next_accum[4] (\next_accum[4] ), 
            .\return_addr[16] (\return_addr[16] )) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(94[14] 130[6])
    
endmodule
//
// Verilog Description of module tinyqv_mem_ctrl
//

module tinyqv_mem_ctrl (instr_active, clk_c, instr_active_N_2106, start_instr, 
            qspi_data_byte_idx, data_txn_len, n26692, qspi_write_done, 
            instr_data, \instr_addr_23__N_318[7] , \addr[8] , \instr_addr_23__N_318[6] , 
            \addr[7] , \instr_addr_23__N_318[8] , \addr[9] , \instr_addr_23__N_318[20] , 
            \addr[21] , \instr_addr_23__N_318[21] , \addr[22] , \instr_addr_23__N_318[2] , 
            \addr[3] , \instr_addr[2] , \addr[2] , \mem_data_from_read[23] , 
            \mem_data_from_read[22] , \mem_data_from_read[21] , \mem_data_from_read[20] , 
            \mem_data_from_read[19] , \mem_data_from_read[18] , \mem_data_from_read[17] , 
            \mem_data_from_read[16] , \qspi_data_buf[15] , clk_c_enable_91, 
            \qspi_data_buf[14] , \qspi_data_buf[13] , \qspi_data_buf[11] , 
            \qspi_data_buf[10] , \qspi_data_buf[9] , \instr_data_7__N_1969[3] , 
            \instr_data_7__N_1969[1] , \instr_addr[1] , \addr[1] , mem_data_ready, 
            \mem_data_from_read[29] , \mem_data_from_read[25] , n32522, 
            \mem_data_from_read[31] , \mem_data_from_read[27] , \mem_data_from_read[28] , 
            \mem_data_from_read[24] , \mem_data_from_read[30] , \mem_data_from_read[26] , 
            n32755, clk_c_enable_432, debug_data_continue, n175, n26691, 
            instr_fetch_running_N_945, n10672, n32537, n11193, qspi_data_ready, 
            data_stall, rst_reg_n, n29887, n32523, n32826, n32712, 
            \addr[24] , n32598, \mem_data_from_read[0] , \mem_data_from_read[7] , 
            \mem_data_from_read[3] , \data_to_write[0] , \mem_data_from_read[5] , 
            \mem_data_from_read[1] , \mem_data_from_read[4] , instr_fetch_stopped, 
            n32531, is_writing_N_2331, \mem_data_from_read[12] , \mem_data_from_read[8] , 
            debug_stop_txn_N_2142, \data_to_write[31] , n32545, n8, 
            n28687, n16, \data_to_write[30] , \data_to_write[29] , \data_to_write[28] , 
            \data_to_write[27] , \data_to_write[26] , \data_to_write[25] , 
            \data_to_write[24] , \data_to_write[23] , \data_to_write[22] , 
            \data_to_write[21] , \data_to_write[20] , \data_to_write[19] , 
            \data_to_write[18] , \data_to_write[17] , \data_to_write[16] , 
            \data_to_write[15] , \data_to_write[14] , \data_to_write[13] , 
            \data_to_write[12] , \data_to_write[11] , \data_to_write[10] , 
            n32787, \data_to_write[9] , \data_to_write[8] , \data_to_write[7] , 
            \data_to_write[6] , \data_to_write[5] , \data_to_write[4] , 
            \data_to_write[2] , \addr[0] , n32711, n32714, continue_txn_N_2131, 
            data_stall_N_2158, n32788, n1, n32771, n32801, n21414, 
            n32689, \addr[23] , instr_fetch_running, n29618, \instr_addr_23__N_318[5] , 
            \addr[6] , \instr_addr_23__N_318[11] , \addr[12] , \instr_addr_23__N_318[14] , 
            \addr[15] , \instr_addr_23__N_318[9] , \addr[10] , \instr_addr_23__N_318[15] , 
            \addr[16] , \instr_addr_23__N_318[16] , \addr[17] , \instr_addr_23__N_318[17] , 
            \addr[18] , \instr_addr_23__N_318[12] , \addr[13] , n32578, 
            \instr_addr_23__N_318[10] , \addr[11] , \instr_addr_23__N_318[13] , 
            \addr[14] , \instr_addr_23__N_318[3] , \addr[4] , is_writing, 
            spi_clk_pos, stop_txn_now_N_2363, \instr_addr_23__N_318[22] , 
            \instr_addr_23__N_318[4] , \addr[5] , \instr_addr_23__N_318[19] , 
            \addr[20] , \instr_addr_23__N_318[18] , \addr[19] , fsm_state, 
            clk_c_enable_340, n32524, clk_c_enable_208, clk_c_enable_66, 
            n29884, n27931, n32681, n32740, n8177, qspi_data_out_3__N_5, 
            \qspi_data_in[3] , \qspi_data_in[2] , \read_cycles_count[1] , 
            n32778, data_req_N_2334, qspi_ram_a_select, qspi_ram_b_select, 
            clk_N_45, stop_txn_reg, n32521, \qspi_data_oe[1] , clk_c_enable_341, 
            n1072, n19867, debug_stop_txn, \writing_N_164[3] , n32542, 
            data_ready_N_2347, n4513, n4501, n32833, n26811, n4503, 
            \addr[20]_adj_15 , \addr[22]_adj_16 , n6218, spi_clk_pos_derived_59, 
            qspi_clk_N_56, n6220, n31866, clk_c_enable_543, n28319, 
            n32874, n28259, \qspi_data_in[0] , n332, n32060, n28111, 
            n32789, n32892) /* synthesis syn_module_defined=1 */ ;
    output instr_active;
    input clk_c;
    input instr_active_N_2106;
    input start_instr;
    output [1:0]qspi_data_byte_idx;
    output [1:0]data_txn_len;
    input n26692;
    output qspi_write_done;
    output [15:0]instr_data;
    input \instr_addr_23__N_318[7] ;
    input \addr[8] ;
    input \instr_addr_23__N_318[6] ;
    input \addr[7] ;
    input \instr_addr_23__N_318[8] ;
    input \addr[9] ;
    input \instr_addr_23__N_318[20] ;
    input \addr[21] ;
    input \instr_addr_23__N_318[21] ;
    input \addr[22] ;
    input \instr_addr_23__N_318[2] ;
    input \addr[3] ;
    input \instr_addr[2] ;
    input \addr[2] ;
    output \mem_data_from_read[23] ;
    output \mem_data_from_read[22] ;
    output \mem_data_from_read[21] ;
    output \mem_data_from_read[20] ;
    output \mem_data_from_read[19] ;
    output \mem_data_from_read[18] ;
    output \mem_data_from_read[17] ;
    output \mem_data_from_read[16] ;
    output \qspi_data_buf[15] ;
    input clk_c_enable_91;
    output \qspi_data_buf[14] ;
    output \qspi_data_buf[13] ;
    output \qspi_data_buf[11] ;
    output \qspi_data_buf[10] ;
    output \qspi_data_buf[9] ;
    input \instr_data_7__N_1969[3] ;
    input \instr_data_7__N_1969[1] ;
    input \instr_addr[1] ;
    input \addr[1] ;
    output mem_data_ready;
    output \mem_data_from_read[29] ;
    output \mem_data_from_read[25] ;
    output n32522;
    output \mem_data_from_read[31] ;
    output \mem_data_from_read[27] ;
    output \mem_data_from_read[28] ;
    output \mem_data_from_read[24] ;
    output \mem_data_from_read[30] ;
    output \mem_data_from_read[26] ;
    output n32755;
    input clk_c_enable_432;
    input debug_data_continue;
    input n175;
    input n26691;
    output instr_fetch_running_N_945;
    input n10672;
    input n32537;
    output n11193;
    output qspi_data_ready;
    output data_stall;
    input rst_reg_n;
    input n29887;
    output n32523;
    output n32826;
    input n32712;
    input \addr[24] ;
    output n32598;
    output \mem_data_from_read[0] ;
    output \mem_data_from_read[7] ;
    output \mem_data_from_read[3] ;
    input \data_to_write[0] ;
    output \mem_data_from_read[5] ;
    output \mem_data_from_read[1] ;
    output \mem_data_from_read[4] ;
    output instr_fetch_stopped;
    input n32531;
    output is_writing_N_2331;
    output \mem_data_from_read[12] ;
    output \mem_data_from_read[8] ;
    input debug_stop_txn_N_2142;
    input \data_to_write[31] ;
    input n32545;
    input n8;
    input n28687;
    output n16;
    input \data_to_write[30] ;
    input \data_to_write[29] ;
    input \data_to_write[28] ;
    input \data_to_write[27] ;
    input \data_to_write[26] ;
    input \data_to_write[25] ;
    input \data_to_write[24] ;
    input \data_to_write[23] ;
    input \data_to_write[22] ;
    input \data_to_write[21] ;
    input \data_to_write[20] ;
    input \data_to_write[19] ;
    input \data_to_write[18] ;
    input \data_to_write[17] ;
    input \data_to_write[16] ;
    input \data_to_write[15] ;
    input \data_to_write[14] ;
    input \data_to_write[13] ;
    input \data_to_write[12] ;
    input \data_to_write[11] ;
    input \data_to_write[10] ;
    input n32787;
    input \data_to_write[9] ;
    input \data_to_write[8] ;
    input \data_to_write[7] ;
    input \data_to_write[6] ;
    input \data_to_write[5] ;
    input \data_to_write[4] ;
    input \data_to_write[2] ;
    input \addr[0] ;
    input n32711;
    input n32714;
    output continue_txn_N_2131;
    output data_stall_N_2158;
    input n32788;
    output n1;
    input n32771;
    input n32801;
    input n21414;
    output n32689;
    input \addr[23] ;
    input instr_fetch_running;
    output n29618;
    input \instr_addr_23__N_318[5] ;
    input \addr[6] ;
    input \instr_addr_23__N_318[11] ;
    input \addr[12] ;
    input \instr_addr_23__N_318[14] ;
    input \addr[15] ;
    input \instr_addr_23__N_318[9] ;
    input \addr[10] ;
    input \instr_addr_23__N_318[15] ;
    input \addr[16] ;
    input \instr_addr_23__N_318[16] ;
    input \addr[17] ;
    input \instr_addr_23__N_318[17] ;
    input \addr[18] ;
    input \instr_addr_23__N_318[12] ;
    input \addr[13] ;
    output n32578;
    input \instr_addr_23__N_318[10] ;
    input \addr[11] ;
    input \instr_addr_23__N_318[13] ;
    input \addr[14] ;
    input \instr_addr_23__N_318[3] ;
    input \addr[4] ;
    output is_writing;
    output spi_clk_pos;
    output stop_txn_now_N_2363;
    input \instr_addr_23__N_318[22] ;
    input \instr_addr_23__N_318[4] ;
    input \addr[5] ;
    input \instr_addr_23__N_318[19] ;
    input \addr[20] ;
    input \instr_addr_23__N_318[18] ;
    input \addr[19] ;
    output [2:0]fsm_state;
    input clk_c_enable_340;
    input n32524;
    input clk_c_enable_208;
    input clk_c_enable_66;
    input n29884;
    input n27931;
    output n32681;
    output n32740;
    input n8177;
    input [3:0]qspi_data_out_3__N_5;
    input \qspi_data_in[3] ;
    input \qspi_data_in[2] ;
    output \read_cycles_count[1] ;
    output n32778;
    output data_req_N_2334;
    output qspi_ram_a_select;
    output qspi_ram_b_select;
    input clk_N_45;
    output stop_txn_reg;
    output n32521;
    output \qspi_data_oe[1] ;
    input clk_c_enable_341;
    output n1072;
    input n19867;
    output debug_stop_txn;
    output \writing_N_164[3] ;
    input n32542;
    input data_ready_N_2347;
    output n4513;
    output n4501;
    output n32833;
    output n26811;
    output n4503;
    output \addr[20]_adj_15 ;
    output \addr[22]_adj_16 ;
    output n6218;
    output spi_clk_pos_derived_59;
    output qspi_clk_N_56;
    output n6220;
    input n31866;
    input clk_c_enable_543;
    output n28319;
    output n32874;
    input n28259;
    input \qspi_data_in[0] ;
    input n332;
    output n32060;
    output n28111;
    input n32789;
    output n32892;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    
    wire clk_c_enable_31, clk_c_enable_144, qspi_data_byte_idx_1__N_2025, 
        n9, clk_c_enable_218, n11684, data_ready_N_2109, clk_c_enable_98;
    wire [31:0]instr_data_7__N_1969;
    wire [24:0]addr_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(57[17:24])
    wire [31:0]qspi_data_buf;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(58[16:29])
    
    wire clk_c_enable_75, clk_c_enable_83, n32648, ram_b_block_N_2303, 
        ram_a_block_N_2299, n482, clk_c_enable_488, n11756, continue_txn, 
        clk_c_enable_118, n32809, n32810, n34272, n6071, n32687, 
        n32669, n32528, data_ready_N_2113;
    wire [1:0]write_qspi_data_byte_idx_1__N_2021;
    
    wire n32649, n29768, n29771, n29774, n29777, n29764, n29761, 
        n29755, n31677, n31646, n31639, n31475, n29752, n29767, 
        n29770, n29773, n29776, n6704, n28383, data_ready_N_2108, 
        n31, n32526, n28127, last_ram_b_sel, n32686, n32534, debug_stop_txn_N_2120, 
        n8205, debug_stop_txn_N_2119, n28419;
    wire [23:0]addr_23__N_2188;
    
    wire n32715, n29319, spi_ram_b_select_N_2313, n3, spi_ram_a_select_N_2309;
    
    FD1P3IX instr_active_180 (.D(start_instr), .SP(clk_c_enable_31), .CD(instr_active_N_2106), 
            .CK(clk_c), .Q(instr_active)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(103[12] 109[8])
    defparam instr_active_180.GSR = "DISABLED";
    FD1P3IX qspi_data_byte_idx__i0 (.D(n9), .SP(clk_c_enable_144), .CD(qspi_data_byte_idx_1__N_2025), 
            .CK(clk_c), .Q(qspi_data_byte_idx[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam qspi_data_byte_idx__i0.GSR = "DISABLED";
    FD1P3AX data_txn_len_i0_i0 (.D(n26692), .SP(clk_c_enable_218), .CK(clk_c), 
            .Q(data_txn_len[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(177[12] 183[8])
    defparam data_txn_len_i0_i0.GSR = "DISABLED";
    FD1S3IX qspi_write_done_185 (.D(data_ready_N_2109), .CK(clk_c), .CD(n11684), 
            .Q(qspi_write_done)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(173[12] 175[8])
    defparam qspi_write_done_185.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i1 (.D(instr_data_7__N_1969[0]), .SP(clk_c_enable_98), 
            .CK(clk_c), .Q(instr_data[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i1.GSR = "DISABLED";
    LUT4 i12917_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr_23__N_318[7] ), 
         .D(\addr[8] ), .Z(addr_in[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i12917_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i8_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[6] ), .D(\addr[7] ), .Z(addr_in[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i8_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX qspi_data_buf_i32 (.D(instr_data_7__N_1969[31]), .SP(clk_c_enable_75), 
            .CK(clk_c), .Q(qspi_data_buf[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i32.GSR = "DISABLED";
    LUT4 i12925_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr_23__N_318[8] ), 
         .D(\addr[9] ), .Z(addr_in[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i12925_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i22_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[20] ), .D(\addr[21] ), .Z(addr_in[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i23_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[21] ), .D(\addr[22] ), .Z(addr_in[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i4_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[2] ), .D(\addr[3] ), .Z(addr_in[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i3_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr[2] ), .D(\addr[2] ), .Z(addr_in[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i3_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX qspi_data_buf_i31 (.D(instr_data_7__N_1969[30]), .SP(clk_c_enable_75), 
            .CK(clk_c), .Q(qspi_data_buf[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i31.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i30 (.D(instr_data_7__N_1969[29]), .SP(clk_c_enable_75), 
            .CK(clk_c), .Q(qspi_data_buf[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i30.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i29 (.D(instr_data_7__N_1969[28]), .SP(clk_c_enable_75), 
            .CK(clk_c), .Q(qspi_data_buf[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i29.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i28 (.D(instr_data_7__N_1969[27]), .SP(clk_c_enable_75), 
            .CK(clk_c), .Q(qspi_data_buf[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i28.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i27 (.D(instr_data_7__N_1969[26]), .SP(clk_c_enable_75), 
            .CK(clk_c), .Q(qspi_data_buf[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i27.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i26 (.D(instr_data_7__N_1969[25]), .SP(clk_c_enable_75), 
            .CK(clk_c), .Q(qspi_data_buf[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i26.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i25 (.D(instr_data_7__N_1969[24]), .SP(clk_c_enable_75), 
            .CK(clk_c), .Q(qspi_data_buf[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i25.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i24 (.D(instr_data_7__N_1969[23]), .SP(clk_c_enable_83), 
            .CK(clk_c), .Q(\mem_data_from_read[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i24.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i23 (.D(instr_data_7__N_1969[22]), .SP(clk_c_enable_83), 
            .CK(clk_c), .Q(\mem_data_from_read[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i23.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i22 (.D(instr_data_7__N_1969[21]), .SP(clk_c_enable_83), 
            .CK(clk_c), .Q(\mem_data_from_read[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i22.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i21 (.D(instr_data_7__N_1969[20]), .SP(clk_c_enable_83), 
            .CK(clk_c), .Q(\mem_data_from_read[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i21.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i20 (.D(instr_data_7__N_1969[19]), .SP(clk_c_enable_83), 
            .CK(clk_c), .Q(\mem_data_from_read[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i20.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i19 (.D(instr_data_7__N_1969[18]), .SP(clk_c_enable_83), 
            .CK(clk_c), .Q(\mem_data_from_read[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i19.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i18 (.D(instr_data_7__N_1969[17]), .SP(clk_c_enable_83), 
            .CK(clk_c), .Q(\mem_data_from_read[17] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i18.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i17 (.D(instr_data_7__N_1969[16]), .SP(clk_c_enable_83), 
            .CK(clk_c), .Q(\mem_data_from_read[16] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i17.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i16 (.D(instr_data_7__N_1969[15]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(\qspi_data_buf[15] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i16.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i15 (.D(instr_data_7__N_1969[14]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(\qspi_data_buf[14] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i15.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i14 (.D(instr_data_7__N_1969[13]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(\qspi_data_buf[13] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i14.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i13 (.D(instr_data_7__N_1969[12]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(qspi_data_buf[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i13.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i12 (.D(instr_data_7__N_1969[11]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(\qspi_data_buf[11] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i12.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i11 (.D(instr_data_7__N_1969[10]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(\qspi_data_buf[10] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i11.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i10 (.D(instr_data_7__N_1969[9]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(\qspi_data_buf[9] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i10.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i9 (.D(instr_data_7__N_1969[8]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(qspi_data_buf[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i9.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i8 (.D(instr_data_7__N_1969[7]), .SP(clk_c_enable_98), 
            .CK(clk_c), .Q(instr_data[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i8.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i7 (.D(instr_data_7__N_1969[6]), .SP(clk_c_enable_98), 
            .CK(clk_c), .Q(instr_data[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i7.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i6 (.D(instr_data_7__N_1969[5]), .SP(clk_c_enable_98), 
            .CK(clk_c), .Q(instr_data[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i6.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i5 (.D(instr_data_7__N_1969[4]), .SP(clk_c_enable_98), 
            .CK(clk_c), .Q(instr_data[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i5.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i4 (.D(\instr_data_7__N_1969[3] ), .SP(clk_c_enable_98), 
            .CK(clk_c), .Q(instr_data[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i4.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i3 (.D(instr_data_7__N_1969[2]), .SP(clk_c_enable_98), 
            .CK(clk_c), .Q(instr_data[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i3.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i2 (.D(\instr_data_7__N_1969[1] ), .SP(clk_c_enable_98), 
            .CK(clk_c), .Q(instr_data[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i2.GSR = "DISABLED";
    LUT4 i12849_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr[1] ), 
         .D(\addr[1] ), .Z(addr_in[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i12849_3_lut_4_lut.init = 16'hf1e0;
    LUT4 qspi_data_buf_29__I_0_3_lut (.A(qspi_data_buf[29]), .B(instr_data[13]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[29] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_29__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_25__I_0_3_lut (.A(qspi_data_buf[25]), .B(instr_data[9]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[25] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_25__I_0_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_507_3_lut_4_lut (.A(n32648), .B(start_instr), .C(ram_b_block_N_2303), 
         .D(ram_a_block_N_2299), .Z(n32522)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i1_2_lut_rep_507_3_lut_4_lut.init = 16'hd000;
    LUT4 qspi_data_buf_31__I_0_189_3_lut (.A(qspi_data_buf[31]), .B(instr_data[15]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[31] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_31__I_0_189_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_27__I_0_3_lut (.A(qspi_data_buf[27]), .B(instr_data[11]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[27] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_27__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_28__I_0_3_lut (.A(qspi_data_buf[28]), .B(instr_data[12]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[28] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_28__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_24__I_0_3_lut (.A(qspi_data_buf[24]), .B(instr_data[8]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_24__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_30__I_0_3_lut (.A(qspi_data_buf[30]), .B(instr_data[14]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[30] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_30__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_26__I_0_3_lut (.A(qspi_data_buf[26]), .B(instr_data[10]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[26] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_26__I_0_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32648), .B(start_instr), .C(n482), 
         .D(n32755), .Z(clk_c_enable_488)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf0fd;
    LUT4 i9048_2_lut_3_lut_4_lut (.A(n32648), .B(start_instr), .C(n482), 
         .D(n32755), .Z(n11756)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i9048_2_lut_3_lut_4_lut.init = 16'hf020;
    FD1P3IX continue_txn_187 (.D(debug_data_continue), .SP(clk_c_enable_118), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(continue_txn)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam continue_txn_187.GSR = "DISABLED";
    FD1P3IX qspi_data_byte_idx__i1 (.D(n175), .SP(clk_c_enable_144), .CD(qspi_data_byte_idx_1__N_2025), 
            .CK(clk_c), .Q(qspi_data_byte_idx[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam qspi_data_byte_idx__i1.GSR = "DISABLED";
    FD1P3AX data_txn_len_i0_i1 (.D(n26691), .SP(clk_c_enable_218), .CK(clk_c), 
            .Q(data_txn_len[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(177[12] 183[8])
    defparam data_txn_len_i0_i1.GSR = "DISABLED";
    FD1S3IX instr_fetch_started_181 (.D(n32537), .CK(clk_c), .CD(n10672), 
            .Q(instr_fetch_running_N_945)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam instr_fetch_started_181.GSR = "DISABLED";
    LUT4 equal_180_i3_2_lut_rep_794 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n32809)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(164[13:59])
    defparam equal_180_i3_2_lut_rep_794.init = 16'hbbbb;
    LUT4 i28388_2_lut_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n11193), .D(qspi_data_ready), .Z(clk_c_enable_83)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C)+!B !((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(164[13:59])
    defparam i28388_2_lut_3_lut_4_lut.init = 16'h40f0;
    LUT4 i15128_2_lut_rep_795 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n32810)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15128_2_lut_rep_795.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_591 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n11193), .D(qspi_data_ready), .Z(clk_c_enable_75)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_591.init = 16'h80f0;
    LUT4 instr_active_I_0_2_lut_rep_840 (.A(instr_active), .B(start_instr), 
         .Z(n34272)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam instr_active_I_0_2_lut_rep_840.init = 16'heeee;
    FD1P3IX data_stall_188 (.D(n29887), .SP(rst_reg_n), .CD(n6071), .CK(clk_c), 
            .Q(data_stall)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam data_stall_188.GSR = "DISABLED";
    LUT4 addr_23__I_201_2_lut_rep_513_3_lut_4_lut (.A(n32687), .B(n32669), 
         .C(n32755), .D(start_instr), .Z(n32528)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (C))) */ ;
    defparam addr_23__I_201_2_lut_rep_513_3_lut_4_lut.init = 16'h0f07;
    LUT4 i1_2_lut_rep_508_3_lut_4_lut (.A(n32687), .B(n32669), .C(ram_a_block_N_2299), 
         .D(start_instr), .Z(n32523)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_rep_508_3_lut_4_lut.init = 16'hf070;
    LUT4 i2_2_lut_4_lut (.A(n32687), .B(n32669), .C(rst_reg_n), .D(start_instr), 
         .Z(qspi_data_byte_idx_1__N_2025)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i2_2_lut_4_lut.init = 16'hff7f;
    LUT4 i1_2_lut_rep_811 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n32826)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam i1_2_lut_rep_811.init = 16'heeee;
    LUT4 i28446_2_lut_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n11193), .D(qspi_data_ready), .Z(clk_c_enable_98)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam i28446_2_lut_3_lut_4_lut.init = 16'h10f0;
    LUT4 i1_2_lut_3_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(data_stall), .Z(data_ready_N_2113)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_3_lut_4_lut (.A(qspi_data_ready), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(start_instr), .D(n32649), .Z(clk_c_enable_144)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[26:60])
    defparam i1_3_lut_4_lut.init = 16'hfeff;
    LUT4 i27059_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[28]), .D(\mem_data_from_read[20] ), .Z(n29768)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27059_3_lut_4_lut.init = 16'hf960;
    LUT4 i27062_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[29]), .D(\mem_data_from_read[21] ), .Z(n29771)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27062_3_lut_4_lut.init = 16'hf960;
    LUT4 i27065_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[30]), .D(\mem_data_from_read[22] ), .Z(n29774)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27065_3_lut_4_lut.init = 16'hf960;
    LUT4 i27068_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[31]), .D(\mem_data_from_read[23] ), .Z(n29777)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27068_3_lut_4_lut.init = 16'hf960;
    LUT4 i27055_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[11] ), .D(instr_data[3]), .Z(n29764)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27055_3_lut_4_lut.init = 16'hf960;
    LUT4 i27052_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[10] ), .D(instr_data[2]), .Z(n29761)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27052_3_lut_4_lut.init = 16'hf960;
    LUT4 i27046_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[9] ), .D(instr_data[1]), .Z(n29755)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27046_3_lut_4_lut.init = 16'hf960;
    LUT4 n5554_bdd_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[25]), .D(\mem_data_from_read[17] ), .Z(n31677)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n5554_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 n18361_bdd_3_lut_29182_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[26]), .D(\mem_data_from_read[18] ), .Z(n31646)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n18361_bdd_3_lut_29182_4_lut.init = 16'hf960;
    LUT4 n18361_bdd_3_lut_28794_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[27]), .D(\mem_data_from_read[19] ), .Z(n31639)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n18361_bdd_3_lut_28794_4_lut.init = 16'hf960;
    LUT4 n18361_bdd_3_lut_28721_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[24]), .D(\mem_data_from_read[16] ), .Z(n31475)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n18361_bdd_3_lut_28721_4_lut.init = 16'hf960;
    LUT4 i27043_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[8]), .D(instr_data[0]), .Z(n29752)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27043_3_lut_4_lut.init = 16'hf960;
    LUT4 i27058_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[12]), .D(instr_data[4]), .Z(n29767)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27058_3_lut_4_lut.init = 16'hf960;
    LUT4 i27061_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[13] ), .D(instr_data[5]), .Z(n29770)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27061_3_lut_4_lut.init = 16'hf960;
    LUT4 i27064_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[14] ), .D(instr_data[6]), .Z(n29773)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27064_3_lut_4_lut.init = 16'hf960;
    LUT4 i27067_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[15] ), .D(instr_data[7]), .Z(n29776)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i27067_3_lut_4_lut.init = 16'hf960;
    LUT4 i4422_2_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .Z(n6704)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i4422_2_lut.init = 16'h8888;
    LUT4 i28397_4_lut (.A(qspi_data_byte_idx[0]), .B(n28383), .C(start_instr), 
         .D(instr_active), .Z(n9)) /* synthesis lut_function=(!(A+!((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(155[17] 157[20])
    defparam i28397_4_lut.init = 16'h5551;
    LUT4 i1_3_lut (.A(data_txn_len[0]), .B(data_txn_len[1]), .C(qspi_data_byte_idx[1]), 
         .Z(n28383)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C)))) */ ;
    defparam i1_3_lut.init = 16'h4141;
    LUT4 data_ready_I_0_206_4_lut (.A(instr_active), .B(data_ready_N_2108), 
         .C(n32712), .D(n31), .Z(mem_data_ready)) /* synthesis lut_function=(!(A+!(B+!(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[25:190])
    defparam data_ready_I_0_206_4_lut.init = 16'h4544;
    LUT4 qspi_data_ready_I_0_202_2_lut (.A(qspi_data_ready), .B(data_ready_N_2109), 
         .Z(data_ready_N_2108)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[43:98])
    defparam qspi_data_ready_I_0_202_2_lut.init = 16'h8888;
    LUT4 i28314_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(data_txn_len[0]), .D(data_txn_len[1]), .Z(data_ready_N_2109)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[64:98])
    defparam i28314_4_lut.init = 16'h8421;
    LUT4 i1_4_lut (.A(start_instr), .B(n32526), .C(\addr[24] ), .D(n28127), 
         .Z(ram_b_block_N_2303)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_4_lut.init = 16'hffbf;
    LUT4 i1_2_lut (.A(instr_active), .B(last_ram_b_sel), .Z(n28127)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 instr_data_7__I_0_i1_3_lut_4_lut (.A(data_txn_len[0]), .B(n32598), 
         .C(instr_data[8]), .D(instr_data[0]), .Z(\mem_data_from_read[0] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i8_3_lut_4_lut (.A(data_txn_len[0]), .B(n32598), 
         .C(instr_data[15]), .D(instr_data[7]), .Z(\mem_data_from_read[7] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_519_3_lut_4_lut (.A(n32712), .B(n32686), .C(start_instr), 
         .D(n32687), .Z(n32534)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam i1_2_lut_rep_519_3_lut_4_lut.init = 16'hf1ff;
    LUT4 instr_data_7__I_0_i4_3_lut_4_lut (.A(data_txn_len[0]), .B(n32598), 
         .C(instr_data[11]), .D(instr_data[3]), .Z(\mem_data_from_read[3] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 i28296_2_lut_3_lut_4_lut (.A(n32712), .B(n32686), .C(rst_reg_n), 
         .D(n32687), .Z(clk_c_enable_218)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam i28296_2_lut_3_lut_4_lut.init = 16'h1fff;
    LUT4 i1_3_lut_rep_634_4_lut (.A(n32712), .B(n32686), .C(rst_reg_n), 
         .D(n32687), .Z(n32649)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i1_3_lut_rep_634_4_lut.init = 16'he000;
    LUT4 instr_data_7__I_173_i1_3_lut (.A(\data_to_write[0] ), .B(instr_data[8]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i1_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_0_i6_3_lut_4_lut (.A(data_txn_len[0]), .B(n32598), 
         .C(instr_data[13]), .D(instr_data[5]), .Z(\mem_data_from_read[5] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i2_3_lut_4_lut (.A(data_txn_len[0]), .B(n32598), 
         .C(instr_data[9]), .D(instr_data[1]), .Z(\mem_data_from_read[1] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i5_3_lut_4_lut (.A(data_txn_len[0]), .B(n32598), 
         .C(instr_data[12]), .D(instr_data[4]), .Z(\mem_data_from_read[4] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut_4_lut (.A(continue_txn), .B(data_ready_N_2109), 
         .C(write_qspi_data_byte_idx_1__N_2021[0]), .D(qspi_data_ready), 
         .Z(debug_stop_txn_N_2120)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[102:115])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h4440;
    FD1S3IX instr_fetch_stopped_182 (.D(debug_stop_txn_N_2119), .CK(clk_c), 
            .CD(n8205), .Q(instr_fetch_stopped)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam instr_fetch_stopped_182.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_592 (.A(start_instr), .B(n32531), .C(n32687), .D(n28419), 
         .Z(is_writing_N_2331)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_592.init = 16'h1000;
    LUT4 qspi_data_buf_15__I_0_i5_3_lut_4_lut (.A(data_txn_len[0]), .B(n32598), 
         .C(instr_data[12]), .D(qspi_data_buf[12]), .Z(\mem_data_from_read[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam qspi_data_buf_15__I_0_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 qspi_data_buf_15__I_0_i1_3_lut_4_lut (.A(data_txn_len[0]), .B(n32598), 
         .C(instr_data[8]), .D(qspi_data_buf[8]), .Z(\mem_data_from_read[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam qspi_data_buf_15__I_0_i1_3_lut_4_lut.init = 16'hf780;
    PFUMX debug_stop_txn_I_182 (.BLUT(debug_stop_txn_N_2120), .ALUT(debug_stop_txn_N_2142), 
          .C0(instr_active), .Z(debug_stop_txn_N_2119)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;
    LUT4 i8889_3_lut (.A(\data_to_write[31] ), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8889_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_593 (.A(instr_fetch_running_N_945), .B(n32545), .C(n8), 
         .D(n28687), .Z(n16)) /* synthesis lut_function=(A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam i1_4_lut_adj_593.init = 16'ha2aa;
    LUT4 i8891_3_lut (.A(\data_to_write[30] ), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8891_3_lut.init = 16'hcaca;
    LUT4 i8893_3_lut (.A(\data_to_write[29] ), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8893_3_lut.init = 16'hcaca;
    LUT4 i8895_3_lut (.A(\data_to_write[28] ), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8895_3_lut.init = 16'hcaca;
    LUT4 i8897_3_lut (.A(\data_to_write[27] ), .B(instr_data[11]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8897_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i27_4_lut (.A(\data_to_write[26] ), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n32810), .Z(instr_data_7__N_1969[26])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i27_4_lut.init = 16'hca0a;
    LUT4 instr_data_7__I_173_i26_4_lut (.A(\data_to_write[25] ), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n32810), .Z(instr_data_7__N_1969[25])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i26_4_lut.init = 16'hca0a;
    LUT4 instr_data_7__I_173_i25_4_lut (.A(\data_to_write[24] ), .B(instr_data[8]), 
         .C(qspi_data_ready), .D(n32810), .Z(instr_data_7__N_1969[24])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i25_4_lut.init = 16'hca0a;
    LUT4 i8899_3_lut (.A(\data_to_write[23] ), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8899_3_lut.init = 16'hcaca;
    LUT4 i8901_3_lut (.A(\data_to_write[22] ), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8901_3_lut.init = 16'hcaca;
    LUT4 i8903_3_lut (.A(\data_to_write[21] ), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8903_3_lut.init = 16'hcaca;
    LUT4 i8905_3_lut (.A(\data_to_write[20] ), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8905_3_lut.init = 16'hcaca;
    LUT4 i8907_3_lut (.A(\data_to_write[19] ), .B(instr_data[11]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8907_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i19_4_lut (.A(\data_to_write[18] ), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n32809), .Z(instr_data_7__N_1969[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i19_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i18_4_lut (.A(\data_to_write[17] ), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n32809), .Z(instr_data_7__N_1969[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i18_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i17_4_lut (.A(\data_to_write[16] ), .B(instr_data[8]), 
         .C(qspi_data_ready), .D(n32809), .Z(instr_data_7__N_1969[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i17_4_lut.init = 16'h0aca;
    LUT4 i8909_3_lut (.A(\data_to_write[15] ), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8909_3_lut.init = 16'hcaca;
    LUT4 i8911_3_lut (.A(\data_to_write[14] ), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8911_3_lut.init = 16'hcaca;
    LUT4 i8913_3_lut (.A(\data_to_write[13] ), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8913_3_lut.init = 16'hcaca;
    LUT4 i8915_3_lut (.A(\data_to_write[12] ), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8915_3_lut.init = 16'hcaca;
    LUT4 i8917_3_lut (.A(\data_to_write[11] ), .B(instr_data[11]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8917_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i11_4_lut (.A(\data_to_write[10] ), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n32787), .Z(instr_data_7__N_1969[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i11_4_lut.init = 16'hca0a;
    LUT4 instr_data_7__I_173_i10_4_lut (.A(\data_to_write[9] ), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n32787), .Z(instr_data_7__N_1969[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i10_4_lut.init = 16'hca0a;
    LUT4 instr_data_7__I_173_i9_4_lut (.A(\data_to_write[8] ), .B(instr_data[8]), 
         .C(qspi_data_ready), .D(n32787), .Z(instr_data_7__N_1969[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i9_4_lut.init = 16'hca0a;
    LUT4 i8919_3_lut (.A(\data_to_write[7] ), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8919_3_lut.init = 16'hcaca;
    LUT4 i8921_3_lut (.A(\data_to_write[6] ), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8921_3_lut.init = 16'hcaca;
    LUT4 i8923_3_lut (.A(\data_to_write[5] ), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8923_3_lut.init = 16'hcaca;
    LUT4 i8925_3_lut (.A(\data_to_write[4] ), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8925_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i3_4_lut (.A(\data_to_write[2] ), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n32826), .Z(instr_data_7__N_1969[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i3_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_594 (.A(n32531), .B(n32528), .C(instr_active), .D(\addr[0] ), 
         .Z(addr_23__N_2188[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_594.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_adj_595 (.A(n32711), .B(n32715), .C(data_ready_N_2113), 
         .D(n32712), .Z(n31)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(91[18] 99[12])
    defparam i1_2_lut_3_lut_4_lut_adj_595.init = 16'hf0f2;
    LUT4 i3913_2_lut (.A(continue_txn), .B(rst_reg_n), .Z(n6071)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i3913_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_596 (.A(n32715), .B(n32714), .C(n28419), 
         .D(n32537), .Z(addr_in[24])) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(95[18] 98[33])
    defparam i1_2_lut_3_lut_4_lut_adj_596.init = 16'hb0f0;
    LUT4 i5572_4_lut (.A(n32648), .B(continue_txn_N_2131), .C(continue_txn), 
         .D(data_stall_N_2158), .Z(clk_c_enable_118)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(198[22] 203[16])
    defparam i5572_4_lut.init = 16'h05c5;
    LUT4 data_ready_N_2113_I_0_4_lut (.A(data_ready_N_2113), .B(n32711), 
         .C(n32712), .D(mem_data_ready), .Z(continue_txn_N_2131)) /* synthesis lut_function=(!((B (C)+!B (C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(194[30:139])
    defparam data_ready_N_2113_I_0_4_lut.init = 16'h0a2a;
    LUT4 continue_txn_I_189_4_lut (.A(n29319), .B(data_ready_N_2108), .C(n32788), 
         .D(data_txn_len[1]), .Z(data_stall_N_2158)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(190[21] 191[76])
    defparam continue_txn_I_189_4_lut.init = 16'hecce;
    LUT4 i1_3_lut_adj_597 (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(data_txn_len[0]), .Z(n29319)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut_adj_597.init = 16'h4848;
    LUT4 equal_58_i1_4_lut (.A(qspi_data_byte_idx[0]), .B(instr_active), 
         .C(start_instr), .D(data_txn_len[0]), .Z(n1)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(155[21:50])
    defparam equal_58_i1_4_lut.init = 16'h5556;
    LUT4 i15783_2_lut_rep_633_3_lut_4_lut_3_lut_4_lut_4_lut (.A(n32771), .B(n32801), 
         .C(n32715), .D(n21414), .Z(n32648)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i15783_2_lut_rep_633_3_lut_4_lut_3_lut_4_lut_4_lut.init = 16'hfefa;
    LUT4 i15652_2_lut_rep_654_3_lut_4_lut_4_lut (.A(n32771), .B(n32801), 
         .C(n32715), .D(n21414), .Z(n32669)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i15652_2_lut_rep_654_3_lut_4_lut_4_lut.init = 16'hfeff;
    LUT4 i2_2_lut_rep_674_4_lut (.A(n32771), .B(n21414), .C(n32801), .D(n32715), 
         .Z(n32689)) /* synthesis lut_function=(A (D)+!A (((D)+!C)+!B)) */ ;
    defparam i2_2_lut_rep_674_4_lut.init = 16'hff15;
    LUT4 i5562_2_lut_rep_671_3_lut_4_lut (.A(n32755), .B(qspi_write_done), 
         .C(n21414), .D(n32771), .Z(n32686)) /* synthesis lut_function=(A+(B+!(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(75[13:41])
    defparam i5562_2_lut_rep_671_3_lut_4_lut.init = 16'heeef;
    LUT4 i15589_2_lut_rep_672_3_lut_4_lut (.A(n32755), .B(qspi_write_done), 
         .C(n21414), .D(n32771), .Z(n32687)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(75[13:41])
    defparam i15589_2_lut_rep_672_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\addr[23] ), .D(\addr[24] ), .Z(spi_ram_b_select_N_2313)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_2_lut_4_lut_3_lut_4_lut.init = 16'hefff;
    LUT4 i26976_2_lut_3_lut_4_lut (.A(n32755), .B(qspi_write_done), .C(instr_fetch_running), 
         .D(n32714), .Z(n29618)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(75[13:41])
    defparam i26976_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 data_addr_24__I_0_i7_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[5] ), .D(\addr[6] ), .Z(addr_in[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i13_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[11] ), .D(\addr[12] ), .Z(addr_in[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i16_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[14] ), .D(\addr[15] ), .Z(addr_in[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i11_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[9] ), .D(\addr[10] ), .Z(addr_in[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr_23__N_318[15] ), 
         .D(\addr[16] ), .Z(n3)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i18_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[16] ), .D(\addr[17] ), .Z(addr_in[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i19_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[17] ), .D(\addr[18] ), .Z(addr_in[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i14_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[12] ), .D(\addr[13] ), .Z(addr_in[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_583 (.A(mem_data_ready), .B(data_txn_len[1]), .Z(n32598)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_583.init = 16'h2222;
    LUT4 i1_2_lut_rep_563_3_lut (.A(mem_data_ready), .B(data_txn_len[1]), 
         .C(data_txn_len[0]), .Z(n32578)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_563_3_lut.init = 16'h2020;
    LUT4 data_addr_24__I_0_i12_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[10] ), .D(\addr[11] ), .Z(addr_in[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i15_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[13] ), .D(\addr[14] ), .Z(addr_in[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i5_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[3] ), .D(\addr[4] ), .Z(addr_in[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_598 (.A(n32715), .B(debug_stop_txn_N_2119), .C(is_writing), 
         .D(spi_clk_pos), .Z(stop_txn_now_N_2363)) /* synthesis lut_function=(A (B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(91[18] 99[12])
    defparam i1_4_lut_adj_598.init = 16'h8808;
    LUT4 data_addr_24__I_0_i24_3_lut_rep_511_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[22] ), .D(\addr[23] ), .Z(n32526)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i24_3_lut_rep_511_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i6_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[4] ), .D(\addr[5] ), .Z(addr_in[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i21_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[19] ), .D(\addr[20] ), .Z(addr_in[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_adj_599 (.A(instr_active), .B(\addr[24] ), .Z(n28419)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_599.init = 16'h4444;
    LUT4 i1_4_lut_adj_600 (.A(start_instr), .B(n32526), .C(\addr[24] ), 
         .D(instr_active), .Z(spi_ram_a_select_N_2309)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_4_lut_adj_600.init = 16'hffef;
    LUT4 data_addr_24__I_0_i20_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[18] ), .D(\addr[19] ), .Z(addr_in[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i20_3_lut_4_lut.init = 16'hf1e0;
    qspi_controller q_ctrl (.fsm_state({fsm_state}), .clk_c(clk_c), .clk_c_enable_340(clk_c_enable_340), 
            .n32524(n32524), .clk_c_enable_208(clk_c_enable_208), .clk_c_enable_66(clk_c_enable_66), 
            .is_writing(is_writing), .ram_b_block_N_2303(ram_b_block_N_2303), 
            .n29884(n29884), .\write_qspi_data_byte_idx_1__N_2021[0] (write_qspi_data_byte_idx_1__N_2021[0]), 
            .n27931(n27931), .n32681(n32681), .n32740(n32740), .qspi_data_ready(qspi_data_ready), 
            .n8177(n8177), .clk_c_enable_432(clk_c_enable_432), .qspi_data_out_3__N_5({qspi_data_out_3__N_5}), 
            .\qspi_data_in[3] (\qspi_data_in[3] ), .rst_reg_n(rst_reg_n), 
            .\qspi_data_in[2] (\qspi_data_in[2] ), .n32755(n32755), .n32534(n32534), 
            .\addr_in[11] (addr_in[11]), .\addr_in[10] (addr_in[10]), .\addr_in[9] (addr_in[9]), 
            .\read_cycles_count[1] (\read_cycles_count[1] ), .\addr_in[8] (addr_in[8]), 
            .spi_clk_pos(spi_clk_pos), .n32778(n32778), .\addr_in[7] (addr_in[7]), 
            .\addr_in[4] (addr_in[4]), .data_req_N_2334(data_req_N_2334), 
            .\addr_in[5] (addr_in[5]), .\addr_in[6] (addr_in[6]), .\addr_in[12] (addr_in[12]), 
            .\addr_in[13] (addr_in[13]), .\addr_in[14] (addr_in[14]), .\addr_in[15] (addr_in[15]), 
            .\instr_data[8] (instr_data[8]), .qspi_ram_a_select(qspi_ram_a_select), 
            .last_ram_b_sel(last_ram_b_sel), .qspi_ram_b_select(qspi_ram_b_select), 
            .clk_N_45(clk_N_45), .n31475(n31475), .n3(n3), .stop_txn_reg(stop_txn_reg), 
            .ram_a_block_N_2299(ram_a_block_N_2299), .n32521(n32521), .\addr_in[17] (addr_in[17]), 
            .\qspi_data_oe[1] (\qspi_data_oe[1] ), .clk_c_enable_341(clk_c_enable_341), 
            .n1072(n1072), .\addr_in[18] (addr_in[18]), .\addr_in[19] (addr_in[19]), 
            .\addr_in[20] (addr_in[20]), .\addr_in[21] (addr_in[21]), .n29752(n29752), 
            .\addr_in[22] (addr_in[22]), .n32526(n32526), .\addr[24] (\addr[24] ), 
            .n34272(n34272), .\instr_data[9] (instr_data[9]), .n29771(n29771), 
            .\instr_data[10] (instr_data[10]), .n29774(n29774), .n19867(n19867), 
            .data_stall(data_stall), .n482(n482), .qspi_write_done(qspi_write_done), 
            .n32715(n32715), .clk_c_enable_488(clk_c_enable_488), .\addr_23__N_2188[0] (addr_23__N_2188[0]), 
            .debug_stop_txn(debug_stop_txn), .clk_c_enable_31(clk_c_enable_31), 
            .\writing_N_164[3] (\writing_N_164[3] ), .n32542(n32542), .data_ready_N_2347(data_ready_N_2347), 
            .n29767(n29767), .n29770(n29770), .n29773(n29773), .\instr_data[11] (instr_data[11]), 
            .n29776(n29776), .n4513(n4513), .\instr_data[13] (instr_data[13]), 
            .\instr_data[14] (instr_data[14]), .n4501(n4501), .n32833(n32833), 
            .n26811(n26811), .\instr_data[12] (instr_data[12]), .n4503(n4503), 
            .\addr[20] (\addr[20]_adj_15 ), .\addr[22] (\addr[22]_adj_16 ), 
            .n11756(n11756), .\addr_in[3] (addr_in[3]), .\addr_in[2] (addr_in[2]), 
            .\addr_in[1] (addr_in[1]), .\instr_data[15] (instr_data[15]), 
            .\qspi_data_byte_idx[1] (qspi_data_byte_idx[1]), .n6704(n6704), 
            .n6218(n6218), .\addr_in[24] (addr_in[24]), .n8205(n8205), 
            .start_instr(start_instr), .instr_active(instr_active), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .qspi_clk_N_56(qspi_clk_N_56), .n11684(n11684), .n32712(n32712), 
            .n32686(n32686), .n11193(n11193), .n32522(n32522), .n6220(n6220), 
            .n31866(n31866), .clk_c_enable_543(clk_c_enable_543), .spi_ram_a_select_N_2309(spi_ram_a_select_N_2309), 
            .n28319(n28319), .spi_ram_b_select_N_2313(spi_ram_b_select_N_2313), 
            .n32874(n32874), .stop_txn_now_N_2363(stop_txn_now_N_2363), 
            .n28259(n28259), .n29768(n29768), .n29777(n29777), .\qspi_data_in[0] (\qspi_data_in[0] ), 
            .n332(n332), .n32060(n32060), .debug_stop_txn_N_2119(debug_stop_txn_N_2119), 
            .n31677(n31677), .n29755(n29755), .n31646(n31646), .n29761(n29761), 
            .n31639(n31639), .n29764(n29764), .n28111(n28111), .n32523(n32523), 
            .n32789(n32789), .n32892(n32892)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(112[21] 136[6])
    
endmodule
//
// Verilog Description of module qspi_controller
//

module qspi_controller (fsm_state, clk_c, clk_c_enable_340, n32524, 
            clk_c_enable_208, clk_c_enable_66, is_writing, ram_b_block_N_2303, 
            n29884, \write_qspi_data_byte_idx_1__N_2021[0] , n27931, n32681, 
            n32740, qspi_data_ready, n8177, clk_c_enable_432, qspi_data_out_3__N_5, 
            \qspi_data_in[3] , rst_reg_n, \qspi_data_in[2] , n32755, 
            n32534, \addr_in[11] , \addr_in[10] , \addr_in[9] , \read_cycles_count[1] , 
            \addr_in[8] , spi_clk_pos, n32778, \addr_in[7] , \addr_in[4] , 
            data_req_N_2334, \addr_in[5] , \addr_in[6] , \addr_in[12] , 
            \addr_in[13] , \addr_in[14] , \addr_in[15] , \instr_data[8] , 
            qspi_ram_a_select, last_ram_b_sel, qspi_ram_b_select, clk_N_45, 
            n31475, n3, stop_txn_reg, ram_a_block_N_2299, n32521, 
            \addr_in[17] , \qspi_data_oe[1] , clk_c_enable_341, n1072, 
            \addr_in[18] , \addr_in[19] , \addr_in[20] , \addr_in[21] , 
            n29752, \addr_in[22] , n32526, \addr[24] , n34272, \instr_data[9] , 
            n29771, \instr_data[10] , n29774, n19867, data_stall, 
            n482, qspi_write_done, n32715, clk_c_enable_488, \addr_23__N_2188[0] , 
            debug_stop_txn, clk_c_enable_31, \writing_N_164[3] , n32542, 
            data_ready_N_2347, n29767, n29770, n29773, \instr_data[11] , 
            n29776, n4513, \instr_data[13] , \instr_data[14] , n4501, 
            n32833, n26811, \instr_data[12] , n4503, \addr[20] , \addr[22] , 
            n11756, \addr_in[3] , \addr_in[2] , \addr_in[1] , \instr_data[15] , 
            \qspi_data_byte_idx[1] , n6704, n6218, \addr_in[24] , n8205, 
            start_instr, instr_active, spi_clk_pos_derived_59, qspi_clk_N_56, 
            n11684, n32712, n32686, n11193, n32522, n6220, n31866, 
            clk_c_enable_543, spi_ram_a_select_N_2309, n28319, spi_ram_b_select_N_2313, 
            n32874, stop_txn_now_N_2363, n28259, n29768, n29777, \qspi_data_in[0] , 
            n332, n32060, debug_stop_txn_N_2119, n31677, n29755, n31646, 
            n29761, n31639, n29764, n28111, n32523, n32789, n32892) /* synthesis syn_module_defined=1 */ ;
    output [2:0]fsm_state;
    input clk_c;
    input clk_c_enable_340;
    input n32524;
    input clk_c_enable_208;
    input clk_c_enable_66;
    output is_writing;
    input ram_b_block_N_2303;
    input n29884;
    output \write_qspi_data_byte_idx_1__N_2021[0] ;
    input n27931;
    output n32681;
    output n32740;
    output qspi_data_ready;
    input n8177;
    input clk_c_enable_432;
    input [3:0]qspi_data_out_3__N_5;
    input \qspi_data_in[3] ;
    input rst_reg_n;
    input \qspi_data_in[2] ;
    output n32755;
    input n32534;
    input \addr_in[11] ;
    input \addr_in[10] ;
    input \addr_in[9] ;
    output \read_cycles_count[1] ;
    input \addr_in[8] ;
    output spi_clk_pos;
    output n32778;
    input \addr_in[7] ;
    input \addr_in[4] ;
    output data_req_N_2334;
    input \addr_in[5] ;
    input \addr_in[6] ;
    input \addr_in[12] ;
    input \addr_in[13] ;
    input \addr_in[14] ;
    input \addr_in[15] ;
    output \instr_data[8] ;
    output qspi_ram_a_select;
    output last_ram_b_sel;
    output qspi_ram_b_select;
    input clk_N_45;
    input n31475;
    input n3;
    output stop_txn_reg;
    output ram_a_block_N_2299;
    output n32521;
    input \addr_in[17] ;
    output \qspi_data_oe[1] ;
    input clk_c_enable_341;
    output n1072;
    input \addr_in[18] ;
    input \addr_in[19] ;
    input \addr_in[20] ;
    input \addr_in[21] ;
    input n29752;
    input \addr_in[22] ;
    input n32526;
    input \addr[24] ;
    input n34272;
    output \instr_data[9] ;
    input n29771;
    output \instr_data[10] ;
    input n29774;
    input n19867;
    input data_stall;
    output n482;
    input qspi_write_done;
    output n32715;
    input clk_c_enable_488;
    input \addr_23__N_2188[0] ;
    output debug_stop_txn;
    output clk_c_enable_31;
    output \writing_N_164[3] ;
    input n32542;
    input data_ready_N_2347;
    input n29767;
    input n29770;
    input n29773;
    output \instr_data[11] ;
    input n29776;
    output n4513;
    output \instr_data[13] ;
    output \instr_data[14] ;
    output n4501;
    output n32833;
    output n26811;
    output \instr_data[12] ;
    output n4503;
    output \addr[20] ;
    output \addr[22] ;
    input n11756;
    input \addr_in[3] ;
    input \addr_in[2] ;
    input \addr_in[1] ;
    output \instr_data[15] ;
    input \qspi_data_byte_idx[1] ;
    input n6704;
    output n6218;
    input \addr_in[24] ;
    output n8205;
    input start_instr;
    input instr_active;
    output spi_clk_pos_derived_59;
    output qspi_clk_N_56;
    output n11684;
    input n32712;
    input n32686;
    output n11193;
    input n32522;
    output n6220;
    input n31866;
    input clk_c_enable_543;
    input spi_ram_a_select_N_2309;
    output n28319;
    input spi_ram_b_select_N_2313;
    output n32874;
    input stop_txn_now_N_2363;
    input n28259;
    input n29768;
    input n29777;
    input \qspi_data_in[0] ;
    input n332;
    output n32060;
    input debug_stop_txn_N_2119;
    input n31677;
    input n29755;
    input n31646;
    input n29761;
    input n31639;
    input n29764;
    output n28111;
    input n32523;
    input n32789;
    output n32892;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    
    wire n1055;
    wire [1:0]read_cycles_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(105[15:32])
    wire [1:0]n396;
    wire [55:0]instr_data_15__N_1959;
    wire [7:0]data_out_7__N_2273;
    
    wire n30226;
    wire [7:0]data_out_7__N_2177;
    wire [2:0]nibbles_remaining;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(86[15:32])
    
    wire n1064, data_req_N_2318, n11068, n18383;
    wire [1:0]delay_cycles_cfg;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(87[15:31])
    
    wire n27898, n27342, n32743, n27343, n32888;
    wire [0:0]n5188;
    
    wire n32887, n26814, n32891, n32890, data_ready_N_2338, n32709;
    wire [3:0]spi_in_buffer;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(91[15:28])
    
    wire n31636, n31643;
    wire [23:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(84[31:35])
    wire [23:0]addr_23__N_2188;
    
    wire n86, n32536, n1164;
    wire [1:0]n381;
    
    wire n32775, n32739, n32752, n32777, n32744, n17865;
    wire [2:0]n4330;
    
    wire n32817, n30110, n26894, n32782, n31476, n31473, clk_c_enable_456, 
        clk_c_enable_507, last_ram_a_sel, spi_clk_neg, n31474, n32674, 
        spi_clk_use_neg, stop_txn_reg_N_2360, n1057, n1056, n31472, 
        n32830, n1042, n32667, clk_c_enable_438, n27903, n29375, 
        n10820, n32823, n32722, n32753, n32820;
    wire [1:0]n127;
    wire [1:0]n333;
    wire [1:0]n181;
    
    wire n29577;
    wire [0:0]n5181;
    wire [3:0]n4499;
    
    wire clk_c_enable_511, n6216;
    wire [2:0]n356;
    
    wire n17882, n28149;
    wire [2:0]n312;
    
    wire n32713, n10, n32059, n31674, n32696, n31645, n31638, 
        n31678, n31675, n31676, n32856, n6, n32857, n31647, n31644, 
        n31640, n31637, n32855;
    
    FD1P3IX fsm_state__i0 (.D(n1055), .SP(clk_c_enable_340), .CD(n32524), 
            .CK(clk_c), .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i0.GSR = "DISABLED";
    FD1P3IX read_cycles_count__i0 (.D(n396[0]), .SP(clk_c_enable_208), .CD(n32524), 
            .CK(clk_c), .Q(read_cycles_count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam read_cycles_count__i0.GSR = "DISABLED";
    PFUMX data_out_7__I_0_242_i8 (.BLUT(instr_data_15__N_1959[31]), .ALUT(data_out_7__N_2273[7]), 
          .C0(n30226), .Z(data_out_7__N_2177[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i7 (.BLUT(instr_data_15__N_1959[30]), .ALUT(data_out_7__N_2273[6]), 
          .C0(n30226), .Z(data_out_7__N_2177[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i6 (.BLUT(instr_data_15__N_1959[29]), .ALUT(data_out_7__N_2273[5]), 
          .C0(n30226), .Z(data_out_7__N_2177[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i5 (.BLUT(instr_data_15__N_1959[28]), .ALUT(data_out_7__N_2273[4]), 
          .C0(n30226), .Z(data_out_7__N_2177[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    FD1P3IX nibbles_remaining__i0 (.D(n1064), .SP(clk_c_enable_66), .CD(n32524), 
            .CK(clk_c), .Q(nibbles_remaining[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i0.GSR = "DISABLED";
    FD1P3IX is_writing_222 (.D(n29884), .SP(ram_b_block_N_2303), .CD(n32524), 
            .CK(clk_c), .Q(is_writing)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam is_writing_222.GSR = "DISABLED";
    FD1S3IX data_req_230 (.D(data_req_N_2318), .CK(clk_c), .CD(n27931), 
            .Q(\write_qspi_data_byte_idx_1__N_2021[0] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam data_req_230.GSR = "DISABLED";
    FD1P3IX nibbles_remaining__i2 (.D(n11068), .SP(clk_c_enable_66), .CD(n32524), 
            .CK(clk_c), .Q(nibbles_remaining[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i2.GSR = "DISABLED";
    FD1P3IX nibbles_remaining__i1 (.D(n18383), .SP(clk_c_enable_66), .CD(n32524), 
            .CK(clk_c), .Q(nibbles_remaining[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i1.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(delay_cycles_cfg[0]), 
         .D(fsm_state[1]), .Z(n27898)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h0020;
    LUT4 i1_4_lut (.A(n32681), .B(n27342), .C(n32743), .D(n32740), .Z(n27343)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut.init = 16'hff7f;
    LUT4 mux_2865_i2_4_lut_then_1_lut (.A(nibbles_remaining[1]), .Z(n32888)) /* synthesis lut_function=(A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_2865_i2_4_lut_then_1_lut.init = 16'haaaa;
    LUT4 mux_2865_i2_4_lut_else_1_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(n5188[0]), .D(fsm_state[0]), .Z(n32887)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_2865_i2_4_lut_else_1_lut.init = 16'h2220;
    LUT4 i1_4_lut_then_3_lut (.A(fsm_state[1]), .B(n26814), .C(fsm_state[2]), 
         .Z(n32891)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(209[30] 211[24])
    defparam i1_4_lut_then_3_lut.init = 16'h0808;
    LUT4 i1_4_lut_else_3_lut (.A(fsm_state[1]), .B(n26814), .C(fsm_state[2]), 
         .D(fsm_state[0]), .Z(n32890)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(209[30] 211[24])
    defparam i1_4_lut_else_3_lut.init = 16'h0800;
    FD1S3IX data_ready_224 (.D(data_ready_N_2338), .CK(clk_c), .CD(n8177), 
            .Q(qspi_data_ready)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam data_ready_224.GSR = "DISABLED";
    FD1P3AX delay_cycles_cfg_i0_i0 (.D(qspi_data_out_3__N_5[0]), .SP(clk_c_enable_432), 
            .CK(clk_c), .Q(delay_cycles_cfg[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(112[12] 117[8])
    defparam delay_cycles_cfg_i0_i0.GSR = "DISABLED";
    LUT4 n9_bdd_4_lut_28791 (.A(n32709), .B(\qspi_data_in[3] ), .C(spi_in_buffer[3]), 
         .D(rst_reg_n), .Z(n31636)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam n9_bdd_4_lut_28791.init = 16'he4a0;
    LUT4 n9_bdd_4_lut_29238 (.A(n32709), .B(\qspi_data_in[2] ), .C(spi_in_buffer[2]), 
         .D(rst_reg_n), .Z(n31643)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam n9_bdd_4_lut_29238.init = 16'he4a0;
    LUT4 addr_23__I_0_i12_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[11] ), 
         .D(addr[7]), .Z(addr_23__N_2188[11])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i11_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[10] ), 
         .D(addr[6]), .Z(addr_23__N_2188[10])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i10_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[9] ), 
         .D(addr[5]), .Z(addr_23__N_2188[9])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 fsm_state_2__bdd_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(fsm_state[0]), 
         .Z(n86)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam fsm_state_2__bdd_3_lut.init = 16'h0202;
    LUT4 mux_114_i1_4_lut_4_lut (.A(read_cycles_count[0]), .B(n32536), .C(n1164), 
         .D(n27898), .Z(n381[0])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam mux_114_i1_4_lut_4_lut.init = 16'h5f5c;
    LUT4 i1_2_lut_rep_760 (.A(fsm_state[1]), .B(fsm_state[0]), .Z(n32775)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_760.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_724_3_lut (.A(fsm_state[1]), .B(fsm_state[0]), .C(fsm_state[2]), 
         .Z(n32739)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_724_3_lut.init = 16'hbfbf;
    FD1P3IX read_cycles_count__i1 (.D(n396[1]), .SP(clk_c_enable_208), .CD(n32524), 
            .CK(clk_c), .Q(\read_cycles_count[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam read_cycles_count__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_737_3_lut (.A(fsm_state[1]), .B(fsm_state[0]), .C(fsm_state[2]), 
         .Z(n32752)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_737_3_lut.init = 16'hfbfb;
    LUT4 i14865_2_lut_rep_762 (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .Z(n32777)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14865_2_lut_rep_762.init = 16'heeee;
    LUT4 i1_3_lut_rep_729_4_lut (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .C(fsm_state[0]), .D(fsm_state[2]), .Z(n32744)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_3_lut_rep_729_4_lut.init = 16'hefff;
    LUT4 addr_23__I_0_i9_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[8] ), 
         .D(addr[4]), .Z(addr_23__N_2188[8])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i9_3_lut_4_lut.init = 16'hfb40;
    LUT4 i27_3_lut_4_lut (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .C(n17865), .D(spi_clk_pos), .Z(n32681)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam i27_3_lut_4_lut.init = 16'hf101;
    LUT4 equal_121_i4_2_lut_rep_763 (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .Z(n32778)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam equal_121_i4_2_lut_rep_763.init = 16'heeee;
    LUT4 equal_121_i5_2_lut_rep_725_3_lut (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .C(nibbles_remaining[0]), .Z(n32740)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam equal_121_i5_2_lut_rep_725_3_lut.init = 16'hfefe;
    LUT4 mux_2865_i3_3_lut_4_lut_4_lut (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .C(n32752), .D(nibbles_remaining[0]), .Z(n4330[2])) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam mux_2865_i3_3_lut_4_lut_4_lut.init = 16'hcccd;
    LUT4 i28583_2_lut_3_lut_4_lut (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .C(n32817), .D(nibbles_remaining[0]), .Z(n30110)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i28583_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .C(n4330[1]), .D(nibbles_remaining[0]), .Z(n26894)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 addr_23__I_0_i8_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[7] ), 
         .D(addr[3]), .Z(addr_23__N_2188[7])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15436_2_lut_rep_767 (.A(fsm_state[2]), .B(fsm_state[1]), .Z(n32782)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15436_2_lut_rep_767.init = 16'h8888;
    L6MUX21 i28698 (.D0(n31476), .D1(n31473), .SD(n30226), .Z(data_out_7__N_2177[0]));
    LUT4 i1_2_lut_rep_728_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(fsm_state[0]), 
         .Z(n32743)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_728_3_lut.init = 16'hf7f7;
    LUT4 addr_23__I_0_i5_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[4] ), 
         .D(addr[0]), .Z(addr_23__N_2188[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 i15717_2_lut_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(fsm_state[0]), 
         .Z(data_req_N_2334)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15717_2_lut_3_lut.init = 16'h8080;
    LUT4 addr_23__I_0_i6_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[5] ), 
         .D(addr[1]), .Z(addr_23__N_2188[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i7_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[6] ), 
         .D(addr[2]), .Z(addr_23__N_2188[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i7_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX spi_in_buffer_i0_i0 (.D(qspi_data_out_3__N_5[0]), .SP(clk_c_enable_456), 
            .CK(clk_c), .Q(spi_in_buffer[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i0.GSR = "DISABLED";
    LUT4 addr_23__I_0_i13_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[12] ), 
         .D(addr[8]), .Z(addr_23__N_2188[12])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i14_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[13] ), 
         .D(addr[9]), .Z(addr_23__N_2188[13])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i15_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[14] ), 
         .D(addr[10]), .Z(addr_23__N_2188[14])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i16_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[15] ), 
         .D(addr[11]), .Z(addr_23__N_2188[15])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i16_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX data_i1 (.D(data_out_7__N_2177[0]), .SP(clk_c_enable_507), .CK(clk_c), 
            .Q(\instr_data[8] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i1.GSR = "DISABLED";
    FD1S3JX last_ram_a_sel_235 (.D(qspi_ram_a_select), .CK(clk_c), .PD(clk_c_enable_432), 
            .Q(last_ram_a_sel)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(272[12] 280[8])
    defparam last_ram_a_sel_235.GSR = "DISABLED";
    FD1S3JX last_ram_b_sel_236 (.D(qspi_ram_b_select), .CK(clk_c), .PD(clk_c_enable_432), 
            .Q(last_ram_b_sel)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(272[12] 280[8])
    defparam last_ram_b_sel_236.GSR = "DISABLED";
    FD1S3AX spi_clk_neg_237 (.D(spi_clk_pos), .CK(clk_N_45), .Q(spi_clk_neg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(286[12:54])
    defparam spi_clk_neg_237.GSR = "DISABLED";
    PFUMX i28696 (.BLUT(n31475), .ALUT(n31474), .C0(n32674), .Z(n31476));
    FD1P3AX spi_clk_use_neg_220 (.D(qspi_data_out_3__N_5[2]), .SP(clk_c_enable_432), 
            .CK(clk_c), .Q(spi_clk_use_neg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(112[12] 117[8])
    defparam spi_clk_use_neg_220.GSR = "DISABLED";
    LUT4 i8_3_lut_4_lut (.A(n32755), .B(n32534), .C(n3), .D(addr[12]), 
         .Z(addr_23__N_2188[16])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam i8_3_lut_4_lut.init = 16'hfb40;
    FD1S3IX stop_txn_reg_218 (.D(stop_txn_reg_N_2360), .CK(clk_c), .CD(clk_c_enable_432), 
            .Q(stop_txn_reg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(98[12] 103[8])
    defparam stop_txn_reg_218.GSR = "DISABLED";
    LUT4 i7180_rep_506_3_lut_4_lut (.A(ram_a_block_N_2299), .B(n32534), 
         .C(n32755), .D(ram_b_block_N_2303), .Z(n32521)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i7180_rep_506_3_lut_4_lut.init = 16'h0800;
    LUT4 addr_23__I_0_i18_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[17] ), 
         .D(addr[13]), .Z(addr_23__N_2188[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i18_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX fsm_state__i2 (.D(n1057), .SP(clk_c_enable_340), .CD(n32524), 
            .CK(clk_c), .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1P3IX fsm_state__i1 (.D(n1056), .SP(clk_c_enable_340), .CD(n32524), 
            .CK(clk_c), .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i1.GSR = "DISABLED";
    FD1P3IX spi_data_oe__i1 (.D(n1072), .SP(clk_c_enable_341), .CD(n32524), 
            .CK(clk_c), .Q(\qspi_data_oe[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_data_oe__i1.GSR = "DISABLED";
    LUT4 addr_23__I_0_i19_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[18] ), 
         .D(addr[14]), .Z(addr_23__N_2188[18])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i20_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[19] ), 
         .D(addr[15]), .Z(addr_23__N_2188[19])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i21_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[20] ), 
         .D(addr[16]), .Z(addr_23__N_2188[20])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i22_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[21] ), 
         .D(addr[17]), .Z(addr_23__N_2188[21])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i22_3_lut_4_lut.init = 16'hfb40;
    PFUMX i28693 (.BLUT(n29752), .ALUT(n31472), .C0(n32830), .Z(n31473));
    LUT4 addr_23__I_0_i23_3_lut_4_lut (.A(n32755), .B(n32534), .C(\addr_in[22] ), 
         .D(addr[18]), .Z(addr_23__N_2188[22])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i23_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i24_3_lut_4_lut (.A(n32755), .B(n32534), .C(n32526), 
         .D(addr[19]), .Z(addr_23__N_2188[23])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i24_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_699_i2_3_lut_4_lut (.A(\addr[24] ), .B(n34272), .C(n1072), 
         .D(n1042), .Z(n1056)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;
    defparam mux_699_i2_3_lut_4_lut.init = 16'hdfd0;
    FD1P3AX delay_cycles_cfg_i0_i1 (.D(qspi_data_out_3__N_5[1]), .SP(clk_c_enable_432), 
            .CK(clk_c), .Q(delay_cycles_cfg[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(112[12] 117[8])
    defparam delay_cycles_cfg_i0_i1.GSR = "DISABLED";
    LUT4 i27970_3_lut_4_lut (.A(\instr_data[9] ), .B(n32667), .C(n32674), 
         .D(n29771), .Z(instr_data_15__N_1959[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(231[22] 237[16])
    defparam i27970_3_lut_4_lut.init = 16'h8f80;
    LUT4 i27972_3_lut_4_lut (.A(\instr_data[10] ), .B(n32667), .C(n32674), 
         .D(n29774), .Z(instr_data_15__N_1959[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(231[22] 237[16])
    defparam i27972_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_rep_802 (.A(fsm_state[2]), .B(fsm_state[0]), .Z(n32817)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_802.init = 16'h8888;
    FD1P3AX spi_clk_pos_225 (.D(n27903), .SP(clk_c_enable_438), .CK(clk_c), 
            .Q(spi_clk_pos)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_clk_pos_225.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_521_3_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), 
         .C(n19867), .D(data_stall), .Z(n32536)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_2_lut_rep_521_3_lut_4_lut.init = 16'h8880;
    LUT4 i1_3_lut_3_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(fsm_state[1]), 
         .Z(n29375)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)+!B !(C)))) */ ;
    defparam i1_3_lut_3_lut.init = 16'h3434;
    LUT4 i1_2_lut_3_lut_4_lut_3_lut (.A(fsm_state[2]), .B(fsm_state[0]), 
         .C(fsm_state[1]), .Z(n10820)) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_3_lut.init = 16'h7373;
    LUT4 i794_2_lut_rep_707_3_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(n32823), .D(fsm_state[0]), .Z(n32722)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(265[13:23])
    defparam i794_2_lut_rep_707_3_lut_4_lut.init = 16'hffdf;
    LUT4 fsm_state_2__I_0_239_i5_2_lut_rep_738_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(fsm_state[0]), .Z(n32753)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(265[13:23])
    defparam fsm_state_2__I_0_239_i5_2_lut_rep_738_3_lut.init = 16'hfdfd;
    LUT4 i171_2_lut_3_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(spi_clk_pos), 
         .D(fsm_state[0]), .Z(n482)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(265[13:23])
    defparam i171_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_805 (.A(fsm_state[1]), .B(fsm_state[0]), .Z(n32820)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(266[13:21])
    defparam i1_2_lut_rep_805.init = 16'heeee;
    LUT4 qspi_busy_I_0_2_lut_rep_700_3_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[0]), 
         .C(qspi_write_done), .D(fsm_state[2]), .Z(n32715)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(266[13:21])
    defparam qspi_busy_I_0_2_lut_rep_700_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_740_3_lut (.A(fsm_state[1]), .B(fsm_state[0]), .C(fsm_state[2]), 
         .Z(n32755)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(266[13:21])
    defparam i1_2_lut_rep_740_3_lut.init = 16'hfefe;
    FD1P3AX addr_i0 (.D(\addr_23__N_2188[0] ), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(fsm_state[2]), .B(n32820), .C(rst_reg_n), 
         .D(debug_stop_txn), .Z(clk_c_enable_31)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_3_lut_4_lut.init = 16'hff1f;
    LUT4 i15254_2_lut_rep_808 (.A(\writing_N_164[3] ), .B(is_writing), .Z(n32823)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15254_2_lut_rep_808.init = 16'heeee;
    LUT4 i15810_2_lut (.A(read_cycles_count[0]), .B(\read_cycles_count[1] ), 
         .Z(n127[1])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(151[22:69])
    defparam i15810_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_577 (.A(delay_cycles_cfg[1]), .B(n86), .C(n32542), 
         .D(n32817), .Z(n333[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(264[13:21])
    defparam i1_4_lut_adj_577.init = 16'ha088;
    FD1P3AX spi_in_buffer_i0_i1 (.D(qspi_data_out_3__N_5[1]), .SP(clk_c_enable_456), 
            .CK(clk_c), .Q(spi_in_buffer[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i1.GSR = "DISABLED";
    LUT4 i10703_1_lut_rep_815 (.A(is_writing), .Z(n32830)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i10703_1_lut_rep_815.init = 16'h5555;
    LUT4 mux_60_i1_4_lut_4_lut_4_lut (.A(is_writing), .B(data_ready_N_2347), 
         .C(delay_cycles_cfg[0]), .D(read_cycles_count[0]), .Z(n181[0])) /* synthesis lut_function=(!(A (B+(D))+!A !(B (C)+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_60_i1_4_lut_4_lut_4_lut.init = 16'h4073;
    LUT4 mux_180_i5_3_lut_3_lut (.A(is_writing), .B(\instr_data[8] ), .C(n29767), 
         .Z(data_out_7__N_2273[4])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i5_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_4_lut_4_lut (.A(is_writing), .B(n29577), .C(fsm_state[0]), 
         .D(read_cycles_count[0]), .Z(clk_c_enable_456)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_4_lut_4_lut.init = 16'h0004;
    LUT4 i15220_2_lut_2_lut (.A(is_writing), .B(\writing_N_164[3] ), .Z(n5188[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i15220_2_lut_2_lut.init = 16'h4444;
    LUT4 mux_180_i6_3_lut_3_lut (.A(is_writing), .B(\instr_data[9] ), .C(n29770), 
         .Z(data_out_7__N_2273[5])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i6_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i7_3_lut_3_lut (.A(is_writing), .B(\instr_data[10] ), .C(n29773), 
         .Z(data_out_7__N_2273[6])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i7_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i8_3_lut_3_lut (.A(is_writing), .B(\instr_data[11] ), .C(n29776), 
         .Z(data_out_7__N_2273[7])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i8_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_2_lut (.A(is_writing), .B(delay_cycles_cfg[1]), .Z(n5181[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 mux_2897_i2_3_lut (.A(addr[21]), .B(n4499[1]), .C(fsm_state[0]), 
         .Z(n4513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2897_i2_3_lut.init = 16'hcaca;
    LUT4 mux_2890_i2_4_lut (.A(nibbles_remaining[0]), .B(\instr_data[13] ), 
         .C(fsm_state[2]), .D(is_writing), .Z(n4499[1])) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B+!(C (D)))) */ ;
    defparam mux_2890_i2_4_lut.init = 16'hc5f5;
    LUT4 i15378_3_lut (.A(\instr_data[14] ), .B(fsm_state[2]), .C(is_writing), 
         .Z(n4501)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i15378_3_lut.init = 16'h8c8c;
    FD1P3AX spi_in_buffer_i0_i2 (.D(qspi_data_out_3__N_5[2]), .SP(clk_c_enable_456), 
            .CK(clk_c), .Q(spi_in_buffer[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX spi_in_buffer_i0_i3 (.D(qspi_data_out_3__N_5[3]), .SP(clk_c_enable_456), 
            .CK(clk_c), .Q(spi_in_buffer[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i3.GSR = "DISABLED";
    LUT4 i13_3_lut_rep_818 (.A(fsm_state[2]), .B(fsm_state[0]), .C(fsm_state[1]), 
         .Z(n32833)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam i13_3_lut_rep_818.init = 16'h1c1c;
    LUT4 i1_2_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(fsm_state[1]), 
         .D(\qspi_data_oe[1] ), .Z(n26811)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C (D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h1c00;
    LUT4 mux_2890_i1_4_lut_4_lut (.A(nibbles_remaining[0]), .B(is_writing), 
         .C(fsm_state[2]), .D(\instr_data[12] ), .Z(n4503)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A ((C (D))+!B)) */ ;
    defparam mux_2890_i1_4_lut_4_lut.init = 16'hf131;
    FD1P3AX addr_i4 (.D(addr_23__N_2188[4]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i4.GSR = "DISABLED";
    FD1P3AX addr_i5 (.D(addr_23__N_2188[5]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i5.GSR = "DISABLED";
    FD1P3AX addr_i6 (.D(addr_23__N_2188[6]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i6.GSR = "DISABLED";
    FD1P3AX addr_i7 (.D(addr_23__N_2188[7]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i7.GSR = "DISABLED";
    FD1P3AX addr_i8 (.D(addr_23__N_2188[8]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i8.GSR = "DISABLED";
    FD1P3AX addr_i9 (.D(addr_23__N_2188[9]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i9.GSR = "DISABLED";
    FD1P3AX addr_i10 (.D(addr_23__N_2188[10]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i10.GSR = "DISABLED";
    FD1P3AX addr_i11 (.D(addr_23__N_2188[11]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i11.GSR = "DISABLED";
    FD1P3AX addr_i12 (.D(addr_23__N_2188[12]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i12.GSR = "DISABLED";
    FD1P3AX addr_i13 (.D(addr_23__N_2188[13]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i13.GSR = "DISABLED";
    FD1P3AX addr_i14 (.D(addr_23__N_2188[14]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i14.GSR = "DISABLED";
    FD1P3AX addr_i15 (.D(addr_23__N_2188[15]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i15.GSR = "DISABLED";
    FD1P3AX addr_i16 (.D(addr_23__N_2188[16]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i16.GSR = "DISABLED";
    FD1P3AX addr_i17 (.D(addr_23__N_2188[17]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i17.GSR = "DISABLED";
    FD1P3AX addr_i18 (.D(addr_23__N_2188[18]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i18.GSR = "DISABLED";
    FD1P3AX addr_i19 (.D(addr_23__N_2188[19]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i19.GSR = "DISABLED";
    FD1P3AX addr_i20 (.D(addr_23__N_2188[20]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(\addr[20] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i20.GSR = "DISABLED";
    FD1P3AX addr_i21 (.D(addr_23__N_2188[21]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i21.GSR = "DISABLED";
    FD1P3AX addr_i22 (.D(addr_23__N_2188[22]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(\addr[22] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i22.GSR = "DISABLED";
    FD1P3AX addr_i23 (.D(addr_23__N_2188[23]), .SP(clk_c_enable_488), .CK(clk_c), 
            .Q(addr[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i23.GSR = "DISABLED";
    FD1P3AX data_i2 (.D(data_out_7__N_2177[1]), .SP(clk_c_enable_507), .CK(clk_c), 
            .Q(\instr_data[9] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i2.GSR = "DISABLED";
    FD1P3IX addr_i3 (.D(\addr_in[3] ), .SP(clk_c_enable_488), .CD(n11756), 
            .CK(clk_c), .Q(addr[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i3.GSR = "DISABLED";
    FD1P3IX addr_i2 (.D(\addr_in[2] ), .SP(clk_c_enable_488), .CD(n11756), 
            .CK(clk_c), .Q(addr[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i2.GSR = "DISABLED";
    FD1P3IX addr_i1 (.D(\addr_in[1] ), .SP(clk_c_enable_488), .CD(n11756), 
            .CK(clk_c), .Q(addr[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i1.GSR = "DISABLED";
    FD1P3AX data_i3 (.D(data_out_7__N_2177[2]), .SP(clk_c_enable_507), .CK(clk_c), 
            .Q(\instr_data[10] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i3.GSR = "DISABLED";
    FD1P3AX data_i4 (.D(data_out_7__N_2177[3]), .SP(clk_c_enable_507), .CK(clk_c), 
            .Q(\instr_data[11] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i4.GSR = "DISABLED";
    FD1P3AX data_i5 (.D(data_out_7__N_2177[4]), .SP(clk_c_enable_511), .CK(clk_c), 
            .Q(\instr_data[12] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i5.GSR = "DISABLED";
    FD1P3AX data_i6 (.D(data_out_7__N_2177[5]), .SP(clk_c_enable_511), .CK(clk_c), 
            .Q(\instr_data[13] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i6.GSR = "DISABLED";
    FD1P3AX data_i7 (.D(data_out_7__N_2177[6]), .SP(clk_c_enable_511), .CK(clk_c), 
            .Q(\instr_data[14] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i7.GSR = "DISABLED";
    FD1P3AX data_i8 (.D(data_out_7__N_2177[7]), .SP(clk_c_enable_511), .CK(clk_c), 
            .Q(\instr_data[15] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i8.GSR = "DISABLED";
    LUT4 i28544_4_lut (.A(is_writing), .B(n32674), .C(\qspi_data_byte_idx[1] ), 
         .D(n6704), .Z(n30226)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(238[18] 244[12])
    defparam i28544_4_lut.init = 16'h7557;
    LUT4 i3180_4_lut (.A(n32681), .B(n6216), .C(n32755), .D(n32743), 
         .Z(n6218)) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i3180_4_lut.init = 16'haccc;
    LUT4 mux_699_i1_4_lut (.A(n356[0]), .B(\addr_in[24] ), .C(n1072), 
         .D(n17882), .Z(n1055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam mux_699_i1_4_lut.init = 16'hcfca;
    LUT4 i28434_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n32820), .C(rst_reg_n), 
         .D(qspi_write_done), .Z(n8205)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i28434_2_lut_3_lut_4_lut.init = 16'h0f1f;
    LUT4 i1_4_lut_adj_578 (.A(ram_a_block_N_2299), .B(ram_b_block_N_2303), 
         .C(n32534), .D(n32755), .Z(n1072)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i1_4_lut_adj_578.init = 16'h0080;
    LUT4 i1_4_lut_adj_579 (.A(start_instr), .B(n32526), .C(\addr[24] ), 
         .D(n28149), .Z(ram_a_block_N_2299)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(109[49:72])
    defparam i1_4_lut_adj_579.init = 16'hffef;
    LUT4 i1_2_lut (.A(instr_active), .B(last_ram_a_sel), .Z(n28149)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(109[49:72])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 spi_clk_pos_I_0_256_3_lut_rep_830 (.A(spi_clk_pos), .B(spi_clk_neg), 
         .C(spi_clk_use_neg), .Z(spi_clk_pos_derived_59)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(287[26:69])
    defparam spi_clk_pos_I_0_256_3_lut_rep_830.init = 16'hcaca;
    LUT4 qspi_clk_I_0_1_lut_3_lut (.A(spi_clk_pos), .B(spi_clk_neg), .C(spi_clk_use_neg), 
         .Z(qspi_clk_N_56)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(287[26:69])
    defparam qspi_clk_I_0_1_lut_3_lut.init = 16'h3535;
    LUT4 fsm_state_2__bdd_4_lut_29315 (.A(fsm_state[2]), .B(fsm_state[0]), 
         .C(fsm_state[1]), .D(n32542), .Z(n27342)) /* synthesis lut_function=(A (B (D)+!B !(C))) */ ;
    defparam fsm_state_2__bdd_4_lut_29315.init = 16'h8a02;
    LUT4 i8976_1_lut (.A(\write_qspi_data_byte_idx_1__N_2021[0] ), .Z(n11684)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i8976_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_580 (.A(qspi_data_ready), .B(data_stall), .C(n32712), 
         .D(n32686), .Z(n11193)) /* synthesis lut_function=(A+!(B (C)+!B (C+(D)))) */ ;
    defparam i1_4_lut_adj_580.init = 16'haeaf;
    LUT4 i3179_4_lut (.A(n32681), .B(n32522), .C(n32755), .D(n32743), 
         .Z(n6220)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i3179_4_lut.init = 16'hac0c;
    LUT4 mux_95_i1_3_lut_4_lut_4_lut_4_lut (.A(fsm_state[0]), .B(n32753), 
         .C(is_writing), .D(\writing_N_164[3] ), .Z(n312[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(266[13:21])
    defparam mux_95_i1_3_lut_4_lut_4_lut_4_lut.init = 16'h7475;
    LUT4 i15226_4_lut (.A(nibbles_remaining[0]), .B(n1072), .C(n31866), 
         .D(n10820), .Z(n1064)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i15226_4_lut.init = 16'hcddd;
    FD1P3JX spi_ram_a_select_228 (.D(spi_ram_a_select_N_2309), .SP(clk_c_enable_543), 
            .PD(n32524), .CK(clk_c), .Q(qspi_ram_a_select)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_ram_a_select_228.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_581 (.A(fsm_state[0]), .B(stop_txn_reg), .C(fsm_state[1]), 
         .D(fsm_state[2]), .Z(n28319)) /* synthesis lut_function=(A (B)+!A (B+(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam i1_4_lut_adj_581.init = 16'hdccd;
    PFUMX mux_129_i1 (.BLUT(n181[0]), .ALUT(n381[0]), .C0(n32743), .Z(n396[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    FD1P3JX spi_ram_b_select_229 (.D(spi_ram_b_select_N_2313), .SP(clk_c_enable_543), 
            .PD(n32524), .CK(clk_c), .Q(qspi_ram_b_select)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_ram_b_select_229.GSR = "DISABLED";
    FD1P3JX spi_flash_select_227 (.D(\addr_in[24] ), .SP(clk_c_enable_543), 
            .PD(n32524), .CK(clk_c), .Q(\writing_N_164[3] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_flash_select_227.GSR = "DISABLED";
    PFUMX i15823 (.BLUT(n333[1]), .ALUT(n127[1]), .C0(n27343), .Z(n396[1]));
    PFUMX mux_687_i2 (.BLUT(n356[1]), .ALUT(n5181[0]), .C0(n17882), .Z(n1042));
    LUT4 mux_706_i3_4_lut (.A(n4330[2]), .B(\addr_in[24] ), .C(n1072), 
         .D(n26894), .Z(n11068)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam mux_706_i3_4_lut.init = 16'h353a;
    LUT4 fsm_state_2__bdd_4_lut_29782 (.A(fsm_state[2]), .B(fsm_state[0]), 
         .C(fsm_state[1]), .D(n32740), .Z(n32874)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+(C+(D))))) */ ;
    defparam fsm_state_2__bdd_4_lut_29782.init = 16'h0021;
    LUT4 i1_2_lut_4_lut_adj_582 (.A(spi_clk_pos), .B(n32777), .C(n17865), 
         .D(n32740), .Z(n26814)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[25:140])
    defparam i1_2_lut_4_lut_adj_582.init = 16'h00a3;
    LUT4 i28535_4_lut (.A(n32743), .B(stop_txn_now_N_2363), .C(n28259), 
         .D(n32755), .Z(n27903)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i28535_4_lut.init = 16'h0200;
    LUT4 i27968_3_lut_4_lut (.A(\instr_data[8] ), .B(n32713), .C(n32674), 
         .D(n29768), .Z(instr_data_15__N_1959[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam i27968_3_lut_4_lut.init = 16'h8f80;
    LUT4 i27974_3_lut_4_lut (.A(\instr_data[11] ), .B(n32713), .C(n32674), 
         .D(n29777), .Z(instr_data_15__N_1959[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam i27974_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_4_lut_adj_583 (.A(n10), .B(n19867), .C(is_writing), .D(data_stall), 
         .Z(data_ready_N_2338)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_583.init = 16'h0002;
    LUT4 i21_4_lut (.A(n32817), .B(\read_cycles_count[1] ), .C(n32743), 
         .D(n26814), .Z(n10)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A !(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(165[26] 212[20])
    defparam i21_4_lut.init = 16'ha303;
    LUT4 n9_bdd_4_lut_28720 (.A(n32709), .B(\qspi_data_in[0] ), .C(spi_in_buffer[0]), 
         .D(rst_reg_n), .Z(n31472)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam n9_bdd_4_lut_28720.init = 16'he4a0;
    PFUMX mux_113_i1 (.BLUT(n312[0]), .ALUT(n332), .C0(n30110), .Z(n356[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 addr_23__bdd_3_lut_29044 (.A(addr[23]), .B(n32059), .C(fsm_state[0]), 
         .Z(n32060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam addr_23__bdd_3_lut_29044.init = 16'hcaca;
    LUT4 addr_23__bdd_4_lut (.A(\instr_data[15] ), .B(fsm_state[2]), .C(is_writing), 
         .D(nibbles_remaining[0]), .Z(n32059)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B (C)+!B (C+(D)))) */ ;
    defparam addr_23__bdd_4_lut.init = 16'h8c8f;
    LUT4 n9_bdd_3_lut_29181_4_lut (.A(fsm_state[1]), .B(n32744), .C(spi_in_buffer[1]), 
         .D(qspi_data_out_3__N_5[1]), .Z(n31674)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[102:126])
    defparam n9_bdd_3_lut_29181_4_lut.init = 16'hf1e0;
    LUT4 i28480_2_lut_4_lut_4_lut (.A(n32744), .B(is_writing), .C(n32674), 
         .D(n32696), .Z(clk_c_enable_511)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (C (D))))) */ ;
    defparam i28480_2_lut_4_lut_4_lut.init = 16'h1ddd;
    LUT4 i14917_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n32820), .C(debug_stop_txn_N_2119), 
         .D(qspi_write_done), .Z(debug_stop_txn)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i14917_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 n18361_bdd_3_lut_28695_4_lut (.A(n32739), .B(n32740), .C(rst_reg_n), 
         .D(\qspi_data_in[0] ), .Z(n31474)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam n18361_bdd_3_lut_28695_4_lut.init = 16'h4000;
    LUT4 n18361_bdd_3_lut_28795_4_lut (.A(n32739), .B(n32740), .C(rst_reg_n), 
         .D(\qspi_data_in[2] ), .Z(n31645)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam n18361_bdd_3_lut_28795_4_lut.init = 16'h4000;
    LUT4 n18361_bdd_3_lut_28786_4_lut (.A(n32739), .B(n32740), .C(rst_reg_n), 
         .D(\qspi_data_in[3] ), .Z(n31638)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam n18361_bdd_3_lut_28786_4_lut.init = 16'h4000;
    L6MUX21 i28823 (.D0(n31678), .D1(n31675), .SD(n30226), .Z(data_out_7__N_2177[1]));
    PFUMX i28821 (.BLUT(n31677), .ALUT(n31676), .C0(n32674), .Z(n31678));
    LUT4 i1_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(\read_cycles_count[1] ), 
         .Z(n29577)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    PFUMX i28819 (.BLUT(n29755), .ALUT(n31674), .C0(n32830), .Z(n31675));
    LUT4 mux_113_i3_4_lut_then_4_lut (.A(n32740), .B(fsm_state[0]), .C(fsm_state[1]), 
         .D(fsm_state[2]), .Z(n32856)) /* synthesis lut_function=(A (B (C (D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_113_i3_4_lut_then_4_lut.init = 16'hd550;
    LUT4 i20_4_lut (.A(n32744), .B(n32674), .C(is_writing), .D(n6), 
         .Z(clk_c_enable_507)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;
    defparam i20_4_lut.init = 16'hf535;
    LUT4 i15466_3_lut_4_lut (.A(n32522), .B(n32755), .C(n17882), .D(n32857), 
         .Z(n1057)) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i15466_3_lut_4_lut.init = 16'hddd0;
    L6MUX21 i28798 (.D0(n31647), .D1(n31644), .SD(n30226), .Z(data_out_7__N_2177[2]));
    LUT4 i15700_3_lut_rep_659_4_lut_3_lut (.A(n32740), .B(n32743), .C(spi_clk_pos), 
         .Z(n32674)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(231[22] 237[16])
    defparam i15700_3_lut_rep_659_4_lut_3_lut.init = 16'h8c8c;
    PFUMX i28796 (.BLUT(n31646), .ALUT(n31645), .C0(n32674), .Z(n31647));
    PFUMX i28792 (.BLUT(n29761), .ALUT(n31643), .C0(n32830), .Z(n31644));
    L6MUX21 i28789 (.D0(n31640), .D1(n31637), .SD(n30226), .Z(data_out_7__N_2177[3]));
    PFUMX i28787 (.BLUT(n31639), .ALUT(n31638), .C0(n32674), .Z(n31640));
    PFUMX i28784 (.BLUT(n29764), .ALUT(n31636), .C0(n32830), .Z(n31637));
    LUT4 mux_113_i3_4_lut_else_4_lut (.A(n32740), .B(fsm_state[0]), .C(fsm_state[1]), 
         .D(fsm_state[2]), .Z(n32855)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_113_i3_4_lut_else_4_lut.init = 16'hd540;
    LUT4 i1_4_lut_4_lut_adj_584 (.A(n32740), .B(n32722), .C(n32536), .D(n29375), 
         .Z(n356[1])) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_4_lut_4_lut_adj_584.init = 16'h5450;
    LUT4 n5554_bdd_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n32775), .C(qspi_data_out_3__N_5[1]), 
         .D(n32740), .Z(n31676)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam n5554_bdd_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_adj_585 (.A(fsm_state[2]), .B(n32775), .C(is_writing), 
         .D(n32740), .Z(data_req_N_2318)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_3_lut_4_lut_adj_585.init = 16'h0020;
    LUT4 i15216_3_lut_4_lut (.A(fsm_state[2]), .B(n32775), .C(is_writing), 
         .D(data_req_N_2334), .Z(n17865)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i15216_3_lut_4_lut.init = 16'h00fd;
    LUT4 i825_2_lut_rep_681_3_lut_4_lut (.A(fsm_state[2]), .B(n32775), .C(spi_clk_pos), 
         .D(n32740), .Z(n32696)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A ((D)+!C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i825_2_lut_rep_681_3_lut_4_lut.init = 16'hdf0f;
    LUT4 i1_2_lut_3_lut_4_lut_adj_586 (.A(fsm_state[2]), .B(n32775), .C(spi_clk_pos), 
         .D(n32740), .Z(n6)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_3_lut_4_lut_adj_586.init = 16'h20f0;
    LUT4 i1_2_lut_rep_652_3_lut_4_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n32775), 
         .C(spi_clk_pos), .D(n32740), .Z(n32667)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_652_3_lut_4_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_adj_587 (.A(nibbles_remaining[0]), .B(n32778), .C(data_req_N_2334), 
         .D(n17882), .Z(n28111)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_3_lut_4_lut_adj_587.init = 16'h000e;
    LUT4 i1_3_lut_4_lut_adj_588 (.A(nibbles_remaining[0]), .B(n32778), .C(n27342), 
         .D(n32681), .Z(n1164)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_3_lut_4_lut_adj_588.init = 16'hefff;
    LUT4 i3440_2_lut_rep_698_3_lut_4_lut (.A(nibbles_remaining[0]), .B(n32778), 
         .C(n32775), .D(fsm_state[2]), .Z(n32713)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i3440_2_lut_rep_698_3_lut_4_lut.init = 16'h0e00;
    LUT4 i3181_3_lut_4_lut (.A(n32523), .B(ram_b_block_N_2303), .C(n32755), 
         .D(data_ready_N_2347), .Z(n6216)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i3181_3_lut_4_lut.init = 16'hf808;
    LUT4 i28374_3_lut_4_lut (.A(fsm_state[0]), .B(n32782), .C(n32789), 
         .D(n19867), .Z(n17882)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(169[58:88])
    defparam i28374_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_3_lut_4_lut_adj_589 (.A(n32523), .B(ram_b_block_N_2303), .C(n32755), 
         .D(n32524), .Z(clk_c_enable_438)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i1_3_lut_4_lut_adj_589.init = 16'hfff8;
    LUT4 i1_2_lut_rep_694_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(n32777), 
         .D(fsm_state[1]), .Z(n32709)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_694_4_lut.init = 16'hfff7;
    LUT4 i1_3_lut_adj_590 (.A(debug_stop_txn), .B(stop_txn_now_N_2363), 
         .C(stop_txn_reg), .Z(stop_txn_reg_N_2360)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut_adj_590.init = 16'h0202;
    LUT4 i28454_3_lut_4_lut (.A(n32778), .B(nibbles_remaining[0]), .C(n1072), 
         .D(n4330[1]), .Z(n18383)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam i28454_3_lut_4_lut.init = 16'h0d02;
    PFUMX i29305 (.BLUT(n32855), .ALUT(n32856), .C0(n32823), .Z(n32857));
    PFUMX i29326 (.BLUT(n32890), .ALUT(n32891), .C0(n5188[0]), .Z(n32892));
    PFUMX i29324 (.BLUT(n32887), .ALUT(n32888), .C0(n32740), .Z(n4330[1]));
    
endmodule
//
// Verilog Description of module tinyqv_cpu
//

module tinyqv_cpu (imm, clk_c, \instr[31] , \imm[13] , n32578, \imm[12] , 
            \imm[11] , \imm[10] , \imm[9] , \imm[8] , \imm[7] , \imm[6] , 
            \imm[5] , \imm[4] , \imm[3] , \imm[2] , \imm[1] , was_early_branch, 
            data_to_write, addr, rd, qv_data_read_n, n29738, \instr_data[3]_adj_13 , 
            \instr_addr_23__N_318[0] , n32656, n26116, debug_data_continue, 
            debug_instr_valid, n32851, n32835, n32723, \gpio_out_func_sel[5][2] , 
            \gpio_out_func_sel[7][2] , \instr_len[2] , \pc[2] , \pc[1] , 
            n2196, n32727, n2191, n32640, instr_data, n32548, n32734, 
            \qspi_data_buf[10] , \qspi_data_buf[14] , n32836, n27888, 
            \gpio_out_func_sel[5][4] , \gpio_out_func_sel[7][4] , n29831, 
            n32655, n34287, instr_fetch_running, n32544, n32537, instr_fetch_running_N_945, 
            n19867, \instr_write_offset[3] , qspi_data_byte_idx, qspi_data_ready, 
            n2150, n2130, n4251, n32685, n19, n32660, \qspi_data_buf[11] , 
            \qspi_data_buf[15] , \peri_data_out[11] , n4, \peri_data_out[10] , 
            n32642, \mem_data_from_read[20] , \mem_data_from_read[16] , 
            n32771, \peri_data_out[9] , rst_reg_n_adj_6, n31796, n31795, 
            n32520, n21414, n32654, \pc[7] , \pc[15] , n32842, \next_pc_for_core[6] , 
            \pc[3] , \pc[11] , n32251, n31706, clk_c_enable_285, n28957, 
            n34285, \pc[6] , \pc[14] , \pc[10] , n3, n3_adj_7, n32638, 
            n29707, qv_data_write_n, n32850, \addr[24] , \addr[23] , 
            \addr[22] , \addr[21] , \imm[21] , \imm[20] , \next_pc_for_core[9] , 
            \next_pc_for_core[13] , \addr[20] , \addr[19] , \addr[18] , 
            \addr[17] , \addr[16] , \pc[5] , \pc[13] , \addr[15] , 
            \pc[9] , \addr[14] , \addr[13] , \addr[12] , \addr[11] , 
            \addr[9] , \addr[8] , \addr[5] , \addr[4] , \addr[1] , 
            \next_pc_for_core[4] , n12, data_ready_r_N_2823, data_ready_r, 
            n32801, n29059, n32598, data_txn_len, n32714, n32689, 
            n32531, rst_reg_n, n32706, n15569, n2211, n17165, VCC_net, 
            n32694, n7, n8854, \next_pc_for_core[10] , \next_pc_for_core[14] , 
            debug_stop_txn_N_2142, \instr_data[0][0] , \instr_data[1][7] , 
            \instr_data[1][0] , \instr_data[2][7] , data_stall, n32542, 
            \next_pc_for_core[8] , \next_pc_for_core[12] , n32787, n32740, 
            data_req_N_2334, n332, instr_active, n11193, clk_c_enable_91, 
            \mem_data_from_read[19] , \mem_data_from_read[23] , n32788, 
            n1, n175, \read_cycles_count[1] , n32789, data_ready_N_2347, 
            \instr_data[2][0] , \instr_data[3][7] , n32545, n32552, 
            n8109, n32695, n32728, n32712, n32745, \next_pc_for_core[3] , 
            \next_pc_for_core[5] , \next_pc_for_core[7] , \next_pc_for_core[11] , 
            \pc[21] , \pc[17] , \next_pc_for_core[20] , \next_pc_for_core[16] , 
            \pc[23] , \pc[19] , \pc[22] , \pc[18] , \pc[20] , \pc[16] , 
            \next_pc_for_core[15] , \next_pc_for_core[21] , \next_pc_for_core[17] , 
            \imm[23] , \imm[22] , \imm[19] , \imm[18] , \next_pc_for_core[22] , 
            \next_pc_for_core[18] , \next_pc_for_core[19] , n28077, \next_pc_for_core[23] , 
            n32819, n32720, n29357, \uo_out_from_user_peri[1][6] , \data_from_user_peri_1__31__N_2455[2] , 
            \uo_out_from_user_peri[1][2] , \uo_out_from_user_peri[1][5] , 
            n29491, \data_from_read[2] , \early_branch_addr[7] , \early_branch_addr[3] , 
            \early_branch_addr[6] , \early_branch_addr[2] , \early_branch_addr[4] , 
            n32822, \early_branch_addr[8] , \early_branch_addr[5] , \early_branch_addr[9] , 
            \early_branch_addr[10] , \early_branch_addr[11] , \early_branch_addr[12] , 
            \early_branch_addr[13] , \early_branch_addr[14] , \early_branch_addr[15] , 
            \early_branch_addr[17] , \early_branch_addr[18] , \early_branch_addr[19] , 
            \early_branch_addr[20] , \early_branch_addr[21] , \early_branch_addr[22] , 
            \early_branch_addr[23] , \early_branch_addr[16] , n16811, 
            n2594, n31883, \pc_23__N_911[13] , \pc[12] , n26838, n10944, 
            n32725, n32761, n32729, \cycle[0] , debug_data_ready, 
            \pc[8] , n27178, n32766, \pc[4] , n32711, n32737, \data_from_peri_31__N_2415[0] , 
            fsm_state, n32778, n31866, n32693, clk_c_enable_50, n32818, 
            clk_c_enable_154, clk_c_enable_283, clk_c_enable_354, \gpio_out_func_sel[0][2] , 
            \gpio_out_func_sel[1][2] , \gpio_out_func_sel[2][2] , \gpio_out_func_sel[3][2] , 
            n32756, n5169, n29618, start_instr, n32825, n29127, 
            n18458, \gpio_out_func_sel[4][2] , \gpio_out_func_sel[6][2] , 
            n8, \uart_rx_buf_data[4] , \baud_divider[4] , instr_fetch_stopped, 
            n16, n32826, \instr_data_7__N_1969[3] , \instr_data_7__N_1969[1] , 
            gpio_out_sel, n14, n14_adj_8, n29293, instr_complete_N_1647, 
            \data_from_read[6] , n32672, n46, \connect_peripheral[1] , 
            \connect_peripheral[0] , \qspi_data_buf[9] , \qspi_data_buf[13] , 
            \instr_addr[2] , n32568, n29741, n29, \uart_rx_buf_data[7] , 
            \baud_divider[7] , n2, n32614, \next_fsm_state_3__N_3046[3] , 
            \ui_in_sync[5] , \ui_in_sync[6] , n32072, n29549, \ui_in_sync[7] , 
            \data_from_user_peri_1__31__N_2455[7] , \uart_rx_buf_data[6] , 
            n26856, \baud_divider[6] , \uart_rx_buf_data[5] , \baud_divider[5] , 
            \mem_data_from_read[4] , \data_from_read[4] , \mem_data_from_read[8] , 
            \data_from_read[8] , \mem_data_from_read[12] , \data_from_read[12] , 
            \mem_data_from_read[1] , \data_from_read[1] , \data_from_user_peri_1__31__N_2455[0] , 
            \uo_out_from_user_peri[1][0] , \mem_data_from_read[5] , \data_from_read[5] , 
            data_out_hold, \mem_data_from_read[3] , \data_from_read[3] , 
            \mem_data_from_read[7] , \data_from_read[7] , \uart_rx_buf_data[3] , 
            \baud_divider[3] , n2_adj_9, \mem_data_from_read[0] , \data_from_read[0] , 
            n32759, \mem_data_from_read[18] , \mem_data_from_read[22] , 
            \mem_data_from_read[26] , \mem_data_from_read[30] , \mem_data_from_read[24] , 
            \mem_data_from_read[28] , \uart_rx_buf_data[2] , \baud_divider[2] , 
            \mem_data_from_read[27] , \mem_data_from_read[31] , \mem_data_from_read[25] , 
            \mem_data_from_read[29] , n10737, n32650, \instr[16] , n32615, 
            n32610, clk_c_enable_342, \ui_in_sync[1] , \ui_in_sync[0] , 
            debug_rd, n29866, n17920, n28687, accum, d_3__N_1868, 
            fsm_state_adj_14, n32791, n32763, n32730, n32834, n32710, 
            n31351, n1152, \mem_data_from_read[17] , \mem_data_from_read[21] , 
            \mul_out[3] , \mul_out[2] , \mul_out[1] , \csr_read_3__N_1447[2] , 
            \next_accum[5] , GND_net, \next_accum[16] , \next_accum[17] , 
            \next_accum[18] , \next_accum[19] , \next_accum[6] , \next_accum[7] , 
            \next_accum[8] , \next_accum[9] , \next_accum[10] , \next_accum[11] , 
            \next_accum[12] , \next_accum[13] , \next_accum[14] , \next_accum[15] , 
            \next_accum[4] , \return_addr[16] ) /* synthesis syn_module_defined=1 */ ;
    output [31:0]imm;
    input clk_c;
    output \instr[31] ;
    output \imm[13] ;
    input n32578;
    output \imm[12] ;
    output \imm[11] ;
    output \imm[10] ;
    output \imm[9] ;
    output \imm[8] ;
    output \imm[7] ;
    output \imm[6] ;
    output \imm[5] ;
    output \imm[4] ;
    output \imm[3] ;
    output \imm[2] ;
    output \imm[1] ;
    output was_early_branch;
    output [31:0]data_to_write;
    output [27:0]addr;
    output [3:0]rd;
    output [1:0]qv_data_read_n;
    input n29738;
    output [15:0]\instr_data[3]_adj_13 ;
    output \instr_addr_23__N_318[0] ;
    output n32656;
    output n26116;
    output debug_data_continue;
    output debug_instr_valid;
    output n32851;
    output n32835;
    output n32723;
    input \gpio_out_func_sel[5][2] ;
    input \gpio_out_func_sel[7][2] ;
    output \instr_len[2] ;
    output \pc[2] ;
    output \pc[1] ;
    output n2196;
    output n32727;
    output n2191;
    output n32640;
    input [15:0]instr_data;
    output n32548;
    output n32734;
    input \qspi_data_buf[10] ;
    input \qspi_data_buf[14] ;
    input n32836;
    output n27888;
    input \gpio_out_func_sel[5][4] ;
    input \gpio_out_func_sel[7][4] ;
    output n29831;
    output n32655;
    input n34287;
    output instr_fetch_running;
    output n32544;
    output n32537;
    input instr_fetch_running_N_945;
    output n19867;
    output \instr_write_offset[3] ;
    input [1:0]qspi_data_byte_idx;
    input qspi_data_ready;
    input n2150;
    input n2130;
    output n4251;
    output n32685;
    output n19;
    output n32660;
    input \qspi_data_buf[11] ;
    input \qspi_data_buf[15] ;
    input \peri_data_out[11] ;
    output n4;
    input \peri_data_out[10] ;
    output n32642;
    input \mem_data_from_read[20] ;
    input \mem_data_from_read[16] ;
    output n32771;
    input \peri_data_out[9] ;
    input rst_reg_n_adj_6;
    input n31796;
    input n31795;
    output n32520;
    output n21414;
    input n32654;
    output \pc[7] ;
    output \pc[15] ;
    output n32842;
    input \next_pc_for_core[6] ;
    output \pc[3] ;
    output \pc[11] ;
    input n32251;
    input n31706;
    output clk_c_enable_285;
    output n28957;
    output n34285;
    output \pc[6] ;
    output \pc[14] ;
    output \pc[10] ;
    output n3;
    output n3_adj_7;
    input n32638;
    input n29707;
    output [1:0]qv_data_write_n;
    output n32850;
    output \addr[24] ;
    output \addr[23] ;
    output \addr[22] ;
    output \addr[21] ;
    output \imm[21] ;
    output \imm[20] ;
    input \next_pc_for_core[9] ;
    input \next_pc_for_core[13] ;
    output \addr[20] ;
    output \addr[19] ;
    output \addr[18] ;
    output \addr[17] ;
    output \addr[16] ;
    output \pc[5] ;
    output \pc[13] ;
    output \addr[15] ;
    output \pc[9] ;
    output \addr[14] ;
    output \addr[13] ;
    output \addr[12] ;
    output \addr[11] ;
    output \addr[9] ;
    output \addr[8] ;
    output \addr[5] ;
    output \addr[4] ;
    output \addr[1] ;
    input \next_pc_for_core[4] ;
    input n12;
    output data_ready_r_N_2823;
    input data_ready_r;
    output n32801;
    output n29059;
    input n32598;
    input [1:0]data_txn_len;
    output n32714;
    input n32689;
    output n32531;
    input rst_reg_n;
    output n32706;
    output n15569;
    output n2211;
    input n17165;
    input VCC_net;
    output n32694;
    output n7;
    input n8854;
    input \next_pc_for_core[10] ;
    input \next_pc_for_core[14] ;
    output debug_stop_txn_N_2142;
    output \instr_data[0][0] ;
    output \instr_data[1][7] ;
    output \instr_data[1][0] ;
    output \instr_data[2][7] ;
    input data_stall;
    output n32542;
    input \next_pc_for_core[8] ;
    input \next_pc_for_core[12] ;
    output n32787;
    input n32740;
    input data_req_N_2334;
    output n332;
    input instr_active;
    input n11193;
    output clk_c_enable_91;
    input \mem_data_from_read[19] ;
    input \mem_data_from_read[23] ;
    output n32788;
    input n1;
    output n175;
    input \read_cycles_count[1] ;
    output n32789;
    output data_ready_N_2347;
    output \instr_data[2][0] ;
    output \instr_data[3][7] ;
    output n32545;
    output n32552;
    output n8109;
    output n32695;
    output n32728;
    output n32712;
    output n32745;
    input \next_pc_for_core[3] ;
    input \next_pc_for_core[5] ;
    input \next_pc_for_core[7] ;
    input \next_pc_for_core[11] ;
    output \pc[21] ;
    output \pc[17] ;
    input \next_pc_for_core[20] ;
    input \next_pc_for_core[16] ;
    output \pc[23] ;
    output \pc[19] ;
    output \pc[22] ;
    output \pc[18] ;
    output \pc[20] ;
    output \pc[16] ;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[21] ;
    input \next_pc_for_core[17] ;
    output \imm[23] ;
    output \imm[22] ;
    output \imm[19] ;
    output \imm[18] ;
    input \next_pc_for_core[22] ;
    input \next_pc_for_core[18] ;
    input \next_pc_for_core[19] ;
    output n28077;
    input \next_pc_for_core[23] ;
    output n32819;
    output n32720;
    output n29357;
    input \uo_out_from_user_peri[1][6] ;
    input \data_from_user_peri_1__31__N_2455[2] ;
    input \uo_out_from_user_peri[1][2] ;
    input \uo_out_from_user_peri[1][5] ;
    output n29491;
    input \data_from_read[2] ;
    input \early_branch_addr[7] ;
    input \early_branch_addr[3] ;
    input \early_branch_addr[6] ;
    input \early_branch_addr[2] ;
    input \early_branch_addr[4] ;
    input n32822;
    input \early_branch_addr[8] ;
    input \early_branch_addr[5] ;
    input \early_branch_addr[9] ;
    input \early_branch_addr[10] ;
    input \early_branch_addr[11] ;
    input \early_branch_addr[12] ;
    input \early_branch_addr[13] ;
    input \early_branch_addr[14] ;
    input \early_branch_addr[15] ;
    input \early_branch_addr[17] ;
    input \early_branch_addr[18] ;
    input \early_branch_addr[19] ;
    input \early_branch_addr[20] ;
    input \early_branch_addr[21] ;
    input \early_branch_addr[22] ;
    input \early_branch_addr[23] ;
    input \early_branch_addr[16] ;
    output n16811;
    input n2594;
    output n31883;
    input \pc_23__N_911[13] ;
    output \pc[12] ;
    output n26838;
    input n10944;
    output n32725;
    output n32761;
    output n32729;
    output \cycle[0] ;
    input debug_data_ready;
    output \pc[8] ;
    output n27178;
    output n32766;
    output \pc[4] ;
    output n32711;
    output n32737;
    output \data_from_peri_31__N_2415[0] ;
    input [2:0]fsm_state;
    input n32778;
    output n31866;
    output n32693;
    output clk_c_enable_50;
    input n32818;
    output clk_c_enable_154;
    output clk_c_enable_283;
    output clk_c_enable_354;
    input \gpio_out_func_sel[0][2] ;
    input \gpio_out_func_sel[1][2] ;
    input \gpio_out_func_sel[2][2] ;
    input \gpio_out_func_sel[3][2] ;
    input n32756;
    output n5169;
    input n29618;
    output start_instr;
    input n32825;
    input n29127;
    output n18458;
    input \gpio_out_func_sel[4][2] ;
    input \gpio_out_func_sel[6][2] ;
    output n8;
    input \uart_rx_buf_data[4] ;
    input \baud_divider[4] ;
    input instr_fetch_stopped;
    input n16;
    input n32826;
    output \instr_data_7__N_1969[3] ;
    output \instr_data_7__N_1969[1] ;
    input [7:6]gpio_out_sel;
    output n14;
    output n14_adj_8;
    output n29293;
    output instr_complete_N_1647;
    input \data_from_read[6] ;
    output n32672;
    output n46;
    output \connect_peripheral[1] ;
    output \connect_peripheral[0] ;
    input \qspi_data_buf[9] ;
    input \qspi_data_buf[13] ;
    output \instr_addr[2] ;
    input n32568;
    output n29741;
    input n29;
    input \uart_rx_buf_data[7] ;
    input \baud_divider[7] ;
    output n2;
    input n32614;
    input \next_fsm_state_3__N_3046[3] ;
    input \ui_in_sync[5] ;
    input \ui_in_sync[6] ;
    input n32072;
    output n29549;
    input \ui_in_sync[7] ;
    output \data_from_user_peri_1__31__N_2455[7] ;
    input \uart_rx_buf_data[6] ;
    input n26856;
    input \baud_divider[6] ;
    input \uart_rx_buf_data[5] ;
    input \baud_divider[5] ;
    input \mem_data_from_read[4] ;
    input \data_from_read[4] ;
    input \mem_data_from_read[8] ;
    input \data_from_read[8] ;
    input \mem_data_from_read[12] ;
    input \data_from_read[12] ;
    input \mem_data_from_read[1] ;
    input \data_from_read[1] ;
    input \data_from_user_peri_1__31__N_2455[0] ;
    input \uo_out_from_user_peri[1][0] ;
    input \mem_data_from_read[5] ;
    input \data_from_read[5] ;
    input data_out_hold;
    input \mem_data_from_read[3] ;
    input \data_from_read[3] ;
    input \mem_data_from_read[7] ;
    input \data_from_read[7] ;
    input \uart_rx_buf_data[3] ;
    input \baud_divider[3] ;
    output n2_adj_9;
    input \mem_data_from_read[0] ;
    input \data_from_read[0] ;
    output n32759;
    input \mem_data_from_read[18] ;
    input \mem_data_from_read[22] ;
    input \mem_data_from_read[26] ;
    input \mem_data_from_read[30] ;
    input \mem_data_from_read[24] ;
    input \mem_data_from_read[28] ;
    input \uart_rx_buf_data[2] ;
    input \baud_divider[2] ;
    input \mem_data_from_read[27] ;
    input \mem_data_from_read[31] ;
    input \mem_data_from_read[25] ;
    input \mem_data_from_read[29] ;
    input n10737;
    output n32650;
    input \instr[16] ;
    input n32615;
    input n32610;
    input clk_c_enable_342;
    input \ui_in_sync[1] ;
    input \ui_in_sync[0] ;
    output [3:0]debug_rd;
    input n29866;
    output n17920;
    output n28687;
    output [15:0]accum;
    output [19:0]d_3__N_1868;
    input [3:0]fsm_state_adj_14;
    output n32791;
    output n32763;
    output n32730;
    output n32834;
    output n32710;
    input n31351;
    output n1152;
    input \mem_data_from_read[17] ;
    input \mem_data_from_read[21] ;
    input \mul_out[3] ;
    input \mul_out[2] ;
    input \mul_out[1] ;
    output \csr_read_3__N_1447[2] ;
    input \next_accum[5] ;
    input GND_net;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[4] ;
    output \return_addr[16] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire clk_c_enable_383, n32022, n32630, n32563, n32540;
    wire [12:0]n4969;
    wire [31:0]n3534;
    wire [31:0]imm_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(100[16:19])
    
    wire n32383, n32382, n32384, clk_c_enable_15;
    wire [3:0]alu_op;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    
    wire clk_c_enable_338, n32840;
    wire [3:0]alu_op_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(64[16:25])
    
    wire clk_c_enable_28, debug_early_branch, clk_c_enable_207;
    wire [3:0]data_out_slice;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(230[16:30])
    wire [2:0]additional_mem_ops;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(120[15:33])
    wire [2:0]additional_mem_ops_2__N_749;
    
    wire clk_c_enable_174;
    wire [27:0]addr_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(131[17:25])
    
    wire clk_c_enable_524, n33740;
    wire [2:1]instr_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(113[15:24])
    
    wire clk_c_enable_41, n32594;
    wire [2:0]mem_op;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(115[15:21])
    
    wire clk_c_enable_365;
    wire [2:0]mem_op_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(65[16:25])
    wire [3:0]rs1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(117[15:18])
    wire [3:0]n2632;
    
    wire clk_c_enable_122, n27629, n32539, clk_c_enable_309;
    wire [63:0]instr_data_0__15__N_638;
    
    wire data_ready_sync, data_ready_core;
    wire [2:0]instr_write_offset_3__N_934;
    
    wire n11, n13, n16_c, n26859, n5, clk_c_enable_52, data_continue_N_963, 
        is_load, clk_c_enable_364, is_load_de, n9, n12_c, n16_adj_3168, 
        n32316, n32314;
    wire [4:2]counter_hi;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(139[15:25])
    
    wire n32317, n32543, n10024, n12_adj_3169, n28527, n28533, n29834, 
        n4271;
    wire [31:0]n3369;
    wire [15:0]n5138;
    wire [31:0]n3410;
    
    wire n31590, n35, n10772, n22, n4_c, n27524, n32393, n32227, 
        n13456, n13_adj_3170, n27364, n13151, n29714, n29702, n32049, 
        n32394, n32541, n32191;
    wire [31:0]n3259;
    wire [31:0]n3292;
    
    wire n32659, n28547, n32252, n32253, n19_c, n32527, n30197, 
        n32551, n29732;
    wire [30:0]n5205;
    
    wire n32550, n28219, n2_c, n27851;
    wire [3:1]next_instr_write_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[16:39])
    
    wire n1_c, n68, n26962;
    wire [15:0]n33;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]n31;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire n32885;
    wire [15:0]n34;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]n36;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire n32884;
    wire [22:0]instr_addr_23__N_318;
    
    wire n32639, n32406;
    wire [3:0]n5658;
    wire [59:0]debug_rd_3__N_405;
    
    wire n32785, n9058;
    wire [59:0]debug_branch_N_446;
    
    wire n32897, n32407, n32896, n32900, n32899, n32268, n32267, 
        n32269, no_write_in_progress, clk_c_enable_99, no_write_in_progress_N_471, 
        n33055, n13_adj_3173, n33056, n30322, n33057, n32641, n28641, 
        n32859, n32651, n32637, n28605, n29700, n29712;
    wire [31:0]instr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(47[17:22])
    
    wire n32858, interrupt_core, clk_c_enable_545, n32546, n4267, 
        n4259;
    wire [31:0]n2970;
    
    wire n29723, debug_instr_valid_N_436, n32716, n32254, n32255, 
        n32525, n30024, n32595, n32488, n31620, n29727;
    wire [15:0]n2151;
    
    wire n32841, n29842, n26, n28669, n28635, n31621, n32533, 
        n29716, n29706, n32180, n33404, n28593, n32643, n28617;
    wire [23:1]return_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(135[17:28])
    wire [1:0]n1768;
    
    wire n31622, n31619, n34281;
    wire [59:0]debug_branch_N_442;
    
    wire stall_core, is_store, n31625, n32769, n8330, n30;
    wire [3:0]alu_op_3__N_1170;
    
    wire n9048, n32768, n32849, n32678, n32226, n32225, n31626, 
        n30920, n32494, n33403, n31627, n31624, n32493, n26857, 
        n21, n29718, n29704, n13140, n4265, n27489, n32222, n32221, 
        n32223, n26858, n20, n28653, n27480;
    wire [31:0]n3183;
    
    wire n30464, n28791, n32566, n32573, n28797, is_system, is_system_de, 
        n32661, n24898, clk_c_enable_513;
    wire [1:0]data_write_n_1__N_369;
    
    wire n27630, n32588;
    wire [3:0]rd_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(119[15:17])
    wire [3:0]n6;
    
    wire n32601, n32877, n28343, n32657, n32177, n32308, n32309;
    wire [27:0]addr_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    
    wire n26863, n25, n30463, n30462, n28763, n28769, n30461, 
        n17747, n37, n30457, n30456, n29710, n32901, n32395, n30365, 
        n32898, n32408, n32409, n28805, n28811, n30455, n28539, 
        n2792, n30454, n29837, n32599, n28777, n28783, n31650, 
        debug_rd_3__N_413, n32653, n28, n30160, n31651, n32812, 
        n27823;
    wire [1:0]n699;
    
    wire clk_c_enable_178, n32644;
    wire [3:2]addr_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(121[15:26])
    wire [1:0]n38;
    
    wire n32668, clk_c_enable_182, n149, clk_c_enable_187, clk_c_enable_191, 
        n32190, n32189, n32990, n29681, n32569, n31652, n31649, 
        n17, n32860, n32385, n32313, n32362, clk_c_enable_195, n32854, 
        n27294, n28851, clk_c_enable_200, n32176, n32178, n32993, 
        n32991, n32994, clk_c_enable_204, n32776, n32783, n28909, 
        n32658, n29661, n29031, n32538, n33737, n4_adj_3177, n28453, 
        n33738, n33735, is_branch, is_branch_de, load_started, address_ready, 
        n829, n26988, n29843, n30423, n30425, n28505, n30327, 
        n30329, n27653, n28889, n209, n32351, n32741, clk_c_enable_232, 
        is_lui, clk_c_enable_234, clk_c_enable_248, clk_c_enable_250, 
        clk_c_enable_292, n30179, n32784, n30172, n157, n32808, 
        n30070, is_jalr, is_jal, n30175;
    wire [3:0]n234;
    
    wire n32742, n28511;
    wire [15:0]n2202;
    
    wire n32585;
    wire [15:0]n2222;
    
    wire n30919, n29758;
    wire [1:0]txn_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(56[16:23])
    
    wire is_jalr_de;
    wire [15:0]n2131;
    
    wire n29840, load_top_bit, data_out_3__N_1385;
    wire [3:0]debug_branch_N_450;
    
    wire n29858, n29917, n29960, n32052, n32053, clk_c_enable_294, 
        clk_c_enable_308, n32796, n32051, n32050, n32797, n32798, 
        is_auipc, is_auipc_de;
    wire [31:0]n3493;
    wire [31:0]n3446;
    
    wire n32032, n32030, n32033, data_ready_latch, clk_c_enable_325, 
        n27854, n9620;
    wire [3:0]n5605;
    wire [3:0]n5640;
    
    wire n27, n29025, n32582, is_timer_addr, timer_data_3__N_631, 
        n29173, n32612, n32633, n32576, is_lui_N_1365;
    wire [3:0]alu_op_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[16:25])
    
    wire n22_adj_3179, n32027, n32024, n32028, n9_adj_3180, n28501, 
        n32664, is_jal_de, is_alu_imm;
    wire [3:0]data_rs2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(84[16:24])
    wire [3:0]n92;
    
    wire n29733, n24, n32611, n32340;
    wire [3:0]rs2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(118[15:18])
    wire [3:0]n2302;
    
    wire n20_adj_3181, n41, n27896, is_jal_N_1374;
    wire [20:0]n1742_adj_3219;
    
    wire n28249;
    wire [3:0]n328;
    
    wire n32581, n27788, n28269, mem_op_increment_reg;
    wire [3:0]n2281;
    
    wire n27430, n28715, is_lui_de, is_alu_reg, is_alu_reg_de, is_store_de, 
        is_alu_imm_de, mem_op_increment_reg_de, n32617, n32570, n28585, 
        n32020, n32017, n32021, clk_c_enable_367, n6396, n32704;
    wire [3:0]data_rs1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(83[16:24])
    
    wire n32702;
    wire [17:16]mip_reg;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(321[17:24])
    
    wire n21667, n34283, n28391, n225, n225_adj_3185, n226, n32034, 
        n32029, n227, n209_adj_3186, n157_adj_3187, n29689, n15_adj_3188, 
        n32754, n28575, n32853, clk_c_enable_538, n32677, n32760, 
        clk_c_enable_321, n32773, n17665, n6634, n32605, n32597, 
        n32629, n32628, n12_adj_3192, n30255, n30256, n30262, n30263, 
        n13156, n32613, n27428, n28407, n29211;
    wire [31:0]n3328;
    
    wire n32627, n32619, n32616, n19_adj_3193, n30132, n28731;
    wire [31:0]data_from_user_peri_1__31__N_2455;
    
    wire n29485;
    wire [3:0]n1708;
    
    wire n4243, n29594;
    wire [3:0]n2590;
    wire [3:0]n1713;
    
    wire n32992, n31589, n29163, n29165, n29161, n29155, n29145, 
        n32821;
    wire [20:0]n1203;
    
    wire n29159, n29141, n29039, n3_adj_3194, n32690;
    wire [1:0]n5017;
    
    wire n30261;
    wire [3:0]n2585;
    
    wire n30260, n32575, n32564, n32829, n8228, n32565, n2557, 
        n27516;
    wire [3:0]n2291;
    
    wire n27523;
    wire [2:0]n39;
    
    wire n30259, n32824, n27502, n28821, n27509, n9394, n32604, 
        n32609, n30258, n32828, load_done, instr_complete_N_1651, 
        n7_adj_3196, n30254, n32589, n32608, n30458, n30459, n30465, 
        n30466, n17_adj_3197, n32623, n31882, n31879, n30253;
    wire [2:0]additional_mem_ops_2__N_1132;
    
    wire n32560, n30252, n31878, n32632, n32602, n30251, clk_c_enable_533;
    wire [20:0]pc_23__N_911;
    
    wire n31588;
    wire [1:0]pc_2__N_932;
    
    wire n32427, n31881, n31880, n32634, n30014, n29696, n32561, 
        n32762, n31698, n8_c, n32875, n32721, n32583, n28435, 
        n32618, n149_adj_3198, n28447, n30007, n32603, n26879, n30037, 
        n32838, n32607;
    wire [1:0]cycle;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(58[15:20])
    
    wire n32767, n32848, n131, instr_complete_N_1652, n28561, n29600, 
        n2798;
    wire [3:0]n2618;
    
    wire n2796;
    wire [3:0]n2609;
    
    wire n28523, n2126, n24_adj_3199, n29605;
    wire [16:0]mie;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(323[16:19])
    
    wire n21665, n8_adj_3200, n793;
    wire [3:1]next_pc_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[16:30])
    
    wire n13152, n29695, n32682;
    wire [2:0]n1764;
    
    wire n29697, n824, n29705, n32549, n29703, n29726, n30084, 
        n29105, n29107, n29097, n29093;
    wire [3:0]n1734;
    wire [3:0]n1742;
    
    wire n29103, n29085, n27567, n2800, n13458, n32026, n30032, 
        n29_c, n28971, n32843, n29836, n10253, n32751, n32846, 
        n43, n2122, n28475, n32847, n24384, n27546, n19_adj_3201, 
        n672, n28733, n27541, n27545, n32547, n30929, n30930, 
        n32735, n24900, n27657, n2124, n27655, n27656, n13165, 
        n2_adj_3202, n4_adj_3203, n27804, n17949, n11066;
    wire [3:0]n2595;
    
    wire n13155, n2559, n28873, n27003, n27585, is_ret_de, n28685, 
        n27483, n27356, n27731, n28827, n32692, n13154;
    wire [31:0]n3222;
    
    wire n32530, n27492, n27427, n32707, n6920, n29725, n30041, 
        n27486, n27495, n58, n28963, n23;
    wire [3:0]n2577;
    
    wire n32806;
    wire [3:0]n155;
    
    wire n29119, n9052, n32487, n1_adj_3208, n32016, n32019, n32179, 
        n32671, n30928, n29745, n30927, n29743, n32025, n32774, 
        n30926, debug_early_branch_N_955, n30925, n28937, n28925, 
        n28919, n30924, n29747, n28647, n32031, n32732, n32733, 
        n32647, n4257, n32765, n28699, n28413, n29685, n28705, 
        n28719, n28553, n28611, n28567, n28599, n32489, n28755, 
        n28577, n29759, n11061;
    wire [59:0]debug_branch_N_840;
    
    wire n28747, n28837, n28429, n28441, n29760, n28739;
    wire [3:0]timer_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(143[16:26])
    
    wire n28673, n29844, n28417, n30320, n30321, n32571, n30_adj_3211, 
        n76, n28659, n33739, n33736, n28285, n30316, n30317, n30318, 
        n30319, n30323, n30324, n7_adj_3212, n29614, n30419, n30420, 
        n22_adj_3213, n32584, n32577, n29838, n32224, n32876, n29748, 
        n926, n28237, n28465, n32360, n32361, n28275, n28483, 
        debug_rd_3__N_1575, n19_adj_3214, n28623, n32, n32580, n27959, 
        n26937;
    wire [3:0]alu_op_3__N_1337;
    
    wire n893, n10, n18098, n28489, n28495, n32596, n29864, n860, 
        time_pulse_r, clk_c_enable_363, n32717;
    wire [31:0]mtimecmp;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(30[16:24])
    
    wire mtimecmp_1__N_1941;
    wire [3:0]mtime_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(29[16:25])
    
    wire timer_interrupt, mtimecmp_3__N_1935, cy, n32663, n32680, 
        mstatus_mie_N_1709, n32670, n32675, mstatus_mie_N_1707, n32758, 
        n32746, clk_c_enable_433, n32691, n29317;
    wire [3:0]\reg_access[4] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(30[16:26])
    wire [3:0]\reg_access[3] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(30[16:26])
    wire [6:0]cycle_count_wide;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(279[16:32])
    
    wire n32652, clk_c_enable_276, n32697, is_double_fault_r, mstatus_mte, 
        n32559, n28363;
    
    FD1P3AX imm_i0_i17 (.D(n32022), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm[17])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i17.GSR = "DISABLED";
    LUT4 mux_3051_i5_4_lut_4_lut (.A(\instr[31] ), .B(n32630), .C(n32563), 
         .D(n32540), .Z(n4969[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3051_i5_4_lut_4_lut.init = 16'ha088;
    FD1P3AX imm_i0_i16 (.D(n3534[16]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm[16])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i16.GSR = "DISABLED";
    FD1P3AX imm_i0_i15 (.D(n3534[15]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i15.GSR = "DISABLED";
    FD1P3AX imm_i0_i14 (.D(n3534[14]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i14.GSR = "DISABLED";
    FD1P3AX imm_i0_i0 (.D(n3534[0]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm_c[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i0.GSR = "DISABLED";
    FD1P3AX imm_i0_i13 (.D(n3534[13]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[13] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i13.GSR = "DISABLED";
    PFUMX i29218 (.BLUT(n32383), .ALUT(n32382), .C0(n32578), .Z(n32384));
    FD1P3AX imm_i0_i12 (.D(n3534[12]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[12] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i12.GSR = "DISABLED";
    FD1P3AX imm_i0_i11 (.D(n3534[11]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[11] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i11.GSR = "DISABLED";
    FD1P3AX imm_i0_i10 (.D(n3534[10]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[10] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i10.GSR = "DISABLED";
    FD1P3AX imm_i0_i9 (.D(n3534[9]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(\imm[9] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i9.GSR = "DISABLED";
    FD1P3AX imm_i0_i8 (.D(n3534[8]), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(\imm[8] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i8.GSR = "DISABLED";
    FD1P3AX imm_i0_i7 (.D(n3534[7]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i7.GSR = "DISABLED";
    FD1P3AX imm_i0_i6 (.D(n3534[6]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[6] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i6.GSR = "DISABLED";
    FD1P3AX imm_i0_i5 (.D(n3534[5]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[5] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i5.GSR = "DISABLED";
    FD1P3AX imm_i0_i4 (.D(n3534[4]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[4] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i4.GSR = "DISABLED";
    FD1P3IX alu_op__i0 (.D(alu_op_de[0]), .SP(clk_c_enable_338), .CD(n32840), 
            .CK(clk_c), .Q(alu_op[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i0.GSR = "DISABLED";
    FD1P3AX imm_i0_i3 (.D(n3534[3]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[3] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i3.GSR = "DISABLED";
    FD1P3AX imm_i0_i2 (.D(n3534[2]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[2] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i2.GSR = "DISABLED";
    FD1P3AX imm_i0_i1 (.D(n3534[1]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[1] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i1.GSR = "DISABLED";
    FD1P3IX was_early_branch_424 (.D(debug_early_branch), .SP(clk_c_enable_28), 
            .CD(n32840), .CK(clk_c), .Q(was_early_branch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(315[12] 320[8])
    defparam was_early_branch_424.GSR = "DISABLED";
    FD1P3IX data_out__i0 (.D(data_out_slice[0]), .SP(clk_c_enable_207), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i0.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i0 (.D(additional_mem_ops_2__N_749[0]), .CK(clk_c), 
            .CD(n32840), .Q(additional_mem_ops[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i0.GSR = "DISABLED";
    FD1P3IX data_addr__i0 (.D(addr_out[0]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(addr[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i0.GSR = "DISABLED";
    FD1P3AX rd_i0_i0 (.D(n33740), .SP(clk_c_enable_524), .CK(clk_c), .Q(rd[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i0.GSR = "DISABLED";
    FD1P3IX instr_len_i1 (.D(n32594), .SP(clk_c_enable_41), .CD(n32840), 
            .CK(clk_c), .Q(instr_len[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_len_i1.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i0 (.D(mem_op_de[0]), .SP(clk_c_enable_365), .CK(clk_c), 
            .Q(mem_op[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i0.GSR = "DISABLED";
    FD1P3AX rs1_i0_i0 (.D(n2632[0]), .SP(clk_c_enable_365), .CK(clk_c), 
            .Q(rs1[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i0.GSR = "DISABLED";
    FD1P3AX data_read_n_i0_i0 (.D(n27629), .SP(clk_c_enable_122), .CK(clk_c), 
            .Q(qv_data_read_n[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_read_n_i0_i0.GSR = "DISABLED";
    LUT4 mux_3051_i10_3_lut_4_lut (.A(\instr[31] ), .B(n32630), .C(n32539), 
         .D(n29738), .Z(n4969[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3051_i10_3_lut_4_lut.init = 16'hf808;
    FD1P3AX instr_data_3__i1 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_309), 
            .CK(clk_c), .Q(\instr_data[3]_adj_13 [0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i1.GSR = "DISABLED";
    FD1S3IX data_ready_sync_415 (.D(data_ready_core), .CK(clk_c), .CD(n32840), 
            .Q(data_ready_sync)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(235[12] 256[8])
    defparam data_ready_sync_415.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i1 (.D(instr_write_offset_3__N_934[0]), .CK(clk_c), 
            .CD(n32840), .Q(\instr_addr_23__N_318[0] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i1.GSR = "DISABLED";
    PFUMX i29 (.BLUT(n11), .ALUT(n13), .C0(n32656), .Z(n16_c));
    PFUMX i13 (.BLUT(n26859), .ALUT(n5), .C0(addr[6]), .Z(n26116));
    FD1P3AX data_continue_420 (.D(data_continue_N_963), .SP(clk_c_enable_52), 
            .CK(clk_c), .Q(debug_data_continue)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_continue_420.GSR = "DISABLED";
    FD1P3IX is_load_393 (.D(is_load_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_load)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_load_393.GSR = "DISABLED";
    PFUMX i29_adj_394 (.BLUT(n9), .ALUT(n12_c), .C0(debug_instr_valid), 
          .Z(n16_adj_3168));
    PFUMX i29176 (.BLUT(n32316), .ALUT(n32314), .C0(counter_hi[4]), .Z(n32317));
    LUT4 i1_4_lut (.A(n32543), .B(n10024), .C(n12_adj_3169), .D(n28527), 
         .Z(n28533)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_rep_708_4_lut (.A(n32851), .B(addr[10]), .C(addr[6]), 
         .D(n32835), .Z(n32723)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_3_lut_rep_708_4_lut.init = 16'hfffd;
    LUT4 i27125_3_lut (.A(\gpio_out_func_sel[5][2] ), .B(\gpio_out_func_sel[7][2] ), 
         .C(addr[3]), .Z(n29834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27125_3_lut.init = 16'hcaca;
    LUT4 mux_2107_i13_3_lut_3_lut (.A(n4271), .B(n3369[11]), .C(n5138[11]), 
         .Z(n3410[12])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2107_i13_3_lut_3_lut.init = 16'he4e4;
    LUT4 i15108_2_lut_3_lut (.A(n31590), .B(n35), .C(n10772), .Z(n3369[0])) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15108_2_lut_3_lut.init = 16'h8080;
    LUT4 i1534_2_lut_3_lut_4_lut_4_lut (.A(\instr_len[2] ), .B(\pc[2] ), 
         .C(\pc[1] ), .D(instr_len[1]), .Z(n2196)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (B+(C (D)+!C !(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1534_2_lut_3_lut_4_lut_4_lut.init = 16'h0990;
    LUT4 i1_3_lut_rep_712_4_lut (.A(n32851), .B(addr[10]), .C(addr[7]), 
         .D(addr[6]), .Z(n32727)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i1_3_lut_rep_712_4_lut.init = 16'hfdff;
    LUT4 i1529_2_lut_3_lut_4_lut_4_lut (.A(\instr_len[2] ), .B(\pc[2] ), 
         .C(\pc[1] ), .D(instr_len[1]), .Z(n2191)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A ((C (D)+!C !(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1529_2_lut_3_lut_4_lut_4_lut.init = 16'h0660;
    LUT4 i1_4_lut_4_lut (.A(n22), .B(n10772), .C(n32640), .D(n4_c), 
         .Z(n27524)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_4_lut_4_lut.init = 16'h0080;
    LUT4 n5568_bdd_3_lut_29222 (.A(counter_hi[2]), .B(instr_data[10]), .C(instr_data[14]), 
         .Z(n32393)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5568_bdd_3_lut_29222.init = 16'he4e4;
    LUT4 i5_2_lut_3_lut (.A(n32548), .B(n32227), .C(additional_mem_ops[2]), 
         .Z(n13456)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(120[15:33])
    defparam i5_2_lut_3_lut.init = 16'h7878;
    LUT4 i30_3_lut_4_lut (.A(n13_adj_3170), .B(n27364), .C(n35), .D(n10772), 
         .Z(n13151)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(47[17:22])
    defparam i30_3_lut_4_lut.init = 16'hcaaa;
    LUT4 n4251_bdd_3_lut_29495 (.A(n29714), .B(n29702), .C(n32734), .Z(n32049)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n4251_bdd_3_lut_29495.init = 16'hacac;
    LUT4 n5568_bdd_3_lut_29230 (.A(counter_hi[2]), .B(\qspi_data_buf[10] ), 
         .C(\qspi_data_buf[14] ), .Z(n32394)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5568_bdd_3_lut_29230.init = 16'he4e4;
    LUT4 i28319_3_lut_4_lut (.A(addr[6]), .B(n32836), .C(addr[7]), .D(addr[3]), 
         .Z(n27888)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i28319_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_4_lut (.A(n32541), .B(n32548), .C(n32191), .D(additional_mem_ops[0]), 
         .Z(additional_mem_ops_2__N_749[0])) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A (B (D)+!B !(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h31ec;
    LUT4 mux_2107_i5_3_lut_4_lut (.A(n3259[4]), .B(n3292[4]), .C(n16_c), 
         .D(n10772), .Z(n3410[4])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2107_i5_3_lut_4_lut.init = 16'hcaaa;
    LUT4 mux_2107_i14_3_lut_3_lut (.A(n4271), .B(n3369[11]), .C(n5138[12]), 
         .Z(n3410[13])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2107_i14_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_2107_i12_3_lut_3_lut (.A(n4271), .B(n3369[11]), .C(n3259[11]), 
         .Z(n3410[11])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2107_i12_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_2107_i8_3_lut_4_lut (.A(n3259[7]), .B(n3292[7]), .C(n16_c), 
         .D(n10772), .Z(n3410[7])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2107_i8_3_lut_4_lut.init = 16'hcaaa;
    LUT4 i27122_3_lut (.A(\gpio_out_func_sel[5][4] ), .B(\gpio_out_func_sel[7][4] ), 
         .C(addr[3]), .Z(n29831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27122_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(n32655), .B(n32659), .C(n34287), .Z(n28547)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4040;
    LUT4 gnd_bdd_2_lut_29153_3_lut_4_lut (.A(addr[6]), .B(n32836), .C(n32252), 
         .D(n32835), .Z(n32253)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam gnd_bdd_2_lut_29153_3_lut_4_lut.init = 16'h0010;
    LUT4 i28612_2_lut_rep_512_3_lut (.A(n16_c), .B(n10772), .C(n19_c), 
         .Z(n32527)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28612_2_lut_rep_512_3_lut.init = 16'hbfbf;
    LUT4 i28552_2_lut_3_lut (.A(n4271), .B(n16_c), .C(n10772), .Z(n30197)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28552_2_lut_3_lut.init = 16'hd5d5;
    LUT4 mux_2107_i17_3_lut_3_lut (.A(n4271), .B(n3369[11]), .C(n5138[15]), 
         .Z(n3410[16])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2107_i17_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_2107_i11_3_lut_3_lut (.A(n4271), .B(n3369[11]), .C(n3259[10]), 
         .Z(n3410[10])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2107_i11_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_3_lut_rep_522_4_lut (.A(n32551), .B(instr_fetch_running), .C(n32544), 
         .D(debug_early_branch), .Z(n32537)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_3_lut_rep_522_4_lut.init = 16'h0002;
    LUT4 mux_2107_i15_3_lut_3_lut (.A(n4271), .B(n3369[11]), .C(n5138[13]), 
         .Z(n3410[14])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2107_i15_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_3151_i31_3_lut_3_lut_4_lut (.A(\instr[31] ), .B(n32630), .C(n29732), 
         .D(n32540), .Z(n5205[30])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3151_i31_3_lut_3_lut_4_lut.init = 16'hf088;
    LUT4 i1_4_lut_adj_395 (.A(debug_early_branch), .B(instr_fetch_running_N_945), 
         .C(n32550), .D(n19867), .Z(n28219)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_395.init = 16'h5010;
    LUT4 i1_4_lut_adj_396 (.A(n2_c), .B(n27851), .C(next_instr_write_offset[3]), 
         .D(n1_c), .Z(n68)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(381[29:75])
    defparam i1_4_lut_adj_396.init = 16'hcc8c;
    FD1S3IX instr_write_offset__i3 (.D(next_instr_write_offset[3]), .CK(clk_c), 
            .CD(n26962), .Q(\instr_write_offset[3] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i3.GSR = "DISABLED";
    LUT4 i1_3_lut_adj_397 (.A(qspi_data_byte_idx[0]), .B(qspi_data_ready), 
         .C(qspi_data_byte_idx[1]), .Z(n27851)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_adj_397.init = 16'hf7f7;
    LUT4 mux_1526_i16_3_lut_then_3_lut (.A(n33[15]), .B(n31[15]), .C(n2150), 
         .Z(n32885)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i16_3_lut_then_3_lut.init = 16'hacac;
    LUT4 mux_1526_i16_3_lut_else_3_lut (.A(n34[15]), .B(n36[15]), .C(n2130), 
         .Z(n32884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i16_3_lut_else_3_lut.init = 16'hcaca;
    LUT4 mux_2107_i16_3_lut_3_lut (.A(n4271), .B(n3369[11]), .C(n5138[14]), 
         .Z(n3410[15])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2107_i16_3_lut_3_lut.init = 16'he4e4;
    FD1S3IX instr_write_offset__i2 (.D(instr_write_offset_3__N_934[1]), .CK(clk_c), 
            .CD(n32840), .Q(instr_addr_23__N_318[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i2.GSR = "DISABLED";
    LUT4 mux_3051_i9_3_lut (.A(n32639), .B(\instr[31] ), .C(n4251), .Z(n4969[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3051_i9_3_lut.init = 16'hcaca;
    LUT4 n5568_bdd_3_lut_29231 (.A(counter_hi[2]), .B(instr_data[11]), .C(instr_data[15]), 
         .Z(n32406)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5568_bdd_3_lut_29231.init = 16'he4e4;
    LUT4 next_pc_for_core_23__I_0_i270_4_lut (.A(n5658[1]), .B(debug_rd_3__N_405[29]), 
         .C(n32785), .D(n9058), .Z(debug_branch_N_446[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i270_4_lut.init = 16'hcac0;
    LUT4 data_from_read_11__bdd_3_lut_then_3_lut (.A(n32685), .B(n19), .C(n32660), 
         .Z(n32897)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam data_from_read_11__bdd_3_lut_then_3_lut.init = 16'hcece;
    LUT4 mux_3051_i8_3_lut (.A(n32656), .B(\instr[31] ), .C(n4251), .Z(n4969[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3051_i8_3_lut.init = 16'hcaca;
    LUT4 n5568_bdd_3_lut_29281 (.A(counter_hi[2]), .B(\qspi_data_buf[11] ), 
         .C(\qspi_data_buf[15] ), .Z(n32407)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5568_bdd_3_lut_29281.init = 16'he4e4;
    LUT4 data_from_read_11__bdd_3_lut_else_3_lut (.A(n32685), .B(n19), .C(\peri_data_out[11] ), 
         .D(n4), .Z(n32896)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam data_from_read_11__bdd_3_lut_else_3_lut.init = 16'heeec;
    LUT4 next_pc_for_core_23__I_0_i271_4_lut (.A(n5658[2]), .B(debug_rd_3__N_405[30]), 
         .C(n32785), .D(n9058), .Z(debug_branch_N_446[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i271_4_lut.init = 16'hcac0;
    LUT4 data_from_read_10__bdd_3_lut_then_3_lut (.A(n32685), .B(n19), .C(n32660), 
         .Z(n32900)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam data_from_read_10__bdd_3_lut_then_3_lut.init = 16'hcece;
    LUT4 data_from_read_10__bdd_3_lut_else_3_lut (.A(n32685), .B(n19), .C(\peri_data_out[10] ), 
         .D(n4), .Z(n32899)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam data_from_read_10__bdd_3_lut_else_3_lut.init = 16'heeec;
    LUT4 mux_3051_i7_3_lut (.A(n32655), .B(\instr[31] ), .C(n4251), .Z(n4969[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3051_i7_3_lut.init = 16'hcaca;
    PFUMX i29151 (.BLUT(n32268), .ALUT(n32267), .C0(n32656), .Z(n32269));
    LUT4 next_pc_for_core_23__I_0_i272_4_lut (.A(n5658[3]), .B(debug_rd_3__N_405[31]), 
         .C(n32785), .D(n9058), .Z(debug_branch_N_446[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i272_4_lut.init = 16'hcac0;
    LUT4 mux_3051_i6_3_lut (.A(n32642), .B(\instr[31] ), .C(n4251), .Z(n4969[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3051_i6_3_lut.init = 16'hcaca;
    FD1P3JX no_write_in_progress_419 (.D(no_write_in_progress_N_471), .SP(clk_c_enable_99), 
            .PD(n32840), .CK(clk_c), .Q(no_write_in_progress)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam no_write_in_progress_419.GSR = "DISABLED";
    LUT4 n32771_bdd_3_lut (.A(counter_hi[2]), .B(\mem_data_from_read[20] ), 
         .C(\mem_data_from_read[16] ), .Z(n33055)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n32771_bdd_3_lut.init = 16'hd8d8;
    LUT4 n33055_bdd_3_lut (.A(n33055), .B(n13_adj_3173), .C(n32771), .Z(n33056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n33055_bdd_3_lut.init = 16'hcaca;
    LUT4 n30322_bdd_3_lut (.A(n30322), .B(n33056), .C(counter_hi[4]), 
         .Z(n33057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30322_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_398 (.A(n32642), .B(n34287), .C(n32641), .D(n32655), 
         .Z(n28641)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_398.init = 16'hc088;
    LUT4 data_from_read_9__bdd_3_lut_then_3_lut (.A(n32685), .B(n19), .C(n32660), 
         .Z(n32859)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam data_from_read_9__bdd_3_lut_then_3_lut.init = 16'hcece;
    LUT4 i1_4_lut_adj_399 (.A(n32651), .B(n34287), .C(n32637), .D(n32655), 
         .Z(n28605)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_399.init = 16'hc088;
    LUT4 mux_1526_i5_3_lut (.A(n29700), .B(n29712), .C(n32734), .Z(instr[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i5_3_lut.init = 16'hcaca;
    LUT4 data_from_read_9__bdd_3_lut_else_3_lut (.A(n32685), .B(n19), .C(\peri_data_out[9] ), 
         .D(n4), .Z(n32858)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam data_from_read_9__bdd_3_lut_else_3_lut.init = 16'heeec;
    FD1P3IX interrupt_core_408 (.D(n32546), .SP(clk_c_enable_545), .CD(n32840), 
            .CK(clk_c), .Q(interrupt_core)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam interrupt_core_408.GSR = "DISABLED";
    LUT4 i28209_3_lut_4_lut (.A(n4267), .B(n4259), .C(n3259[8]), .D(n2970[8]), 
         .Z(n3410[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28209_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_514_3_lut (.A(n32541), .B(n32548), .C(n34287), .Z(clk_c_enable_365)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i1_2_lut_rep_514_3_lut.init = 16'h2020;
    LUT4 mux_2107_i10_3_lut_4_lut (.A(n4267), .B(n4259), .C(n3259[9]), 
         .D(n29723), .Z(n3410[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2107_i10_3_lut_4_lut.init = 16'hf4b0;
    FD1P3IX instr_valid_392 (.D(debug_instr_valid_N_436), .SP(clk_c_enable_545), 
            .CD(n32840), .CK(clk_c), .Q(debug_instr_valid)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_valid_392.GSR = "DISABLED";
    LUT4 i28448_2_lut_3_lut (.A(n32541), .B(n32548), .C(rst_reg_n_adj_6), 
         .Z(clk_c_enable_15)) /* synthesis lut_function=(!(A (B (C))+!A (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i28448_2_lut_3_lut.init = 16'h2f2f;
    LUT4 n31796_bdd_4_lut (.A(n31796), .B(n31795), .C(addr[2]), .D(n32716), 
         .Z(n32520)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n31796_bdd_4_lut.init = 16'hca00;
    PFUMX i29142 (.BLUT(n32254), .ALUT(n32253), .C0(addr[7]), .Z(n32255));
    LUT4 i1_2_lut (.A(qv_data_read_n[0]), .B(qv_data_read_n[1]), .Z(n21414)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i28613_2_lut_3_lut_4_lut (.A(n4267), .B(n4259), .C(n32525), .D(n4271), 
         .Z(n30024)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28613_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 n23_bdd_4_lut (.A(n32656), .B(n32639), .C(n32595), .D(n32654), 
         .Z(n32488)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;
    defparam n23_bdd_4_lut.init = 16'hc800;
    LUT4 pc_3__bdd_3_lut_28777 (.A(\pc[7] ), .B(\pc[15] ), .C(counter_hi[3]), 
         .Z(n31620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_3__bdd_3_lut_28777.init = 16'hcaca;
    LUT4 mux_1526_i11_3_lut (.A(n29727), .B(n2151[10]), .C(n32734), .Z(instr[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i11_3_lut.init = 16'hcaca;
    LUT4 i27133_3_lut_4_lut (.A(n32842), .B(n32841), .C(counter_hi[2]), 
         .D(\next_pc_for_core[6] ), .Z(n29842)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i27133_3_lut_4_lut.init = 16'hf606;
    LUT4 i1_2_lut_adj_400 (.A(n26), .B(n28669), .Z(n28635)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_400.init = 16'h8888;
    LUT4 pc_3__bdd_3_lut_29256 (.A(\pc[3] ), .B(\pc[11] ), .C(counter_hi[3]), 
         .Z(n31621)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_3__bdd_3_lut_29256.init = 16'hcaca;
    LUT4 mux_1526_i7_rep_87_3_lut_3_lut (.A(n32533), .B(n32640), .C(n29716), 
         .Z(n29706)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1526_i7_rep_87_3_lut_3_lut.init = 16'he4e4;
    LUT4 n32191_bdd_3_lut (.A(n32541), .B(n32180), .C(additional_mem_ops[1]), 
         .Z(n33404)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n32191_bdd_3_lut.init = 16'hd8d8;
    LUT4 i1_4_lut_adj_401 (.A(n32642), .B(n34287), .C(n32640), .D(n32655), 
         .Z(n28593)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_401.init = 16'hc088;
    PFUMX i29140 (.BLUT(n32251), .ALUT(n31706), .C0(addr[3]), .Z(n32252));
    LUT4 i1_4_lut_adj_402 (.A(n32642), .B(n34287), .C(n32643), .D(n32655), 
         .Z(n28617)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_402.init = 16'hc088;
    LUT4 mux_347_i2_3_lut_4_lut (.A(n32842), .B(n32841), .C(n32544), .D(return_addr[2]), 
         .Z(n1768[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam mux_347_i2_3_lut_4_lut.init = 16'hf606;
    LUT4 n31622_bdd_3_lut (.A(n31622), .B(n31619), .C(n34281), .Z(debug_branch_N_442[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31622_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_403 (.A(stall_core), .B(clk_c_enable_285), .C(n32771), 
         .D(is_load), .Z(n28957)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_403.init = 16'h8000;
    LUT4 i28266_4_lut (.A(n34285), .B(is_store), .C(no_write_in_progress), 
         .D(is_load), .Z(stall_core)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(149[50:61])
    defparam i28266_4_lut.init = 16'ha0a2;
    LUT4 pc_2__bdd_3_lut_28781 (.A(\pc[6] ), .B(\pc[14] ), .C(counter_hi[3]), 
         .Z(n31625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_2__bdd_3_lut_28781.init = 16'hcaca;
    LUT4 stall_core_I_0_438_2_lut_rep_754 (.A(stall_core), .B(interrupt_core), 
         .Z(n32769)) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(340[19:48])
    defparam stall_core_I_0_438_2_lut_rep_754.init = 16'h1111;
    LUT4 i6367_4_lut_4_lut (.A(n32654), .B(n8330), .C(n30), .D(alu_op_3__N_1170[1]), 
         .Z(n9048)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i6367_4_lut_4_lut.init = 16'hd850;
    LUT4 i1_2_lut_rep_663_3_lut_4_lut_4_lut (.A(stall_core), .B(interrupt_core), 
         .C(n32768), .D(n32849), .Z(n32678)) /* synthesis lut_function=((B+!((D)+!C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(340[19:48])
    defparam i1_2_lut_rep_663_3_lut_4_lut_4_lut.init = 16'hddfd;
    PFUMX i29130 (.BLUT(n32226), .ALUT(n32225), .C0(clk_c_enable_41), 
          .Z(n32227));
    LUT4 pc_2__bdd_3_lut_29250 (.A(\pc[2] ), .B(\pc[10] ), .C(counter_hi[3]), 
         .Z(n31626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_2__bdd_3_lut_29250.init = 16'hcaca;
    LUT4 n30920_bdd_4_lut (.A(n30920), .B(n32656), .C(n32654), .D(n32655), 
         .Z(n32494)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam n30920_bdd_4_lut.init = 16'h0204;
    LUT4 n32191_bdd_2_lut (.A(additional_mem_ops[1]), .B(additional_mem_ops[0]), 
         .Z(n33403)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam n32191_bdd_2_lut.init = 16'h9999;
    LUT4 n31627_bdd_3_lut (.A(n31627), .B(n31624), .C(n34281), .Z(debug_branch_N_442[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31627_bdd_3_lut.init = 16'hcaca;
    LUT4 n30920_bdd_3_lut (.A(n30920), .B(n32656), .C(n32655), .Z(n32493)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;
    defparam n30920_bdd_3_lut.init = 16'h4545;
    PFUMX i10 (.BLUT(n26857), .ALUT(n21), .C0(addr[6]), .Z(n3));
    LUT4 mux_1526_i8_rep_85_3_lut_3_lut (.A(n32533), .B(n32641), .C(n29718), 
         .Z(n29704)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1526_i8_rep_85_3_lut_3_lut.init = 16'he4e4;
    LUT4 i28181_3_lut_4_lut (.A(n13140), .B(n32643), .C(n4265), .D(n27489), 
         .Z(n3369[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i28181_3_lut_4_lut.init = 16'hf808;
    PFUMX i29128 (.BLUT(n32222), .ALUT(n32221), .C0(n32654), .Z(n32223));
    PFUMX i8 (.BLUT(n26858), .ALUT(n20), .C0(addr[6]), .Z(n3_adj_7));
    LUT4 i1_4_lut_adj_404 (.A(n32642), .B(n34287), .C(n32638), .D(n32655), 
         .Z(n28653)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_404.init = 16'hc088;
    LUT4 i28171_3_lut_4_lut (.A(n32638), .B(n13140), .C(n4265), .D(n27480), 
         .Z(n3183[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i28171_3_lut_4_lut.init = 16'hf808;
    LUT4 i27755_3_lut (.A(imm_c[25]), .B(imm_c[29]), .C(counter_hi[2]), 
         .Z(n30464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27755_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_405 (.A(n10024), .B(n28791), .C(n32566), .D(n32573), 
         .Z(n28797)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_405.init = 16'h0004;
    FD1P3IX is_system_402 (.D(is_system_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_system)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_system_402.GSR = "DISABLED";
    LUT4 mux_1526_i8_3_lut (.A(n29707), .B(n29718), .C(n32734), .Z(instr[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i8_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32656), .B(n32655), .C(n32661), .D(n32639), 
         .Z(n24898)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3AX data_write_n_i0 (.D(data_write_n_1__N_369[0]), .SP(clk_c_enable_513), 
            .CK(clk_c), .Q(qv_data_write_n[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_write_n_i0.GSR = "DISABLED";
    FD1P3AX data_read_n_i0_i1 (.D(n27630), .SP(clk_c_enable_122), .CK(clk_c), 
            .Q(qv_data_read_n[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_read_n_i0_i1.GSR = "DISABLED";
    FD1P3AX rs1_i0_i3 (.D(n2632[3]), .SP(clk_c_enable_365), .CK(clk_c), 
            .Q(rs1[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i3.GSR = "DISABLED";
    FD1P3AX rs1_i0_i2 (.D(n2632[2]), .SP(clk_c_enable_365), .CK(clk_c), 
            .Q(rs1[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i2.GSR = "DISABLED";
    FD1P3AX rs1_i0_i1 (.D(n2632[1]), .SP(clk_c_enable_365), .CK(clk_c), 
            .Q(rs1[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i1.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i2 (.D(mem_op_de[2]), .SP(clk_c_enable_365), .CK(clk_c), 
            .Q(mem_op[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i2.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i1 (.D(mem_op_de[1]), .SP(clk_c_enable_365), .CK(clk_c), 
            .Q(mem_op[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i1.GSR = "DISABLED";
    FD1P3AX instr_len_i2 (.D(n32588), .SP(clk_c_enable_338), .CK(clk_c), 
            .Q(\instr_len[2] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_len_i2.GSR = "DISABLED";
    FD1P3AX rd_i0_i3 (.D(n6[3]), .SP(clk_c_enable_524), .CK(clk_c), .Q(rd_c[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i3.GSR = "DISABLED";
    FD1P3AX rd_i0_i2 (.D(n6[2]), .SP(clk_c_enable_524), .CK(clk_c), .Q(rd_c[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i2.GSR = "DISABLED";
    FD1P3AX rd_i0_i1 (.D(n6[1]), .SP(clk_c_enable_524), .CK(clk_c), .Q(rd_c[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_586_3_lut (.A(n32656), .B(n32655), .C(n32639), .Z(n32601)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_586_3_lut.init = 16'h8080;
    LUT4 i1_3_lut_3_lut (.A(n32548), .B(n32877), .C(n10024), .Z(n28343)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_3_lut_3_lut.init = 16'h0404;
    LUT4 n10904_bdd_2_lut_29274_3_lut_4_lut (.A(n32656), .B(n32655), .C(n32657), 
         .D(n32639), .Z(n32177)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam n10904_bdd_2_lut_29274_3_lut_4_lut.init = 16'h8000;
    LUT4 n32308_bdd_3_lut_4_lut (.A(addr[27]), .B(n32850), .C(n13_adj_3173), 
         .D(n32308), .Z(n32309)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n32308_bdd_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX data_addr__i27 (.D(addr_out[27]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(addr[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i27.GSR = "DISABLED";
    FD1P3IX data_addr__i26 (.D(addr_out[26]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(addr_c[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i26.GSR = "DISABLED";
    FD1P3IX data_addr__i25 (.D(addr_out[25]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(addr_c[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i25.GSR = "DISABLED";
    FD1P3IX data_addr__i24 (.D(addr_out[24]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[24] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i24.GSR = "DISABLED";
    FD1P3IX data_addr__i23 (.D(addr_out[23]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i23.GSR = "DISABLED";
    FD1P3IX data_addr__i22 (.D(addr_out[22]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i22.GSR = "DISABLED";
    FD1P3IX data_addr__i21 (.D(addr_out[21]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i21.GSR = "DISABLED";
    LUT4 i31_4_lut_4_lut (.A(n32639), .B(n32656), .C(n26863), .D(n32655), 
         .Z(n25)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(C+(D))))) */ ;
    defparam i31_4_lut_4_lut.init = 16'h11fc;
    LUT4 i27754_3_lut (.A(imm[17]), .B(\imm[21] ), .C(counter_hi[2]), 
         .Z(n30463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27754_3_lut.init = 16'hcaca;
    LUT4 i27753_3_lut (.A(\imm[9] ), .B(\imm[13] ), .C(counter_hi[2]), 
         .Z(n30462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27753_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_406 (.A(n10024), .B(n28763), .C(n32566), .D(n32573), 
         .Z(n28769)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_406.init = 16'h0004;
    LUT4 i27752_3_lut (.A(\imm[1] ), .B(\imm[5] ), .C(counter_hi[2]), 
         .Z(n30461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27752_3_lut.init = 16'hcaca;
    LUT4 i52_4_lut_4_lut (.A(n32654), .B(n32655), .C(n17747), .D(n32656), 
         .Z(n37)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (D)+!B !(C+(D))))) */ ;
    defparam i52_4_lut_4_lut.init = 16'h4403;
    LUT4 i27748_3_lut (.A(imm_c[24]), .B(imm_c[28]), .C(counter_hi[2]), 
         .Z(n30457)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27748_3_lut.init = 16'hcaca;
    LUT4 i27747_3_lut (.A(imm[16]), .B(\imm[20] ), .C(counter_hi[2]), 
         .Z(n30456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27747_3_lut.init = 16'hcaca;
    LUT4 mux_1526_i7_3_lut (.A(n29710), .B(n29716), .C(n32734), .Z(instr[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i7_3_lut.init = 16'hcaca;
    LUT4 n32395_bdd_3_lut_4_lut (.A(addr[27]), .B(n32850), .C(n32901), 
         .D(n32395), .Z(n30365)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n32395_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32408_bdd_3_lut_4_lut (.A(addr[27]), .B(n32850), .C(n32898), 
         .D(n32408), .Z(n32409)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n32408_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_407 (.A(n10024), .B(n28805), .C(n32566), .D(n32573), 
         .Z(n28811)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_407.init = 16'h0004;
    LUT4 mux_1526_i6_3_lut (.A(n29702), .B(n29714), .C(n32734), .Z(instr[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i6_3_lut.init = 16'hcaca;
    LUT4 i27746_3_lut (.A(\imm[8] ), .B(\imm[12] ), .C(counter_hi[2]), 
         .Z(n30455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27746_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n32548), .B(n32543), .C(n28539), .D(n32546), 
         .Z(n2792)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i27745_3_lut (.A(imm_c[0]), .B(\imm[4] ), .C(counter_hi[2]), 
         .Z(n30454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27745_3_lut.init = 16'hcaca;
    LUT4 i27128_3_lut (.A(\next_pc_for_core[9] ), .B(\next_pc_for_core[13] ), 
         .C(counter_hi[2]), .Z(n29837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27128_3_lut.init = 16'hcaca;
    FD1P3IX data_addr__i20 (.D(addr_out[20]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i20.GSR = "DISABLED";
    FD1P3IX data_addr__i19 (.D(addr_out[19]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i19.GSR = "DISABLED";
    FD1P3IX data_addr__i18 (.D(addr_out[18]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i18.GSR = "DISABLED";
    FD1P3IX data_addr__i17 (.D(addr_out[17]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[17] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i17.GSR = "DISABLED";
    LUT4 i15527_2_lut_3_lut_4_lut (.A(n32654), .B(n32656), .C(n32655), 
         .D(n32639), .Z(n30)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i15527_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i28290_2_lut_rep_584_3_lut (.A(n32654), .B(n32656), .C(n32639), 
         .Z(n32599)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i28290_2_lut_rep_584_3_lut.init = 16'h1010;
    FD1P3IX data_addr__i16 (.D(addr_out[16]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[16] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i16.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_408 (.A(n10024), .B(n28777), .C(n32566), .D(n32573), 
         .Z(n28783)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_408.init = 16'h0004;
    LUT4 pc_1__bdd_3_lut_28801 (.A(\pc[5] ), .B(\pc[13] ), .C(counter_hi[3]), 
         .Z(n31650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_1__bdd_3_lut_28801.init = 16'hcaca;
    FD1P3IX data_addr__i15 (.D(addr_out[15]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[15] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i15.GSR = "DISABLED";
    LUT4 i1_3_lut_adj_409 (.A(no_write_in_progress), .B(debug_instr_valid), 
         .C(is_store), .Z(debug_rd_3__N_413)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_3_lut_adj_409.init = 16'h8080;
    LUT4 i49_3_lut_3_lut (.A(n32654), .B(n32656), .C(n32653), .Z(n28)) /* synthesis lut_function=(!(A (C)+!A (B+!(C)))) */ ;
    defparam i49_3_lut_3_lut.init = 16'h1a1a;
    LUT4 i28587_3_lut_4_lut (.A(addr[27]), .B(n32850), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n30160)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i28587_3_lut_4_lut.init = 16'hefff;
    LUT4 pc_1__bdd_3_lut_29234 (.A(\pc[1] ), .B(\pc[9] ), .C(counter_hi[3]), 
         .Z(n31651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_1__bdd_3_lut_29234.init = 16'hcaca;
    FD1P3IX data_addr__i14 (.D(addr_out[14]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[14] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i14.GSR = "DISABLED";
    FD1P3IX data_addr__i13 (.D(addr_out[13]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[13] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i13.GSR = "DISABLED";
    FD1P3IX data_addr__i12 (.D(addr_out[12]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[12] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i12.GSR = "DISABLED";
    FD1P3IX data_addr__i11 (.D(addr_out[11]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[11] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i11.GSR = "DISABLED";
    FD1P3IX data_addr__i10 (.D(addr_out[10]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(addr[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i10.GSR = "DISABLED";
    FD1P3IX data_addr__i9 (.D(addr_out[9]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[9] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i9.GSR = "DISABLED";
    FD1P3IX data_addr__i8 (.D(addr_out[8]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[8] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i8.GSR = "DISABLED";
    FD1P3IX data_addr__i7 (.D(addr_out[7]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(addr[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i7.GSR = "DISABLED";
    FD1P3IX data_addr__i6 (.D(addr_out[6]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(addr[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i6.GSR = "DISABLED";
    FD1P3IX data_addr__i5 (.D(addr_out[5]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[5] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i5.GSR = "DISABLED";
    FD1P3IX data_addr__i4 (.D(addr_out[4]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[4] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i4.GSR = "DISABLED";
    FD1S3IX counter_hi_3544__i2 (.D(n32812), .CK(clk_c), .CD(n32840), 
            .Q(counter_hi[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3544__i2.GSR = "DISABLED";
    FD1P3IX data_addr__i3 (.D(n27823), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(addr[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i3.GSR = "DISABLED";
    FD1P3IX data_addr__i2 (.D(n699[0]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(addr[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i2.GSR = "DISABLED";
    FD1P3IX data_addr__i1 (.D(addr_out[1]), .SP(clk_c_enable_174), .CD(n32840), 
            .CK(clk_c), .Q(\addr[1] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i1.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i2 (.D(additional_mem_ops_2__N_749[2]), .CK(clk_c), 
            .CD(n32840), .Q(additional_mem_ops[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i2.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i1 (.D(additional_mem_ops_2__N_749[1]), .CK(clk_c), 
            .CD(n32840), .Q(additional_mem_ops[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i1.GSR = "DISABLED";
    FD1P3IX data_out__i31 (.D(n32644), .SP(clk_c_enable_178), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i31.GSR = "DISABLED";
    FD1P3IX data_out__i30 (.D(data_out_slice[2]), .SP(clk_c_enable_178), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i30.GSR = "DISABLED";
    FD1S3IX addr_offset_3545__i2 (.D(n38[0]), .CK(clk_c), .CD(n32840), 
            .Q(addr_offset[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam addr_offset_3545__i2.GSR = "DISABLED";
    FD1P3IX data_out__i29 (.D(n32668), .SP(clk_c_enable_178), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i29.GSR = "DISABLED";
    FD1P3IX data_out__i28 (.D(data_out_slice[0]), .SP(clk_c_enable_178), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i28.GSR = "DISABLED";
    FD1P3IX data_out__i27 (.D(n32644), .SP(clk_c_enable_182), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i27.GSR = "DISABLED";
    FD1P3IX data_out__i26 (.D(data_out_slice[2]), .SP(clk_c_enable_182), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i26.GSR = "DISABLED";
    FD1P3IX data_out__i25 (.D(n32668), .SP(clk_c_enable_182), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i25.GSR = "DISABLED";
    FD1P3IX data_out__i24 (.D(data_out_slice[0]), .SP(clk_c_enable_182), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i24.GSR = "DISABLED";
    LUT4 i15161_2_lut (.A(\next_pc_for_core[4] ), .B(counter_hi[2]), .Z(n149)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i15161_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_410 (.A(addr[27]), .B(n32850), .C(n12), 
         .D(n21414), .Z(data_ready_r_N_2823)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_4_lut_adj_410.init = 16'h00e0;
    FD1P3IX data_out__i23 (.D(n32644), .SP(clk_c_enable_187), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[23])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i23.GSR = "DISABLED";
    FD1P3IX data_out__i22 (.D(data_out_slice[2]), .SP(clk_c_enable_187), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[22])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i22.GSR = "DISABLED";
    FD1P3IX data_out__i21 (.D(n32668), .SP(clk_c_enable_187), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[21])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i21.GSR = "DISABLED";
    FD1P3IX data_out__i20 (.D(data_out_slice[0]), .SP(clk_c_enable_187), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[20])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i20.GSR = "DISABLED";
    FD1P3IX data_out__i19 (.D(n32644), .SP(clk_c_enable_191), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[19])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i19.GSR = "DISABLED";
    FD1P3IX data_out__i18 (.D(data_out_slice[2]), .SP(clk_c_enable_191), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[18])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i18.GSR = "DISABLED";
    FD1P3IX data_out__i17 (.D(n32668), .SP(clk_c_enable_191), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[17])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i17.GSR = "DISABLED";
    FD1P3IX data_out__i16 (.D(data_out_slice[0]), .SP(clk_c_enable_191), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[16])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i16.GSR = "DISABLED";
    PFUMX i29112 (.BLUT(n32190), .ALUT(n32189), .C0(n32653), .Z(n32191));
    LUT4 i1_2_lut_3_lut_4_lut_adj_411 (.A(addr[27]), .B(n32850), .C(data_ready_r), 
         .D(n32801), .Z(n29059)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_4_lut_adj_411.init = 16'hf0fe;
    LUT4 data_from_read_6__bdd_4_lut (.A(n32598), .B(data_txn_len[0]), .C(instr_data[14]), 
         .D(instr_data[6]), .Z(n32990)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam data_from_read_6__bdd_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_rep_554_4_lut (.A(n32639), .B(n32655), .C(n32656), .D(n29681), 
         .Z(n32569)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_3_lut_rep_554_4_lut.init = 16'h0002;
    LUT4 n31652_bdd_3_lut (.A(n31652), .B(n31649), .C(n34281), .Z(debug_branch_N_442[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31652_bdd_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut (.A(n32653), .B(n32654), .C(n32639), .Z(n11)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_2_lut_3_lut.init = 16'h2020;
    LUT4 i2_2_lut_3_lut_adj_412 (.A(n32653), .B(n32654), .C(n32655), .Z(n17)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_2_lut_3_lut_adj_412.init = 16'h2020;
    LUT4 i1_3_lut_rep_699_4_lut (.A(addr[27]), .B(n32850), .C(n32801), 
         .D(n21414), .Z(n32714)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_3_lut_rep_699_4_lut.init = 16'hfeee;
    LUT4 n32384_bdd_3_lut_4_lut (.A(addr[27]), .B(n32850), .C(n32860), 
         .D(n32384), .Z(n32385)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n32384_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32313_bdd_3_lut_4_lut (.A(addr[27]), .B(n32850), .C(n13_adj_3173), 
         .D(n32313), .Z(n32314)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n32313_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15012_2_lut_3_lut (.A(n32653), .B(n32654), .C(n32362), .Z(mem_op_de[0])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i15012_2_lut_3_lut.init = 16'hd0d0;
    FD1P3IX data_out__i15 (.D(n32644), .SP(clk_c_enable_195), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i15.GSR = "DISABLED";
    FD1P3IX data_out__i14 (.D(data_out_slice[2]), .SP(clk_c_enable_195), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i14.GSR = "DISABLED";
    FD1P3IX data_out__i13 (.D(n32668), .SP(clk_c_enable_195), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i13.GSR = "DISABLED";
    FD1P3IX data_out__i12 (.D(data_out_slice[0]), .SP(clk_c_enable_195), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i12.GSR = "DISABLED";
    LUT4 i1_rep_516_4_lut (.A(debug_early_branch), .B(n32544), .C(n32550), 
         .D(n32689), .Z(n32531)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_rep_516_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_4_lut_adj_413 (.A(n32851), .B(addr[10]), .C(rst_reg_n), 
         .D(n32706), .Z(n15569)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_413.init = 16'hd000;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n32854), .B(counter_hi[4]), .C(debug_instr_valid), 
         .D(n27294), .Z(n28851)) /* synthesis lut_function=(A (B ((D)+!C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h8808;
    FD1P3IX data_out__i11 (.D(n32644), .SP(clk_c_enable_200), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i11.GSR = "DISABLED";
    PFUMX i29107 (.BLUT(n32177), .ALUT(n32176), .C0(n32653), .Z(n32178));
    FD1P3IX data_out__i10 (.D(data_out_slice[2]), .SP(clk_c_enable_200), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i10.GSR = "DISABLED";
    FD1P3IX data_out__i9 (.D(n32668), .SP(clk_c_enable_200), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i9.GSR = "DISABLED";
    FD1P3IX data_out__i8 (.D(data_out_slice[0]), .SP(clk_c_enable_200), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i8.GSR = "DISABLED";
    L6MUX21 i29387 (.D0(n32993), .D1(n32991), .SD(counter_hi[2]), .Z(n32994));
    FD1P3IX data_out__i7 (.D(n32644), .SP(clk_c_enable_204), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i7.GSR = "DISABLED";
    FD1P3IX data_out__i6 (.D(data_out_slice[2]), .SP(clk_c_enable_204), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i6.GSR = "DISABLED";
    FD1P3IX data_out__i5 (.D(n32668), .SP(clk_c_enable_204), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i5.GSR = "DISABLED";
    FD1P3IX data_out__i4 (.D(data_out_slice[0]), .SP(clk_c_enable_204), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i4.GSR = "DISABLED";
    FD1P3IX data_out__i3 (.D(n32644), .SP(clk_c_enable_207), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i3.GSR = "DISABLED";
    FD1P3IX data_out__i2 (.D(data_out_slice[2]), .SP(clk_c_enable_207), 
            .CD(n32840), .CK(clk_c), .Q(data_to_write[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i2.GSR = "DISABLED";
    FD1P3IX data_out__i1 (.D(n32668), .SP(clk_c_enable_207), .CD(n32840), 
            .CK(clk_c), .Q(data_to_write[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i1.GSR = "DISABLED";
    LUT4 i4374_2_lut_rep_761 (.A(rd_c[1]), .B(rd[0]), .Z(n32776)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(180[19:31])
    defparam i4374_2_lut_rep_761.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(rd_c[1]), .B(rd[0]), .C(n32783), .D(rd_c[2]), 
         .Z(n28909)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)))+!A !(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(180[19:31])
    defparam i1_3_lut_4_lut.init = 16'h7080;
    LUT4 i27018_3_lut_4_lut (.A(n32658), .B(n32657), .C(n32641), .D(n32642), 
         .Z(n29661)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i27018_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_414 (.A(n32658), .B(n32657), .C(n32661), .D(n32642), 
         .Z(n29031)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_414.init = 16'hfffe;
    LUT4 n2122_bdd_4_lut_29733 (.A(n32538), .B(n2211), .C(n17165), .D(n32734), 
         .Z(n33737)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;
    defparam n2122_bdd_4_lut_29733.init = 16'hfaee;
    LUT4 n2122_bdd_4_lut (.A(n4_adj_3177), .B(n32546), .C(n28453), .D(n32543), 
         .Z(n33738)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam n2122_bdd_4_lut.init = 16'h2000;
    LUT4 n2124_bdd_4_lut (.A(n2211), .B(n17165), .C(n32734), .D(n32653), 
         .Z(n33735)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n2124_bdd_4_lut.init = 16'hffca;
    FD1P3IX is_branch_399 (.D(is_branch_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_branch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_branch_399.GSR = "DISABLED";
    FD1P3IX load_started_422 (.D(VCC_net), .SP(address_ready), .CD(n829), 
            .CK(clk_c), .Q(load_started)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam load_started_422.GSR = "DISABLED";
    LUT4 i24592_4_lut (.A(n32694), .B(n7), .C(n26988), .D(n8854), .Z(n13_adj_3173)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam i24592_4_lut.init = 16'hcddd;
    LUT4 i27134_3_lut (.A(\next_pc_for_core[10] ), .B(\next_pc_for_core[14] ), 
         .C(counter_hi[2]), .Z(n29843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27134_3_lut.init = 16'hcaca;
    LUT4 i27716_3_lut (.A(n30423), .B(n32409), .C(counter_hi[3]), .Z(n30425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27716_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_rep_525 (.A(n32543), .B(n32546), .C(n32548), .D(n28505), 
         .Z(n32540)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_rep_525.init = 16'h0200;
    LUT4 i27620_3_lut (.A(n30327), .B(n32385), .C(counter_hi[3]), .Z(n30329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27620_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_768 (.A(additional_mem_ops[1]), .B(additional_mem_ops[0]), 
         .C(additional_mem_ops[2]), .Z(n32783)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_768.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_415 (.A(n32543), .B(n32546), .C(n10024), .D(n27653), 
         .Z(clk_c_enable_364)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_415.init = 16'h0002;
    LUT4 i1_2_lut_4_lut_adj_416 (.A(additional_mem_ops[1]), .B(additional_mem_ops[0]), 
         .C(additional_mem_ops[2]), .D(n34287), .Z(n28889)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_416.init = 16'hfe00;
    LUT4 next_pc_for_core_23__I_0_i269_4_lut (.A(n209), .B(n32351), .C(n32741), 
         .D(n9058), .Z(debug_branch_N_446[28])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i269_4_lut.init = 16'haca0;
    FD1P3AX instr_data_3__i64 (.D(instr_data[15]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i64.GSR = "DISABLED";
    FD1P3AX instr_data_3__i63 (.D(instr_data[14]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i63.GSR = "DISABLED";
    FD1P3AX instr_data_3__i62 (.D(instr_data[13]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i62.GSR = "DISABLED";
    FD1P3AX instr_data_3__i61 (.D(instr_data[12]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i61.GSR = "DISABLED";
    FD1P3AX instr_data_3__i60 (.D(instr_data[11]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i60.GSR = "DISABLED";
    FD1P3AX instr_data_3__i59 (.D(instr_data[10]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i59.GSR = "DISABLED";
    FD1P3AX instr_data_3__i58 (.D(instr_data[9]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i58.GSR = "DISABLED";
    FD1P3AX instr_data_3__i57 (.D(instr_data[8]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i57.GSR = "DISABLED";
    FD1P3AX instr_data_3__i56 (.D(instr_data[7]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i56.GSR = "DISABLED";
    FD1P3AX instr_data_3__i55 (.D(instr_data[6]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i55.GSR = "DISABLED";
    FD1P3AX instr_data_3__i54 (.D(instr_data[5]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i54.GSR = "DISABLED";
    FD1P3AX instr_data_3__i53 (.D(instr_data[4]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i53.GSR = "DISABLED";
    FD1P3AX instr_data_3__i52 (.D(instr_data[3]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i52.GSR = "DISABLED";
    FD1P3AX instr_data_3__i51 (.D(instr_data[2]), .SP(clk_c_enable_232), 
            .CK(clk_c), .Q(n33[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i51.GSR = "DISABLED";
    LUT4 i1_rep_520_4_lut (.A(n32543), .B(n32546), .C(n10024), .D(n32548), 
         .Z(clk_c_enable_41)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_rep_520_4_lut.init = 16'h0002;
    LUT4 i14916_4_lut_4_lut (.A(n32544), .B(n68), .C(n28219), .D(n32714), 
         .Z(debug_stop_txn_N_2142)) /* synthesis lut_function=(!(A (B+(D))+!A !(B (C)+!B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(435[108:115])
    defparam i14916_4_lut_4_lut.init = 16'h5073;
    LUT4 is_lui_I_0_473_2_lut_rep_770 (.A(is_lui), .B(debug_instr_valid), 
         .Z(n32785)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam is_lui_I_0_473_2_lut_rep_770.init = 16'h8888;
    FD1P3AX instr_data_3__i50 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_234), 
            .CK(clk_c), .Q(n33[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i50.GSR = "DISABLED";
    FD1P3AX instr_data_3__i49 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_234), 
            .CK(clk_c), .Q(\instr_data[0][0] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i49.GSR = "DISABLED";
    FD1P3AX instr_data_3__i48 (.D(instr_data[15]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i48.GSR = "DISABLED";
    FD1P3AX instr_data_3__i47 (.D(instr_data[14]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i47.GSR = "DISABLED";
    FD1P3AX instr_data_3__i46 (.D(instr_data[13]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i46.GSR = "DISABLED";
    FD1P3AX instr_data_3__i45 (.D(instr_data[12]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i45.GSR = "DISABLED";
    FD1P3AX instr_data_3__i44 (.D(instr_data[11]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i44.GSR = "DISABLED";
    FD1P3AX instr_data_3__i43 (.D(instr_data[10]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i43.GSR = "DISABLED";
    FD1P3AX instr_data_3__i42 (.D(instr_data[9]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i42.GSR = "DISABLED";
    FD1P3AX instr_data_3__i41 (.D(instr_data[8]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i41.GSR = "DISABLED";
    FD1P3AX instr_data_3__i40 (.D(instr_data[7]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(\instr_data[1][7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i40.GSR = "DISABLED";
    FD1P3AX instr_data_3__i39 (.D(instr_data[6]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i39.GSR = "DISABLED";
    FD1P3AX instr_data_3__i38 (.D(instr_data[5]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i38.GSR = "DISABLED";
    FD1P3AX instr_data_3__i37 (.D(instr_data[4]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i37.GSR = "DISABLED";
    FD1P3AX instr_data_3__i36 (.D(instr_data[3]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i36.GSR = "DISABLED";
    FD1P3AX instr_data_3__i35 (.D(instr_data[2]), .SP(clk_c_enable_248), 
            .CK(clk_c), .Q(n34[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i35.GSR = "DISABLED";
    FD1P3AX instr_data_3__i34 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_250), 
            .CK(clk_c), .Q(n34[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i34.GSR = "DISABLED";
    FD1P3AX instr_data_3__i33 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_250), 
            .CK(clk_c), .Q(\instr_data[1][0] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i33.GSR = "DISABLED";
    FD1P3AX instr_data_3__i32 (.D(instr_data[15]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i32.GSR = "DISABLED";
    FD1P3AX instr_data_3__i31 (.D(instr_data[14]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i31.GSR = "DISABLED";
    FD1P3AX instr_data_3__i30 (.D(instr_data[13]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i30.GSR = "DISABLED";
    FD1P3AX instr_data_3__i29 (.D(instr_data[12]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i29.GSR = "DISABLED";
    FD1P3AX instr_data_3__i28 (.D(instr_data[11]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i28.GSR = "DISABLED";
    FD1P3AX instr_data_3__i27 (.D(instr_data[10]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i27.GSR = "DISABLED";
    FD1P3AX instr_data_3__i26 (.D(instr_data[9]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i26.GSR = "DISABLED";
    FD1P3AX instr_data_3__i25 (.D(instr_data[8]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i25.GSR = "DISABLED";
    FD1P3AX instr_data_3__i24 (.D(instr_data[7]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(\instr_data[2][7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i24.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_527 (.A(data_stall), .B(n19867), .Z(n32542)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_527.init = 16'heeee;
    LUT4 i27463_3_lut_4_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(n30179), 
         .D(n32784), .Z(n30172)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i27463_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 next_pc_for_core_23__I_0_i157_3_lut (.A(\next_pc_for_core[8] ), .B(\next_pc_for_core[12] ), 
         .C(counter_hi[2]), .Z(n157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i157_3_lut.init = 16'hcaca;
    LUT4 i28595_3_lut_4_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(n32808), 
         .D(n32784), .Z(n30070)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i28595_3_lut_4_lut_4_lut.init = 16'hc888;
    LUT4 i28566_2_lut_3_lut_4_lut_4_lut (.A(is_lui), .B(debug_instr_valid), 
         .C(is_jalr), .D(is_jal), .Z(n30175)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i28566_2_lut_3_lut_4_lut_4_lut.init = 16'hbbbf;
    LUT4 mux_91_i1_3_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(debug_rd_3__N_405[28]), 
         .D(n157), .Z(n234[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam mux_91_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_772 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n32787)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_2_lut_rep_772.init = 16'h2222;
    LUT4 mux_105_i1_3_lut_4_lut (.A(data_stall), .B(n19867), .C(n32740), 
         .D(data_req_N_2334), .Z(n332)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_105_i1_3_lut_4_lut.init = 16'hf101;
    LUT4 i1_2_lut_rep_727_3_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(instr_active), .Z(n32742)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_2_lut_rep_727_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_417 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(qspi_data_ready), .D(instr_active), .Z(n28511)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_2_lut_3_lut_4_lut_adj_417.init = 16'h0200;
    LUT4 mux_1539_i5_3_lut (.A(n33[4]), .B(n34[4]), .C(n2130), .Z(n2202[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i5_3_lut.init = 16'hcaca;
    LUT4 i28370_2_lut_rep_570_3_lut_4_lut (.A(n32654), .B(n32639), .C(n32655), 
         .D(n32656), .Z(n32585)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i28370_2_lut_rep_570_3_lut_4_lut.init = 16'h0001;
    LUT4 mux_1549_i2_rep_133_3_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .Z(n30919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i2_rep_133_3_lut.init = 16'hcaca;
    LUT4 mux_1543_i5_3_lut (.A(n36[4]), .B(n31[4]), .C(n2150), .Z(n2222[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i5_3_lut.init = 16'hcaca;
    LUT4 i28478_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n11193), .D(qspi_data_ready), .Z(clk_c_enable_91)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i28478_3_lut_4_lut.init = 16'h20f0;
    LUT4 i27049_3_lut (.A(\mem_data_from_read[19] ), .B(\mem_data_from_read[23] ), 
         .C(counter_hi[2]), .Z(n29758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27049_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_2_lut_rep_773 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n32788)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_3_lut_2_lut_rep_773.init = 16'h6666;
    LUT4 i15009_4_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(txn_len[1]), .D(n1), .Z(n175)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i15009_4_lut_4_lut.init = 16'h6624;
    LUT4 i30_3_lut_4_lut_3_lut (.A(n32654), .B(n32639), .C(n32653), .Z(n13)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam i30_3_lut_4_lut_3_lut.init = 16'h1818;
    LUT4 i1_2_lut_rep_774 (.A(\read_cycles_count[1] ), .B(data_stall), .Z(n32789)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_774.init = 16'heeee;
    LUT4 i28365_2_lut_3_lut (.A(\read_cycles_count[1] ), .B(data_stall), 
         .C(n19867), .Z(data_ready_N_2347)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i28365_2_lut_3_lut.init = 16'h0101;
    FD1P3IX is_jalr_400 (.D(is_jalr_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_jalr)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_jalr_400.GSR = "DISABLED";
    PFUMX mux_1526_i4 (.BLUT(n2131[3]), .ALUT(n2151[3]), .C0(n32734), 
          .Z(instr[19]));
    PFUMX mux_1526_i9 (.BLUT(n2131[8]), .ALUT(n2151[8]), .C0(n32734), 
          .Z(instr[24]));
    LUT4 debug_branch_I_48_i1_3_lut (.A(n29840), .B(load_top_bit), .C(data_out_3__N_1385), 
         .Z(debug_branch_N_450[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_48_i1_3_lut.init = 16'hcaca;
    PFUMX mux_1526_i10 (.BLUT(n2131[9]), .ALUT(n2151[9]), .C0(n32734), 
          .Z(instr[25]));
    PFUMX mux_1526_i13 (.BLUT(n2131[12]), .ALUT(n2151[12]), .C0(n32734), 
          .Z(instr[28]));
    PFUMX mux_1526_i14 (.BLUT(n2131[13]), .ALUT(n2151[13]), .C0(n32734), 
          .Z(instr[29]));
    LUT4 debug_branch_I_48_i2_3_lut (.A(n29858), .B(load_top_bit), .C(data_out_3__N_1385), 
         .Z(debug_branch_N_450[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_48_i2_3_lut.init = 16'hcaca;
    LUT4 i28438_3_lut_4_lut (.A(n32563), .B(n32734), .C(n32540), .D(n32525), 
         .Z(n29917)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28438_3_lut_4_lut.init = 16'h10ff;
    LUT4 i28422_3_lut_4_lut (.A(n32563), .B(n32734), .C(n32540), .D(n32525), 
         .Z(n29960)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28422_3_lut_4_lut.init = 16'h1fff;
    LUT4 n32052_bdd_3_lut_4_lut (.A(n32563), .B(n32643), .C(n32540), .D(n32052), 
         .Z(n32053)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n32052_bdd_3_lut_4_lut.init = 16'h8f80;
    FD1P3AX instr_data_3__i23 (.D(instr_data[6]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i23.GSR = "DISABLED";
    FD1P3AX instr_data_3__i22 (.D(instr_data[5]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i22.GSR = "DISABLED";
    FD1P3AX instr_data_3__i21 (.D(instr_data[4]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i21.GSR = "DISABLED";
    FD1P3AX instr_data_3__i20 (.D(instr_data[3]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i20.GSR = "DISABLED";
    FD1P3AX instr_data_3__i19 (.D(instr_data[2]), .SP(clk_c_enable_292), 
            .CK(clk_c), .Q(n36[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i19.GSR = "DISABLED";
    FD1P3AX instr_data_3__i18 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_294), 
            .CK(clk_c), .Q(n36[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i18.GSR = "DISABLED";
    FD1P3AX instr_data_3__i17 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_294), 
            .CK(clk_c), .Q(\instr_data[2][0] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i17.GSR = "DISABLED";
    FD1P3AX instr_data_3__i16 (.D(instr_data[15]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i16.GSR = "DISABLED";
    FD1P3AX instr_data_3__i15 (.D(instr_data[14]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i15.GSR = "DISABLED";
    FD1P3AX instr_data_3__i14 (.D(instr_data[13]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i14.GSR = "DISABLED";
    FD1P3AX instr_data_3__i13 (.D(instr_data[12]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i13.GSR = "DISABLED";
    FD1P3AX instr_data_3__i12 (.D(instr_data[11]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i12.GSR = "DISABLED";
    FD1P3AX instr_data_3__i11 (.D(instr_data[10]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i11.GSR = "DISABLED";
    FD1P3AX instr_data_3__i10 (.D(instr_data[9]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i10.GSR = "DISABLED";
    FD1P3AX instr_data_3__i9 (.D(instr_data[8]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i9.GSR = "DISABLED";
    FD1P3AX instr_data_3__i8 (.D(instr_data[7]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(\instr_data[3][7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i8.GSR = "DISABLED";
    FD1P3AX instr_data_3__i7 (.D(instr_data[6]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i7.GSR = "DISABLED";
    FD1P3AX instr_data_3__i6 (.D(instr_data[5]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i6.GSR = "DISABLED";
    FD1P3AX instr_data_3__i5 (.D(instr_data[4]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i5.GSR = "DISABLED";
    FD1P3AX instr_data_3__i4 (.D(instr_data[3]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i4.GSR = "DISABLED";
    FD1P3AX instr_data_3__i3 (.D(instr_data[2]), .SP(clk_c_enable_308), 
            .CK(clk_c), .Q(n31[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i3.GSR = "DISABLED";
    FD1P3AX instr_data_3__i2 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_309), 
            .CK(clk_c), .Q(n31[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i2.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_781 (.A(\instr_addr_23__N_318[0] ), .B(instr_addr_23__N_318[1]), 
         .Z(n32796)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_rep_781.init = 16'hbbbb;
    PFUMX i29037 (.BLUT(n32051), .ALUT(n32050), .C0(n32539), .Z(n32052));
    LUT4 i1_2_lut_rep_782 (.A(\instr_addr_23__N_318[0] ), .B(instr_addr_23__N_318[1]), 
         .Z(n32797)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_782.init = 16'hdddd;
    LUT4 i1_2_lut_rep_783 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .Z(n32798)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_783.init = 16'heeee;
    FD1P3IX is_auipc_395 (.D(is_auipc_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_auipc)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_auipc_395.GSR = "DISABLED";
    LUT4 mux_2111_i28_3_lut_3_lut (.A(n32525), .B(n3493[17]), .C(n2131[11]), 
         .Z(n3446[27])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2111_i28_3_lut_3_lut.init = 16'he4e4;
    PFUMX i29027 (.BLUT(n32032), .ALUT(n32030), .C0(n32540), .Z(n32033));
    FD1P3AX data_ready_latch_416 (.D(n27854), .SP(clk_c_enable_325), .CK(clk_c), 
            .Q(data_ready_latch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(235[12] 256[8])
    defparam data_ready_latch_416.GSR = "DISABLED";
    LUT4 i27905_3_lut_3_lut (.A(\imm[10] ), .B(n9620), .C(n5605[2]), .Z(n5640[2])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i27905_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_3_lut_rep_526_4_lut (.A(n32545), .B(n32552), .C(n10024), .D(n32546), 
         .Z(n32541)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i1_3_lut_rep_526_4_lut.init = 16'h000e;
    LUT4 i14893_2_lut_rep_786 (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .Z(n32801)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14893_2_lut_rep_786.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n32639), .B(n27), .C(n32653), .D(n32654), 
         .Z(n29025)) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'hf444;
    LUT4 i15639_2_lut_rep_680_3_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(n8109), .Z(n32695)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i15639_2_lut_rep_680_3_lut.init = 16'h8f8f;
    LUT4 is_alu_imm_N_1367_bdd_3_lut_29150_4_lut_4_lut (.A(n32639), .B(n32655), 
         .C(n32582), .D(n32643), .Z(n32267)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam is_alu_imm_N_1367_bdd_3_lut_29150_4_lut_4_lut.init = 16'h0400;
    LUT4 i15576_2_lut_rep_713_3_lut_4_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(n32850), .D(addr[27]), .Z(n32728)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(C+(D))) */ ;
    defparam i15576_2_lut_rep_713_3_lut_4_lut.init = 16'h888f;
    LUT4 i1_3_lut_4_lut_adj_418 (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(addr[2]), .D(is_timer_addr), .Z(timer_data_3__N_631)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_418.init = 16'h7000;
    LUT4 i1_2_lut_3_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(data_ready_sync), .Z(n29173)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i15659_2_lut_rep_697_3_lut_4_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(n32850), .D(addr[27]), .Z(n32712)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i15659_2_lut_rep_697_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_4_lut_4_lut_adj_419 (.A(n32639), .B(n32612), .C(n32633), .D(n32576), 
         .Z(is_lui_N_1365)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_419.init = 16'h4000;
    FD1P3IX alu_op__i3 (.D(alu_op_de[3]), .SP(clk_c_enable_338), .CD(n32840), 
            .CK(clk_c), .Q(alu_op[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i3.GSR = "DISABLED";
    FD1P3IX alu_op__i2 (.D(alu_op_de[2]), .SP(clk_c_enable_338), .CD(n32840), 
            .CK(clk_c), .Q(alu_op_in[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i2.GSR = "DISABLED";
    FD1P3IX alu_op__i1 (.D(alu_op_de[1]), .SP(clk_c_enable_338), .CD(n32840), 
            .CK(clk_c), .Q(alu_op[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i1.GSR = "DISABLED";
    LUT4 i24568_2_lut_rep_730_3_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(addr[2]), .Z(n32745)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i24568_2_lut_rep_730_3_lut.init = 16'hf8f8;
    LUT4 i14936_2_lut_3_lut_3_lut (.A(n32639), .B(n32655), .C(n32656), 
         .Z(n22_adj_3179)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;
    defparam i14936_2_lut_3_lut_3_lut.init = 16'h5454;
    PFUMX i29022 (.BLUT(n32027), .ALUT(n32024), .C0(n32540), .Z(n32028));
    LUT4 i1_3_lut_4_lut_adj_420 (.A(n32563), .B(n9_adj_3180), .C(n28501), 
         .D(n10024), .Z(n28505)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_adj_420.init = 16'h0070;
    LUT4 i1_2_lut_rep_649_3_lut_4_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(is_timer_addr), .D(addr[2]), .Z(n32664)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_2_lut_rep_649_3_lut_4_lut.init = 16'h0070;
    FD1P3IX is_jal_401 (.D(is_jal_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_jal)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_jal_401.GSR = "DISABLED";
    LUT4 mux_40_i1_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[28]), 
         .D(data_rs2[0]), .Z(n92[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_40_i2_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[29]), 
         .D(data_rs2[1]), .Z(n92[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2111_i31_3_lut_3_lut (.A(n32525), .B(n3493[17]), .C(n29733), 
         .Z(n3446[30])) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2111_i31_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_2135_i30_3_lut_4_lut (.A(n32525), .B(n32540), .C(n3446[24]), 
         .D(n5205[29]), .Z(n3534[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2135_i30_3_lut_4_lut.init = 16'hf870;
    LUT4 i38_4_lut_3_lut_rep_596 (.A(n32654), .B(n24), .C(n32653), .Z(n32611)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i38_4_lut_3_lut_rep_596.init = 16'ha4a4;
    LUT4 mux_40_i3_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[30]), 
         .D(data_rs2[2]), .Z(n92[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_40_i4_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[31]), 
         .D(data_rs2[3]), .Z(n92[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i28441_2_lut_3_lut (.A(n32654), .B(n32653), .C(n32340), .Z(mem_op_de[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A (C))) */ ;
    defparam i28441_2_lut_3_lut.init = 16'h0d0d;
    FD1P3AX rs2_i0_i0 (.D(n2302[0]), .SP(clk_c_enable_524), .CK(clk_c), 
            .Q(rs2[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_3_lut (.A(n32654), .B(n32653), .C(n32639), .Z(n20_adj_3181)) /* synthesis lut_function=(A (B+(C))+!A !(B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'hb9b9;
    LUT4 i46_3_lut_3_lut (.A(n32656), .B(n32655), .C(n32639), .Z(n41)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;
    defparam i46_3_lut_3_lut.init = 16'h4a4a;
    LUT4 i1_3_lut_3_lut_4_lut (.A(n32656), .B(n32655), .C(n32653), .D(n32639), 
         .Z(n27896)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_3_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 mux_1549_i2_rep_134_3_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .Z(n30920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i2_rep_134_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_421 (.A(n32656), .B(n32655), .C(n32653), 
         .D(n32654), .Z(is_jal_N_1374)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_421.init = 16'h0400;
    LUT4 mux_2135_i25_3_lut_4_lut (.A(n32525), .B(n32540), .C(n3446[24]), 
         .D(n5205[24]), .Z(n3534[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2135_i25_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_2135_i26_3_lut_4_lut (.A(n32525), .B(n32540), .C(n3446[24]), 
         .D(n5205[25]), .Z(n3534[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2135_i26_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_345_i1_3_lut (.A(\next_pc_for_core[3] ), .B(return_addr[3]), 
         .C(n32544), .Z(n1742_adj_3219[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i1_3_lut.init = 16'hcaca;
    LUT4 i16_4_lut (.A(n28249), .B(clk_c_enable_41), .C(rst_reg_n_adj_6), 
         .D(n32525), .Z(clk_c_enable_383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i16_4_lut.init = 16'hcfca;
    LUT4 i1_4_lut_4_lut_4_lut_adj_422 (.A(n32641), .B(n32637), .C(n328[1]), 
         .D(n32581), .Z(n27788)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_4_lut_4_lut_4_lut_adj_422.init = 16'h00c4;
    LUT4 i1_2_lut_3_lut_adj_423 (.A(n32641), .B(n34287), .C(n32656), .Z(n28269)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i1_2_lut_3_lut_adj_423.init = 16'h8080;
    LUT4 mux_1562_i1_4_lut (.A(n32658), .B(rs2[0]), .C(n32548), .D(mem_op_increment_reg), 
         .Z(n2281[0])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1562_i1_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_3_lut_adj_424 (.A(n32641), .B(rst_reg_n_adj_6), .C(n13140), 
         .Z(n27430)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i1_2_lut_3_lut_adj_424.init = 16'h8080;
    LUT4 i1_4_lut_adj_425 (.A(n4271), .B(n32543), .C(n32546), .D(n28715), 
         .Z(n28249)) /* synthesis lut_function=(A+!((C+!(D))+!B)) */ ;
    defparam i1_4_lut_adj_425.init = 16'haeaa;
    FD1P3IX is_lui_398 (.D(is_lui_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_lui)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_lui_398.GSR = "DISABLED";
    LUT4 mux_345_i2_3_lut (.A(\next_pc_for_core[4] ), .B(return_addr[4]), 
         .C(n32544), .Z(n1742_adj_3219[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i2_3_lut.init = 16'hcaca;
    FD1P3IX is_alu_reg_397 (.D(is_alu_reg_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_alu_reg)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_alu_reg_397.GSR = "DISABLED";
    FD1P3IX is_store_396 (.D(is_store_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_store)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_store_396.GSR = "DISABLED";
    LUT4 mux_345_i3_3_lut (.A(\next_pc_for_core[5] ), .B(return_addr[5]), 
         .C(n32544), .Z(n1742_adj_3219[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i3_3_lut.init = 16'hcaca;
    FD1P3IX is_alu_imm_394 (.D(is_alu_imm_de), .SP(clk_c_enable_364), .CD(n32840), 
            .CK(clk_c), .Q(is_alu_imm)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_alu_imm_394.GSR = "DISABLED";
    FD1P3AX mem_op_increment_reg_413 (.D(mem_op_increment_reg_de), .SP(clk_c_enable_365), 
            .CK(clk_c), .Q(mem_op_increment_reg)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_increment_reg_413.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_426 (.A(n32617), .B(n32569), .C(rst_reg_n_adj_6), 
         .D(n32570), .Z(n28585)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_426.init = 16'h0080;
    LUT4 mux_345_i4_3_lut (.A(\next_pc_for_core[6] ), .B(return_addr[6]), 
         .C(n32544), .Z(n1742_adj_3219[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i4_3_lut.init = 16'hcaca;
    LUT4 mux_345_i5_3_lut (.A(\next_pc_for_core[7] ), .B(return_addr[7]), 
         .C(n32544), .Z(n1742_adj_3219[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i5_3_lut.init = 16'hcaca;
    PFUMX i29018 (.BLUT(n32020), .ALUT(n32017), .C0(n32540), .Z(n32021));
    LUT4 mux_345_i6_3_lut (.A(\next_pc_for_core[8] ), .B(return_addr[8]), 
         .C(n32544), .Z(n1742_adj_3219[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i6_3_lut.init = 16'hcaca;
    FD1P3AX instr_fetch_running_429 (.D(n6396), .SP(clk_c_enable_367), .CK(clk_c), 
            .Q(instr_fetch_running)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_fetch_running_429.GSR = "DISABLED";
    LUT4 mux_1539_i6_3_lut (.A(n33[5]), .B(n34[5]), .C(n2130), .Z(n2202[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1543_i6_3_lut (.A(n36[5]), .B(n31[5]), .C(n2150), .Z(n2222[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i6_3_lut.init = 16'hcaca;
    LUT4 mux_345_i7_3_lut (.A(\next_pc_for_core[9] ), .B(return_addr[9]), 
         .C(n32544), .Z(n1742_adj_3219[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i7_3_lut.init = 16'hcaca;
    LUT4 mux_345_i8_3_lut (.A(\next_pc_for_core[10] ), .B(return_addr[10]), 
         .C(n32544), .Z(n1742_adj_3219[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1539_i3_3_lut (.A(n33[2]), .B(n34[2]), .C(n2130), .Z(n2202[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i3_3_lut.init = 16'hcaca;
    LUT4 mux_345_i9_3_lut (.A(\next_pc_for_core[11] ), .B(return_addr[11]), 
         .C(n32544), .Z(n1742_adj_3219[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i9_3_lut.init = 16'hcaca;
    LUT4 mux_345_i10_3_lut (.A(\next_pc_for_core[12] ), .B(return_addr[12]), 
         .C(n32544), .Z(n1742_adj_3219[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1543_i3_3_lut (.A(n36[2]), .B(n31[2]), .C(n2150), .Z(n2222[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i3_3_lut.init = 16'hcaca;
    LUT4 i19156_4_lut (.A(n32704), .B(data_rs1[0]), .C(n32702), .D(mip_reg[16]), 
         .Z(n21667)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(78[10:20])
    defparam i19156_4_lut.init = 16'hf2c0;
    LUT4 mux_345_i11_3_lut (.A(\next_pc_for_core[13] ), .B(return_addr[13]), 
         .C(n32544), .Z(n1742_adj_3219[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i11_3_lut.init = 16'hcaca;
    LUT4 c_2__N_1861_1__bdd_4_lut_4_lut (.A(n34283), .B(counter_hi[2]), 
         .C(\pc[21] ), .D(\pc[17] ), .Z(n31649)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam c_2__N_1861_1__bdd_4_lut_4_lut.init = 16'h5140;
    LUT4 mux_345_i12_3_lut (.A(\next_pc_for_core[14] ), .B(return_addr[14]), 
         .C(n32544), .Z(n1742_adj_3219[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i12_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_427 (.A(n32543), .B(n32546), .C(n32548), .D(n28391), 
         .Z(n13140)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_427.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_428 (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[20] ), 
         .D(\next_pc_for_core[16] ), .Z(n225)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i1_4_lut_4_lut_adj_428.init = 16'h5140;
    LUT4 c_2__N_1861_1__bdd_4_lut_28780_4_lut (.A(n34283), .B(counter_hi[2]), 
         .C(\pc[23] ), .D(\pc[19] ), .Z(n31619)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam c_2__N_1861_1__bdd_4_lut_28780_4_lut.init = 16'h5140;
    LUT4 mux_1539_i4_3_lut (.A(n33[3]), .B(n34[3]), .C(n2130), .Z(n2202[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i4_3_lut.init = 16'hcaca;
    LUT4 c_2__N_1861_1__bdd_4_lut_28800_4_lut (.A(n34283), .B(counter_hi[2]), 
         .C(\pc[22] ), .D(\pc[18] ), .Z(n31624)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam c_2__N_1861_1__bdd_4_lut_28800_4_lut.init = 16'h5140;
    LUT4 i15141_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\pc[20] ), 
         .D(\pc[16] ), .Z(n225_adj_3185)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i15141_4_lut_4_lut.init = 16'h5140;
    FD1P3AX imm_i0_i31 (.D(n3446[24]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm_c[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i31.GSR = "DISABLED";
    LUT4 mux_1543_i4_3_lut (.A(n36[3]), .B(n31[3]), .C(n2150), .Z(n2222[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i4_3_lut.init = 16'hcaca;
    LUT4 mux_345_i13_3_lut (.A(\next_pc_for_core[15] ), .B(return_addr[15]), 
         .C(n32544), .Z(n1742_adj_3219[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i13_3_lut.init = 16'hcaca;
    LUT4 i15171_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[21] ), 
         .D(\next_pc_for_core[17] ), .Z(n226)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i15171_4_lut_4_lut.init = 16'h5140;
    FD1P3AX imm_i0_i30 (.D(n3534[30]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm_c[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i30.GSR = "DISABLED";
    FD1P3AX imm_i0_i29 (.D(n3534[29]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm_c[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i29.GSR = "DISABLED";
    FD1P3AX imm_i0_i28 (.D(n3534[28]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm_c[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i28.GSR = "DISABLED";
    FD1P3AX imm_i0_i27 (.D(n3534[27]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm_c[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i27.GSR = "DISABLED";
    FD1P3AX imm_i0_i26 (.D(n3534[26]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm_c[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i26.GSR = "DISABLED";
    FD1P3AX imm_i0_i25 (.D(n3534[25]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm_c[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i25.GSR = "DISABLED";
    FD1P3AX imm_i0_i24 (.D(n3534[24]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(imm_c[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i24.GSR = "DISABLED";
    FD1P3AX imm_i0_i23 (.D(n3534[23]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i23.GSR = "DISABLED";
    FD1P3AX imm_i0_i22 (.D(n3534[22]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i22.GSR = "DISABLED";
    FD1P3AX imm_i0_i21 (.D(n3534[21]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i21.GSR = "DISABLED";
    FD1P3AX imm_i0_i20 (.D(n3534[20]), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i20.GSR = "DISABLED";
    FD1P3AX imm_i0_i19 (.D(n32034), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i19.GSR = "DISABLED";
    FD1P3AX imm_i0_i18 (.D(n32029), .SP(clk_c_enable_383), .CK(clk_c), 
            .Q(\imm[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i18.GSR = "DISABLED";
    LUT4 i15172_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[22] ), 
         .D(\next_pc_for_core[18] ), .Z(n227)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i15172_4_lut_4_lut.init = 16'h5140;
    LUT4 mux_345_i15_3_lut (.A(\next_pc_for_core[17] ), .B(return_addr[17]), 
         .C(n32544), .Z(n1742_adj_3219[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i15_3_lut.init = 16'hcaca;
    LUT4 mux_345_i16_3_lut (.A(\next_pc_for_core[18] ), .B(return_addr[18]), 
         .C(n32544), .Z(n1742_adj_3219[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i16_3_lut.init = 16'hcaca;
    LUT4 i27350_2_lut_rep_793 (.A(n34281), .B(n34283), .Z(n32808)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i27350_2_lut_rep_793.init = 16'h4444;
    LUT4 pc_23__I_0_450_i269_rep_70_3_lut_4_lut (.A(counter_hi[4]), .B(counter_hi[3]), 
         .C(n209_adj_3186), .D(n157_adj_3187), .Z(n29689)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam pc_23__I_0_450_i269_rep_70_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_345_i17_3_lut (.A(\next_pc_for_core[19] ), .B(return_addr[19]), 
         .C(n32544), .Z(n1742_adj_3219[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i17_3_lut.init = 16'hcaca;
    LUT4 mux_345_i18_3_lut (.A(\next_pc_for_core[20] ), .B(return_addr[20]), 
         .C(n32544), .Z(n1742_adj_3219[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i18_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_3_lut_adj_429 (.A(addr[6]), .B(n15_adj_3188), .C(n32754), 
         .Z(n28077)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_3_lut_3_lut_adj_429.init = 16'h4040;
    LUT4 mux_345_i19_3_lut (.A(\next_pc_for_core[21] ), .B(return_addr[21]), 
         .C(n32544), .Z(n1742_adj_3219[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i19_3_lut.init = 16'hcaca;
    LUT4 mux_2135_i29_3_lut_4_lut (.A(n32525), .B(n32540), .C(n3446[24]), 
         .D(n5205[28]), .Z(n3534[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2135_i29_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_345_i20_3_lut (.A(\next_pc_for_core[22] ), .B(return_addr[22]), 
         .C(n32544), .Z(n1742_adj_3219[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i20_3_lut.init = 16'hcaca;
    LUT4 mux_345_i21_3_lut (.A(\next_pc_for_core[23] ), .B(return_addr[23]), 
         .C(n32544), .Z(n1742_adj_3219[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i21_3_lut.init = 16'hcaca;
    LUT4 i15485_4_lut (.A(n2131[11]), .B(n32563), .C(n2151[11]), .D(n32734), 
         .Z(n5205[7])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15485_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_430 (.A(n32548), .B(n35), .C(n28575), .D(n32611), 
         .Z(n28715)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_430.init = 16'h5040;
    LUT4 mux_1562_i2_4_lut (.A(n32657), .B(rs2[1]), .C(n32548), .D(n32853), 
         .Z(n2281[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1562_i2_4_lut.init = 16'h3aca;
    LUT4 i21711_1_lut_rep_797 (.A(counter_hi[2]), .Z(n32812)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i21711_1_lut_rep_797.init = 16'h5555;
    LUT4 i1_4_lut_4_lut_adj_431 (.A(counter_hi[2]), .B(clk_c_enable_538), 
         .C(n32677), .D(n32760), .Z(clk_c_enable_321)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i1_4_lut_4_lut_adj_431.init = 16'h0100;
    LUT4 mux_1562_i3_4_lut (.A(n32661), .B(rs2[2]), .C(n32548), .D(n32773), 
         .Z(n2281[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1562_i3_4_lut.init = 16'h3aca;
    LUT4 mux_1549_i12_3_lut_rep_622 (.A(n2202[11]), .B(n2222[11]), .C(n32734), 
         .Z(n32637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i12_3_lut_rep_622.init = 16'hcaca;
    LUT4 i15018_2_lut_4_lut (.A(n2202[11]), .B(n2222[11]), .C(n32734), 
         .D(n32656), .Z(n17665)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15018_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_1539_i15_3_lut (.A(n33[14]), .B(n34[14]), .C(n2130), .Z(n2202[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1562_i4_4_lut (.A(n32659), .B(rs2[3]), .C(n32548), .D(n6634), 
         .Z(n2281[3])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1562_i4_4_lut.init = 16'h3aca;
    LUT4 i1_2_lut_rep_590_4_lut (.A(n2202[11]), .B(n2222[11]), .C(n32734), 
         .D(n32641), .Z(n32605)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_590_4_lut.init = 16'hca00;
    LUT4 i15355_2_lut_2_lut_4_lut (.A(n2202[11]), .B(n2222[11]), .C(n32734), 
         .D(n32656), .Z(n5138[3])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15355_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_1543_i15_3_lut (.A(n36[14]), .B(n31[14]), .C(n2150), .Z(n2222[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1539_i14_3_lut (.A(n33[13]), .B(n34[13]), .C(n2130), .Z(n2202[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1543_i14_3_lut (.A(n36[13]), .B(n31[13]), .C(n2150), .Z(n2222[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1549_i16_3_lut_rep_624 (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .Z(n32639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i16_3_lut_rep_624.init = 16'hcaca;
    LUT4 i1_2_lut_rep_582_2_lut_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32655), .Z(n32597)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_582_2_lut_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_rep_614_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32654), .Z(n32629)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_614_4_lut.init = 16'hca00;
    LUT4 i28257_2_lut_rep_613_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32654), .Z(n32628)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i28257_2_lut_rep_613_4_lut.init = 16'h0035;
    LUT4 i15346_2_lut_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32651), .Z(n2970[4])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15346_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_2_lut_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32654), .Z(n12_adj_3192)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_2_lut_4_lut.init = 16'h3500;
    L6MUX21 i27548 (.D0(n30255), .D1(n30256), .SD(counter_hi[4]), .Z(debug_rd_3__N_405[30]));
    L6MUX21 i27555 (.D0(n30262), .D1(n30263), .SD(n34281), .Z(debug_rd_3__N_405[31]));
    LUT4 i10453_3_lut (.A(n13156), .B(n32053), .C(n32525), .Z(n3534[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i10453_3_lut.init = 16'hcaca;
    LUT4 i14875_2_lut_rep_598_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32656), .Z(n32613)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i14875_2_lut_rep_598_4_lut.init = 16'hffca;
    LUT4 i1_3_lut_adj_432 (.A(n32640), .B(n13140), .C(rst_reg_n_adj_6), 
         .Z(n27428)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i1_3_lut_adj_432.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_433 (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n34287), .Z(n28407)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_433.init = 16'hca00;
    LUT4 i1_2_lut_4_lut_adj_434 (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32654), .Z(n29211)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_434.init = 16'h00ca;
    LUT4 i1_2_lut_rep_804 (.A(addr[2]), .B(addr[3]), .Z(n32819)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_804.init = 16'heeee;
    LUT4 i6610_4_lut (.A(n29727), .B(instr[26]), .C(n32540), .D(n32563), 
         .Z(n3328[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i6610_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_rep_612_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32655), .Z(n32627)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_612_4_lut.init = 16'hffca;
    LUT4 i15349_2_lut_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32657), .Z(n2970[7])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15349_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_rep_705_3_lut_4_lut (.A(addr[2]), .B(addr[3]), .C(n32835), 
         .D(n32836), .Z(n32720)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_705_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_435 (.A(addr[2]), .B(addr[3]), .C(\addr[5] ), 
         .Z(n29357)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_435.init = 16'h1010;
    LUT4 i1_2_lut_rep_604_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32656), .Z(n32619)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_604_4_lut.init = 16'hca00;
    LUT4 i1_2_lut_rep_601_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32655), .Z(n32616)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_601_4_lut.init = 16'h00ca;
    LUT4 i1_4_lut_4_lut_adj_436 (.A(addr[7]), .B(n32720), .C(n19_adj_3193), 
         .D(\uo_out_from_user_peri[1][6] ), .Z(n20)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_4_lut_4_lut_adj_436.init = 16'h5140;
    LUT4 i28578_2_lut_4_lut (.A(n2202[15]), .B(n2222[15]), .C(n32734), 
         .D(n32653), .Z(n30132)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i28578_2_lut_4_lut.init = 16'hff35;
    LUT4 i1_4_lut_4_lut_adj_437 (.A(addr[7]), .B(n32720), .C(\data_from_user_peri_1__31__N_2455[2] ), 
         .D(\uo_out_from_user_peri[1][2] ), .Z(n5)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_4_lut_4_lut_adj_437.init = 16'h5140;
    LUT4 mux_1549_i10_3_lut_rep_625 (.A(n2202[9]), .B(n2222[9]), .C(n32734), 
         .Z(n32640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i10_3_lut_rep_625.init = 16'hcaca;
    LUT4 i1_4_lut_adj_438 (.A(n10024), .B(n32617), .C(n32566), .D(n34287), 
         .Z(n28731)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_438.init = 16'h1000;
    LUT4 i1_4_lut_4_lut_adj_439 (.A(addr[7]), .B(n32720), .C(data_from_user_peri_1__31__N_2455[5]), 
         .D(\uo_out_from_user_peri[1][5] ), .Z(n21)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_4_lut_4_lut_adj_439.init = 16'h5140;
    LUT4 i1_4_lut_4_lut_adj_440 (.A(addr[7]), .B(n32851), .C(n29485), 
         .D(n32771), .Z(n29491)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_4_lut_4_lut_adj_440.init = 16'hf7ff;
    LUT4 i14957_2_lut_2_lut_4_lut (.A(n2202[9]), .B(n2222[9]), .C(n32734), 
         .D(n32538), .Z(n1708[2])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i14957_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 i26955_3_lut (.A(n32641), .B(n13140), .C(n4243), .Z(n29594)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(47[17:22])
    defparam i26955_3_lut.init = 16'hecec;
    LUT4 mux_1539_i2_3_lut (.A(n33[1]), .B(n34[1]), .C(n2130), .Z(n2202[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i2_3_lut.init = 16'hcaca;
    LUT4 i15343_2_lut_4_lut (.A(n2202[9]), .B(n2222[9]), .C(n32734), .D(n32656), 
         .Z(n2590[2])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15343_2_lut_4_lut.init = 16'h00ca;
    LUT4 i14975_2_lut_2_lut_4_lut (.A(n2202[9]), .B(n2222[9]), .C(n32734), 
         .D(n32653), .Z(n1713[2])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i14975_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_1549_i11_3_lut_rep_626 (.A(n2202[10]), .B(n2222[10]), .C(n32734), 
         .Z(n32641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i11_3_lut_rep_626.init = 16'hcaca;
    PFUMX i29385 (.BLUT(n32992), .ALUT(\data_from_read[2] ), .C0(n32771), 
          .Z(n32993));
    LUT4 mux_1543_i2_3_lut (.A(n36[1]), .B(n31[1]), .C(n2150), .Z(n2222[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i2_3_lut.init = 16'hcaca;
    LUT4 i14974_2_lut_2_lut_4_lut (.A(n2202[10]), .B(n2222[10]), .C(n32734), 
         .D(n32653), .Z(n1713[3])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i14974_2_lut_2_lut_4_lut.init = 16'hcaff;
    LUT4 i14956_2_lut_2_lut_4_lut (.A(n2202[10]), .B(n2222[10]), .C(n32734), 
         .D(n32538), .Z(n1708[3])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i14956_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 n14_bdd_2_lut_29192_4_lut (.A(n2202[10]), .B(n2222[10]), .C(n32734), 
         .D(n32651), .Z(n31589)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam n14_bdd_2_lut_29192_4_lut.init = 16'h3500;
    LUT4 i1_4_lut_adj_441 (.A(n29163), .B(n27888), .C(n29165), .D(n29161), 
         .Z(is_timer_addr)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_441.init = 16'h8000;
    LUT4 i1_4_lut_adj_442 (.A(\addr[23] ), .B(n29155), .C(n29145), .D(\addr[20] ), 
         .Z(n29163)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_442.init = 16'h8000;
    LUT4 is_branch_I_0_475_2_lut_rep_806 (.A(is_branch), .B(n34285), .Z(n32821)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam is_branch_I_0_475_2_lut_rep_806.init = 16'h8888;
    LUT4 mux_832_i5_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[7] ), 
         .D(addr_out[7]), .Z(n1203[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_443 (.A(n29159), .B(addr_c[26]), .C(n29141), .D(addr_c[25]), 
         .Z(n29165)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_443.init = 16'h8000;
    LUT4 i1_4_lut_adj_444 (.A(addr[10]), .B(\addr[8] ), .C(\addr[24] ), 
         .D(\addr[16] ), .Z(n29161)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_444.init = 16'h8000;
    LUT4 i15344_2_lut_4_lut (.A(n2202[10]), .B(n2222[10]), .C(n32734), 
         .D(n32656), .Z(n2590[3])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15344_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_1549_i13_3_lut_rep_627 (.A(n2202[12]), .B(n2222[12]), .C(n32734), 
         .Z(n32642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i13_3_lut_rep_627.init = 16'hcaca;
    LUT4 i1_4_lut_adj_445 (.A(\addr[12] ), .B(\addr[21] ), .C(\addr[13] ), 
         .D(\addr[15] ), .Z(n29155)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_445.init = 16'h8000;
    LUT4 mux_832_i1_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[3] ), 
         .D(addr_out[3]), .Z(n1203[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_446 (.A(n2202[12]), .B(n2222[12]), .C(n32734), 
         .D(n32655), .Z(n29039)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_446.init = 16'hca00;
    LUT4 equal_25_i3_2_lut_4_lut (.A(n2202[12]), .B(n2222[12]), .C(n32734), 
         .D(n32655), .Z(n3_adj_3194)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam equal_25_i3_2_lut_4_lut.init = 16'hff35;
    LUT4 mux_832_i4_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[6] ), 
         .D(addr_out[6]), .Z(n1203[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3069_i2_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[2] ), .D(n32690), .Z(n5017[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_3069_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i2_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[4] ), 
         .D(addr_out[4]), .Z(n1203[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1549_i9_3_lut_rep_628 (.A(n2202[8]), .B(n2222[8]), .C(n32734), 
         .Z(n32643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i9_3_lut_rep_628.init = 16'hcaca;
    LUT4 i14958_2_lut_2_lut_4_lut (.A(n2202[8]), .B(n2222[8]), .C(n32734), 
         .D(n32538), .Z(n1708[1])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i14958_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 i14976_2_lut_2_lut_4_lut (.A(n2202[8]), .B(n2222[8]), .C(n32734), 
         .D(n32653), .Z(n1713[1])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i14976_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_3069_i1_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(n32822), .D(addr_out[1]), .Z(n5017[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_3069_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i6_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[8] ), 
         .D(addr_out[8]), .Z(n1203[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i3_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[5] ), 
         .D(addr_out[5]), .Z(n1203[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_447 (.A(\addr[22] ), .B(\addr[14] ), .Z(n29145)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_447.init = 16'h8888;
    LUT4 i27552_3_lut (.A(imm_c[27]), .B(imm_c[31]), .C(counter_hi[2]), 
         .Z(n30261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27552_3_lut.init = 16'hcaca;
    LUT4 i15351_2_lut_4_lut (.A(n2202[8]), .B(n2222[8]), .C(n32734), .D(n2792), 
         .Z(n2585[1])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15351_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_4_lut_adj_448 (.A(\addr[9] ), .B(\addr[17] ), .C(addr[27]), 
         .D(\addr[11] ), .Z(n29159)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_448.init = 16'h8000;
    LUT4 i27551_3_lut (.A(\imm[19] ), .B(\imm[23] ), .C(counter_hi[2]), 
         .Z(n30260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27551_3_lut.init = 16'hcaca;
    LUT4 mux_832_i7_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[9] ), 
         .D(addr_out[9]), .Z(n1203[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_449 (.A(\addr[19] ), .B(\addr[18] ), .Z(n29141)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_449.init = 16'h8888;
    LUT4 mux_832_i8_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[10] ), 
         .D(addr_out[10]), .Z(n1203[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i9_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[11] ), 
         .D(addr_out[11]), .Z(n1203[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i28203_3_lut (.A(n3328[12]), .B(n5205[12]), .C(n32540), .Z(n3446[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28203_3_lut.init = 16'hcaca;
    LUT4 mux_832_i10_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[12] ), .D(addr_out[12]), .Z(n1203[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i28201_3_lut (.A(n3328[13]), .B(n5205[13]), .C(n32540), .Z(n3446[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28201_3_lut.init = 16'hcaca;
    LUT4 i28199_3_lut (.A(n3328[14]), .B(n5205[14]), .C(n32540), .Z(n3446[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28199_3_lut.init = 16'hcaca;
    LUT4 mux_832_i11_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[13] ), .D(addr_out[13]), .Z(n1203[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i12_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[14] ), .D(addr_out[14]), .Z(n1203[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i13_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[15] ), .D(addr_out[15]), .Z(n1203[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i15_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[17] ), .D(addr_out[17]), .Z(n1203[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i16_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[18] ), .D(addr_out[18]), .Z(n1203[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i17_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[19] ), .D(addr_out[19]), .Z(n1203[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i18_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[20] ), .D(addr_out[20]), .Z(n1203[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_rep_549 (.A(is_timer_addr), .B(n32575), .C(data_ready_latch), 
         .Z(n32564)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(258[53:106])
    defparam i1_3_lut_rep_549.init = 16'hfefe;
    LUT4 i5568_2_lut_4_lut (.A(is_timer_addr), .B(n32575), .C(data_ready_latch), 
         .D(n32829), .Z(n8228)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(258[53:106])
    defparam i5568_2_lut_4_lut.init = 16'hfe00;
    LUT4 i28165_3_lut_4_lut (.A(n32658), .B(n32565), .C(n2557), .D(n27516), 
         .Z(n2291[0])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28165_3_lut_4_lut.init = 16'hefe0;
    LUT4 i28161_3_lut_4_lut_4_lut (.A(n32565), .B(n27523), .C(n2557), 
         .D(n32661), .Z(n2291[2])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam i28161_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i28197_3_lut (.A(n3328[15]), .B(n5205[15]), .C(n32540), .Z(n3446[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28197_3_lut.init = 16'hcaca;
    LUT4 mux_1539_i7_3_lut (.A(n33[6]), .B(n34[6]), .C(n2130), .Z(n2202[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1520_i14_3_lut (.A(n31[13]), .B(n33[13]), .C(n2150), .Z(n2151[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i14_3_lut.init = 16'hcaca;
    FD1S3IX counter_hi_3544__i3 (.D(n39[1]), .CK(clk_c), .CD(n32840), 
            .Q(counter_hi[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3544__i3.GSR = "DISABLED";
    FD1S3IX counter_hi_3544__i4 (.D(n39[2]), .CK(clk_c), .CD(n32840), 
            .Q(counter_hi[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3544__i4.GSR = "DISABLED";
    FD1S3IX addr_offset_3545__i3 (.D(n38[1]), .CK(clk_c), .CD(n32840), 
            .Q(addr_offset[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam addr_offset_3545__i3.GSR = "DISABLED";
    LUT4 mux_832_i19_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[21] ), .D(addr_out[21]), .Z(n1203[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i20_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[22] ), .D(addr_out[22]), .Z(n1203[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_832_i21_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[23] ), .D(addr_out[23]), .Z(n1203[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_832_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 i15373_4_lut (.A(n32641), .B(n32656), .C(n32659), .D(n32653), 
         .Z(n3292[3])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15373_4_lut.init = 16'hc088;
    LUT4 mux_1543_i7_3_lut (.A(n36[6]), .B(n31[6]), .C(n2150), .Z(n2222[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i7_3_lut.init = 16'hcaca;
    LUT4 i28214_3_lut (.A(n3259[3]), .B(n3292[3]), .C(n4267), .Z(n3410[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i28214_3_lut.init = 16'hcaca;
    LUT4 i14153_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[16] ), 
         .D(addr_out[16]), .Z(n16811)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam i14153_3_lut_4_lut.init = 16'hf780;
    LUT4 i15374_4_lut (.A(n32637), .B(n32656), .C(n32651), .D(n32653), 
         .Z(n3292[4])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15374_4_lut.init = 16'hc088;
    LUT4 i15375_4_lut (.A(n32658), .B(n32656), .C(n32642), .D(n32653), 
         .Z(n3292[5])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15375_4_lut.init = 16'hc088;
    LUT4 i27550_3_lut (.A(\imm[11] ), .B(imm[15]), .C(counter_hi[2]), 
         .Z(n30259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27550_3_lut.init = 16'hcaca;
    LUT4 i15376_4_lut (.A(n32659), .B(n32656), .C(n32658), .D(n32653), 
         .Z(n3292[6])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15376_4_lut.init = 16'hc088;
    LUT4 mux_2084_i7_4_lut (.A(n2594), .B(n32659), .C(n4259), .D(n32639), 
         .Z(n3259[6])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2084_i7_4_lut.init = 16'hfaca;
    LUT4 i1_2_lut_rep_809 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .Z(n32824)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_809.init = 16'h8888;
    LUT4 i15377_4_lut (.A(n32651), .B(n32656), .C(n32657), .D(n32653), 
         .Z(n3292[7])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15377_4_lut.init = 16'hc088;
    LUT4 i28163_3_lut_4_lut_4_lut (.A(n32565), .B(n27502), .C(n2557), 
         .D(n32657), .Z(n2291[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam i28163_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i1_2_lut_3_lut_adj_450 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .C(n34287), .Z(n28821)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_450.init = 16'h8080;
    LUT4 i28159_3_lut_4_lut_4_lut (.A(n32565), .B(n27509), .C(n2557), 
         .D(n32659), .Z(n2291[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam i28159_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 mux_2126_i9_4_lut (.A(n3369[8]), .B(instr[28]), .C(n32525), .D(n9394), 
         .Z(n3493[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2126_i9_4_lut.init = 16'hca0a;
    LUT4 mux_1549_i7_3_lut_rep_636 (.A(n2202[6]), .B(n2222[6]), .C(n32734), 
         .Z(n32651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i7_3_lut_rep_636.init = 16'hcaca;
    LUT4 i15118_2_lut_rep_589_4_lut (.A(n2202[6]), .B(n2222[6]), .C(n32734), 
         .D(n32659), .Z(n32604)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15118_2_lut_rep_589_4_lut.init = 16'hca00;
    LUT4 mux_1516_i14_3_lut (.A(n34[13]), .B(n36[13]), .C(n2130), .Z(n2131[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i14_3_lut.init = 16'hcaca;
    LUT4 instr_6__I_0_128_i7_2_lut_rep_594_4_lut (.A(n2202[6]), .B(n2222[6]), 
         .C(n32734), .D(n32659), .Z(n32609)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_6__I_0_128_i7_2_lut_rep_594_4_lut.init = 16'hffca;
    LUT4 i27549_3_lut (.A(\imm[3] ), .B(\imm[7] ), .C(counter_hi[2]), 
         .Z(n30258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27549_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_813 (.A(debug_instr_valid), .B(no_write_in_progress), 
         .Z(n32828)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_2_lut_rep_813.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_451 (.A(debug_instr_valid), .B(no_write_in_progress), 
         .C(load_done), .D(is_load), .Z(instr_complete_N_1651)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_3_lut_4_lut_adj_451.init = 16'h8000;
    LUT4 instr_6__I_0_127_i7_2_lut_4_lut (.A(n2202[6]), .B(n2222[6]), .C(n32734), 
         .D(n32659), .Z(n7_adj_3196)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_6__I_0_127_i7_2_lut_4_lut.init = 16'hcaff;
    LUT4 i15357_2_lut_2_lut_4_lut (.A(n2202[6]), .B(n2222[6]), .C(n32734), 
         .D(n32656), .Z(n5138[6])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15357_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 i27545_3_lut (.A(imm_c[26]), .B(imm_c[30]), .C(counter_hi[2]), 
         .Z(n30254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27545_3_lut.init = 16'hcaca;
    LUT4 mux_1549_i2_3_lut_rep_638 (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .Z(n32653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i2_3_lut_rep_638.init = 16'hcaca;
    LUT4 i1_2_lut_rep_602_4_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .D(n32654), .Z(n32617)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_602_4_lut.init = 16'h00ca;
    LUT4 i24528_2_lut_rep_574_3_lut_2_lut_4_lut (.A(n2202[1]), .B(n2222[1]), 
         .C(n32734), .D(n32654), .Z(n32589)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i24528_2_lut_rep_574_3_lut_2_lut_4_lut.init = 16'h35ca;
    LUT4 i28495_2_lut_rep_593_4_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .D(n32656), .Z(n32608)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i28495_2_lut_rep_593_4_lut.init = 16'h3500;
    L6MUX21 i27751 (.D0(n30458), .D1(n30459), .SD(n34281), .Z(debug_rd_3__N_405[28]));
    L6MUX21 i27758 (.D0(n30465), .D1(n30466), .SD(n34281), .Z(debug_rd_3__N_405[29]));
    LUT4 i1_2_lut_2_lut_4_lut_adj_452 (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .D(n32269), .Z(n17_adj_3197)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_2_lut_4_lut_adj_452.init = 16'h3500;
    LUT4 i15031_2_lut_rep_615_4_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .D(n32654), .Z(n32630)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15031_2_lut_rep_615_4_lut.init = 16'hca00;
    LUT4 i166_2_lut_rep_608_4_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .D(n32654), .Z(n32623)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i166_2_lut_rep_608_4_lut.init = 16'h3500;
    L6MUX21 i28965 (.D0(n31882), .D1(n31879), .SD(\addr[4] ), .Z(n31883));
    LUT4 i15032_1_lut_rep_579_2_lut_4_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .D(n32654), .Z(n32594)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15032_1_lut_rep_579_2_lut_4_lut.init = 16'h35ff;
    LUT4 i27544_3_lut (.A(\imm[18] ), .B(\imm[22] ), .C(counter_hi[2]), 
         .Z(n30253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27544_3_lut.init = 16'hcaca;
    LUT4 n8539_bdd_1_lut_2_lut_4_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .D(additional_mem_ops_2__N_1132[0]), .Z(n32221)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam n8539_bdd_1_lut_2_lut_4_lut.init = 16'h35ff;
    LUT4 i1_2_lut_rep_618_4_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .D(n32654), .Z(n32633)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_618_4_lut.init = 16'h3500;
    LUT4 i15446_2_lut_rep_545_4_lut (.A(n2202[1]), .B(n2222[1]), .C(n32734), 
         .D(additional_mem_ops_2__N_1132[0]), .Z(n32560)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15446_2_lut_rep_545_4_lut.init = 16'hca00;
    LUT4 i27543_3_lut (.A(\imm[10] ), .B(imm[14]), .C(counter_hi[2]), 
         .Z(n30252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27543_3_lut.init = 16'hcaca;
    LUT4 mux_1549_i14_3_lut_rep_640 (.A(n2202[13]), .B(n2222[13]), .C(n32734), 
         .Z(n32655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i14_3_lut_rep_640.init = 16'hcaca;
    LUT4 i1_2_lut_rep_597_4_lut (.A(n2202[13]), .B(n2222[13]), .C(n32734), 
         .D(n32656), .Z(n32612)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_597_4_lut.init = 16'hca00;
    PFUMX i28960 (.BLUT(n31878), .ALUT(n29834), .C0(addr[2]), .Z(n31879));
    LUT4 i14940_2_lut_rep_617_4_lut (.A(n2202[13]), .B(n2222[13]), .C(n32734), 
         .D(n32656), .Z(n32632)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i14940_2_lut_rep_617_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_rep_587_4_lut (.A(n2202[13]), .B(n2222[13]), .C(n32734), 
         .D(n32656), .Z(n32602)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_587_4_lut.init = 16'hffca;
    LUT4 i27542_3_lut (.A(\imm[2] ), .B(\imm[6] ), .C(counter_hi[2]), 
         .Z(n30251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27542_3_lut.init = 16'hcaca;
    FD1P3IX pc_offset__i23 (.D(pc_23__N_911[20]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[23] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i23.GSR = "DISABLED";
    FD1P3IX pc_offset__i22 (.D(pc_23__N_911[19]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[22] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i22.GSR = "DISABLED";
    FD1P3IX pc_offset__i21 (.D(pc_23__N_911[18]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[21] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i21.GSR = "DISABLED";
    FD1P3IX pc_offset__i20 (.D(pc_23__N_911[17]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[20] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i20.GSR = "DISABLED";
    FD1P3IX pc_offset__i19 (.D(pc_23__N_911[16]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[19] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i19.GSR = "DISABLED";
    FD1P3IX pc_offset__i18 (.D(pc_23__N_911[15]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[18] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i18.GSR = "DISABLED";
    FD1P3IX pc_offset__i17 (.D(pc_23__N_911[14]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[17] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i17.GSR = "DISABLED";
    FD1P3IX pc_offset__i16 (.D(\pc_23__N_911[13] ), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[16] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i16.GSR = "DISABLED";
    FD1P3IX pc_offset__i15 (.D(pc_23__N_911[12]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[15] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i15.GSR = "DISABLED";
    FD1P3IX pc_offset__i14 (.D(pc_23__N_911[11]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[14] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i14.GSR = "DISABLED";
    LUT4 n14_bdd_2_lut_28756_2_lut_4_lut (.A(n2202[13]), .B(n2222[13]), 
         .C(n32734), .D(n32658), .Z(n31588)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam n14_bdd_2_lut_28756_2_lut_4_lut.init = 16'h3500;
    LUT4 mux_1549_i15_3_lut_rep_641 (.A(n2202[14]), .B(n2222[14]), .C(n32734), 
         .Z(n32656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i15_3_lut_rep_641.init = 16'hcaca;
    FD1P3IX pc_offset__i1 (.D(pc_2__N_932[0]), .SP(clk_c_enable_533), .CD(n32840), 
            .CK(clk_c), .Q(\pc[1] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i1.GSR = "DISABLED";
    FD1P3AX data_write_n_i1 (.D(data_write_n_1__N_369[1]), .SP(clk_c_enable_513), 
            .CK(clk_c), .Q(qv_data_write_n[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_write_n_i1.GSR = "DISABLED";
    FD1P3IX pc_offset__i13 (.D(pc_23__N_911[10]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[13] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i13.GSR = "DISABLED";
    LUT4 i15372_2_lut_4_lut (.A(n2202[14]), .B(n2222[14]), .C(n32734), 
         .D(n32661), .Z(n3292[2])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15372_2_lut_4_lut.init = 16'hca00;
    LUT4 additional_mem_ops_2__N_1132_0__bdd_2_lut_4_lut (.A(n2202[14]), .B(n2222[14]), 
         .C(n32734), .D(additional_mem_ops_2__N_1132[0]), .Z(n32427)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam additional_mem_ops_2__N_1132_0__bdd_2_lut_4_lut.init = 16'h00ca;
    FD1P3IX pc_offset__i12 (.D(pc_23__N_911[9]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[12] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i12.GSR = "DISABLED";
    FD1P3IX pc_offset__i11 (.D(pc_23__N_911[8]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[11] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i11.GSR = "DISABLED";
    FD1P3IX pc_offset__i10 (.D(pc_23__N_911[7]), .SP(clk_c_enable_533), 
            .CD(n32840), .CK(clk_c), .Q(\pc[10] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i10.GSR = "DISABLED";
    PFUMX i28963 (.BLUT(n31881), .ALUT(n31880), .C0(addr[3]), .Z(n31882));
    LUT4 i24_1_lut_rep_619_3_lut (.A(n2202[14]), .B(n2222[14]), .C(n32734), 
         .Z(n32634)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i24_1_lut_rep_619_3_lut.init = 16'h3535;
    LUT4 mux_2089_i5_3_lut (.A(n32637), .B(instr[24]), .C(n32533), .Z(n3328[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2089_i5_3_lut.init = 16'hcaca;
    LUT4 i28277_3_lut_4_lut (.A(n4251), .B(n32734), .C(n32539), .D(n32540), 
         .Z(n30014)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28277_3_lut_4_lut.init = 16'hff1f;
    LUT4 i41_2_lut_rep_820 (.A(\addr[1] ), .B(addr[0]), .Z(n32835)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i41_2_lut_rep_820.init = 16'heeee;
    LUT4 mux_1526_i5_rep_77_3_lut (.A(n29712), .B(n32638), .C(n4251), 
         .Z(n29696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i5_rep_77_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_546_4_lut (.A(n32616), .B(n29681), .C(n32656), .D(n32617), 
         .Z(n32561)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_546_4_lut.init = 16'h0200;
    LUT4 i28205_3_lut (.A(n29696), .B(n3328[11]), .C(n30014), .Z(n3446[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28205_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_453 (.A(\addr[1] ), .B(addr[0]), .C(\addr[5] ), 
         .Z(n26838)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_453.init = 16'h1010;
    LUT4 mux_1549_i4_3_lut_rep_642 (.A(n2202[3]), .B(n2222[3]), .C(n32734), 
         .Z(n32657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i4_3_lut_rep_642.init = 16'hcaca;
    LUT4 i28311_2_lut_rep_701_3_lut_4_lut (.A(\addr[1] ), .B(addr[0]), .C(n32836), 
         .D(addr[6]), .Z(n32716)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i28311_2_lut_rep_701_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_454 (.A(n32771), .B(n32762), .C(addr[6]), .D(addr[7]), 
         .Z(n8109)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_454.init = 16'h0200;
    LUT4 i28561_3_lut_rep_739_4_lut (.A(\addr[1] ), .B(addr[0]), .C(addr[2]), 
         .D(n32836), .Z(n32754)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i28561_3_lut_rep_739_4_lut.init = 16'h0001;
    LUT4 is_jalr_N_1372_bdd_2_lut_28839_4_lut (.A(n32616), .B(n29681), .C(n32656), 
         .D(n32570), .Z(n31698)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam is_jalr_N_1372_bdd_2_lut_28839_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_710_3_lut_4_lut (.A(\addr[1] ), .B(addr[0]), .C(n10944), 
         .D(n32836), .Z(n32725)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_710_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_else_4_lut (.A(n8_c), .B(n2202[3]), .C(n28501), .D(n32658), 
         .Z(n32875)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4010;
    LUT4 i1_2_lut_rep_746_3_lut (.A(\addr[1] ), .B(addr[0]), .C(\addr[5] ), 
         .Z(n32761)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_746_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_714_3_lut_4_lut (.A(\addr[1] ), .B(addr[0]), .C(\addr[4] ), 
         .D(\addr[5] ), .Z(n32729)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_2_lut_rep_714_3_lut_4_lut.init = 16'hefff;
    LUT4 i1_2_lut_rep_706_3_lut_4_lut (.A(\addr[1] ), .B(addr[0]), .C(\addr[4] ), 
         .D(\addr[5] ), .Z(n32721)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_2_lut_rep_706_3_lut_4_lut.init = 16'hfeff;
    LUT4 instr_6__I_0_126_i6_2_lut_rep_568_2_lut_4_lut (.A(n2202[3]), .B(n2222[3]), 
         .C(n32734), .D(n32658), .Z(n32583)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_6__I_0_126_i6_2_lut_rep_568_2_lut_4_lut.init = 16'hcaff;
    LUT4 i1_2_lut_4_lut_adj_455 (.A(n2202[3]), .B(n2222[3]), .C(n32734), 
         .D(n34287), .Z(n28435)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_455.init = 16'hca00;
    LUT4 mux_2135_i7_3_lut (.A(n3493[6]), .B(n3446[6]), .C(n32525), .Z(n3534[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2135_i7_3_lut.init = 16'hcaca;
    LUT4 instr_6__I_0_i6_2_lut_rep_603_4_lut (.A(n2202[3]), .B(n2222[3]), 
         .C(n32734), .D(n32658), .Z(n32618)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_6__I_0_i6_2_lut_rep_603_4_lut.init = 16'hffca;
    PFUMX pc_23__I_0_450_i209 (.BLUT(n149_adj_3198), .ALUT(n225_adj_3185), 
          .C0(counter_hi[4]), .Z(n209_adj_3186)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 mux_1549_i3_3_lut_rep_643 (.A(n2202[2]), .B(n2222[2]), .C(n32734), 
         .Z(n32658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i3_3_lut_rep_643.init = 16'hcaca;
    LUT4 mux_2135_i6_3_lut (.A(n3493[5]), .B(n3446[5]), .C(n32525), .Z(n3534[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2135_i6_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_456 (.A(n2202[2]), .B(n2222[2]), .C(n32734), 
         .D(n34287), .Z(n28447)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_456.init = 16'hca00;
    LUT4 mux_2126_i16_3_lut (.A(n3259[12]), .B(n3410[15]), .C(n30007), 
         .Z(n3493[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2126_i16_3_lut.init = 16'hcaca;
    LUT4 i24409_2_lut_rep_588_4_lut (.A(n2202[2]), .B(n2222[2]), .C(n32734), 
         .D(n32661), .Z(n32603)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i24409_2_lut_rep_588_4_lut.init = 16'hca00;
    LUT4 mux_1549_i6_3_lut_rep_644 (.A(n2202[5]), .B(n2222[5]), .C(n32734), 
         .Z(n32659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i6_3_lut_rep_644.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_457 (.A(n2202[5]), .B(n2222[5]), .C(n32734), 
         .D(n32661), .Z(n26879)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_457.init = 16'h00ca;
    LUT4 mux_2126_i15_3_lut (.A(n3259[12]), .B(n3410[14]), .C(n30007), 
         .Z(n3493[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2126_i15_3_lut.init = 16'hcaca;
    LUT4 i28607_2_lut_4_lut (.A(n2202[5]), .B(n2222[5]), .C(n32734), .D(n4265), 
         .Z(n30037)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i28607_2_lut_4_lut.init = 16'hff35;
    LUT4 mux_2126_i14_3_lut (.A(n3259[12]), .B(n3410[13]), .C(n30007), 
         .Z(n3493[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2126_i14_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_823 (.A(alu_op[1]), .B(alu_op[0]), .Z(n32838)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_rep_823.init = 16'hbbbb;
    LUT4 mux_1549_i5_3_lut_rep_646 (.A(n2202[4]), .B(n2222[4]), .C(n32734), 
         .Z(n32661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1549_i5_3_lut_rep_646.init = 16'hcaca;
    LUT4 mux_2126_i13_3_lut (.A(n3259[12]), .B(n3410[12]), .C(n30007), 
         .Z(n3493[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2126_i13_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_592_4_lut (.A(n2202[4]), .B(n2222[4]), .C(n32734), 
         .D(n34287), .Z(n32607)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_592_4_lut.init = 16'hca00;
    LUT4 equal_3528_i7_2_lut_rep_752_3_lut_4_lut (.A(alu_op[1]), .B(alu_op[0]), 
         .C(cycle[1]), .D(\cycle[0] ), .Z(n32767)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam equal_3528_i7_2_lut_rep_752_3_lut_4_lut.init = 16'hfbff;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(alu_op[1]), .B(alu_op[0]), .C(data_rs1[3]), 
         .D(n32848), .Z(n131)) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'he400;
    LUT4 mux_2126_i11_4_lut (.A(n29723), .B(instr[30]), .C(n32525), .D(n9394), 
         .Z(n3493[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2126_i11_4_lut.init = 16'hca0a;
    LUT4 i1_3_lut_4_lut_4_lut_adj_458 (.A(alu_op[1]), .B(alu_op[0]), .C(\cycle[0] ), 
         .D(alu_op_in[2]), .Z(instr_complete_N_1652)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_4_lut_4_lut_adj_458.init = 16'h4be1;
    LUT4 mux_2111_i27_3_lut_4_lut (.A(n32525), .B(n32540), .C(n3446[24]), 
         .D(n29727), .Z(n3446[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2111_i27_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_2_lut_3_lut_adj_459 (.A(n32661), .B(n34287), .C(n32655), .Z(n28561)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_459.init = 16'h0808;
    LUT4 mux_2126_i10_4_lut (.A(n3369[9]), .B(instr[29]), .C(n32525), 
         .D(n9394), .Z(n3493[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2126_i10_4_lut.init = 16'hca0a;
    L6MUX21 mux_2135_i1 (.D0(n3493[0]), .D1(n3446[0]), .SD(n32525), .Z(n3534[0]));
    PFUMX mux_2126_i1 (.BLUT(n3369[0]), .ALUT(n29600), .C0(n4271), .Z(n3493[0]));
    LUT4 i1_3_lut_adj_460 (.A(n32548), .B(n34287), .C(n32541), .Z(clk_c_enable_524)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(35[19:36])
    defparam i1_3_lut_adj_460.init = 16'hc8c8;
    LUT4 mux_1867_i1_4_lut (.A(n2594), .B(n32639), .C(n2798), .D(n32630), 
         .Z(n2618[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam mux_1867_i1_4_lut.init = 16'hca0a;
    LUT4 i15103_3_lut (.A(n2792), .B(n2796), .C(n32638), .Z(n2609[0])) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam i15103_3_lut.init = 16'hc8c8;
    LUT4 i1_4_lut_adj_461 (.A(clk_c_enable_524), .B(n32548), .C(n28523), 
         .D(n32546), .Z(n2126)) /* synthesis lut_function=(A (B+!((D)+!C))) */ ;
    defparam i1_4_lut_adj_461.init = 16'h88a8;
    LUT4 i1_4_lut_adj_462 (.A(n32543), .B(n24_adj_3199), .C(n10024), .D(n29605), 
         .Z(n28523)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_462.init = 16'h0008;
    LUT4 i1_3_lut_adj_463 (.A(mie[2]), .B(n21665), .C(n8_adj_3200), .Z(n793)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_463.init = 16'hcece;
    LUT4 n5568_bdd_3_lut_29217 (.A(counter_hi[2]), .B(instr_data[9]), .C(instr_data[13]), 
         .Z(n32382)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5568_bdd_3_lut_29217.init = 16'he4e4;
    LUT4 instr_len_2__bdd_4_lut (.A(\instr_len[2] ), .B(\pc[1] ), .C(instr_len[1]), 
         .D(\pc[2] ), .Z(next_pc_offset[3])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B (C (D)))) */ ;
    defparam instr_len_2__bdd_4_lut.init = 16'hea80;
    FD1P3AX rs2_i0_i1 (.D(n2302[1]), .SP(clk_c_enable_524), .CK(clk_c), 
            .Q(rs2[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i1.GSR = "DISABLED";
    L6MUX21 i10449 (.D0(n13152), .D1(n3446[3]), .SD(n32525), .Z(n3534[3]));
    PFUMX mux_2135_i21 (.BLUT(n29695), .ALUT(n3446[20]), .C0(n29960), 
          .Z(n3534[20]));
    LUT4 mux_346_i2_3_lut_4_lut (.A(instr_addr_23__N_318[1]), .B(n32682), 
         .C(n32544), .D(return_addr[2]), .Z(n1764[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam mux_346_i2_3_lut_4_lut.init = 16'hf606;
    PFUMX mux_2135_i22 (.BLUT(n29697), .ALUT(n3446[21]), .C0(n29960), 
          .Z(n3534[21]));
    LUT4 data_ready_I_0_3_lut_rep_560 (.A(debug_data_ready), .B(addr[27]), 
         .C(addr_c[26]), .Z(n32575)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(231[27:66])
    defparam data_ready_I_0_3_lut_rep_560.init = 16'h2a2a;
    LUT4 i243_2_lut_4_lut (.A(debug_data_ready), .B(addr[27]), .C(addr_c[26]), 
         .D(load_started), .Z(n824)) /* synthesis lut_function=(!((B (C+!(D))+!B !(D))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(231[27:66])
    defparam i243_2_lut_4_lut.init = 16'h2a00;
    PFUMX mux_2135_i23 (.BLUT(n29705), .ALUT(n3446[22]), .C0(n29960), 
          .Z(n3534[22]));
    LUT4 mux_1867_i4_4_lut (.A(n2590[3]), .B(instr[18]), .C(n2798), .D(n32630), 
         .Z(n2618[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam mux_1867_i4_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_464 (.A(n824), .B(n32549), .C(address_ready), .D(is_load), 
         .Z(clk_c_enable_122)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_464.init = 16'hfeff;
    LUT4 i1_4_lut_adj_465 (.A(n824), .B(n32549), .C(is_load), .D(mem_op[0]), 
         .Z(n27629)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_4_lut_adj_465.init = 16'hffef;
    PFUMX mux_2135_i24 (.BLUT(n29703), .ALUT(n3446[23]), .C0(n29960), 
          .Z(n3534[23]));
    LUT4 mux_2089_i3_4_lut (.A(n29710), .B(n32640), .C(n32540), .D(n32563), 
         .Z(n3328[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2089_i3_4_lut.init = 16'hca0a;
    PFUMX mux_2135_i27 (.BLUT(n29726), .ALUT(n3446[26]), .C0(n29960), 
          .Z(n3534[26]));
    PFUMX mux_2111_i4 (.BLUT(n29704), .ALUT(n3328[3]), .C0(n30084), .Z(n3446[3]));
    FD1P3AX rs2_i0_i2 (.D(n2302[2]), .SP(clk_c_enable_524), .CK(clk_c), 
            .Q(rs2[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i2.GSR = "DISABLED";
    FD1P3AX rs2_i0_i3 (.D(n2302[3]), .SP(clk_c_enable_524), .CK(clk_c), 
            .Q(rs2[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i3.GSR = "DISABLED";
    LUT4 mux_2111_i24_3_lut_4_lut (.A(n32525), .B(n32540), .C(n3446[24]), 
         .D(n29707), .Z(n3446[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2111_i24_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_2089_i4_4_lut (.A(n29707), .B(n32641), .C(n32540), .D(n32563), 
         .Z(n3328[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2089_i4_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_466 (.A(n29105), .B(addr[27]), .C(n29107), .D(n32850), 
         .Z(n7)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_466.init = 16'hfffb;
    PFUMX mux_2111_i3 (.BLUT(n29706), .ALUT(n3328[2]), .C0(n30084), .Z(n3446[2]));
    L6MUX21 mux_2126_i7 (.D0(n3369[6]), .D1(n3410[6]), .SD(n4271), .Z(n3493[6]));
    LUT4 i1_4_lut_adj_467 (.A(\addr[13] ), .B(n29097), .C(n29093), .D(\addr[12] ), 
         .Z(n29105)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_467.init = 16'hfffe;
    L6MUX21 mux_1141_i4 (.D0(n1734[3]), .D1(n1742[3]), .SD(n2126), .Z(n6[3]));
    LUT4 i1_4_lut_adj_468 (.A(\addr[15] ), .B(n29103), .C(n29085), .D(\addr[14] ), 
         .Z(n29107)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_468.init = 16'hfffe;
    L6MUX21 mux_1141_i3 (.D0(n1734[2]), .D1(n1742[2]), .SD(n2126), .Z(n6[2]));
    L6MUX21 mux_1141_i2 (.D0(n1734[1]), .D1(n1742[1]), .SD(n2126), .Z(n6[1]));
    PFUMX mux_1877_i4 (.BLUT(n27567), .ALUT(n2618[3]), .C0(n2800), .Z(n2632[3]));
    LUT4 i1_2_lut_adj_469 (.A(\addr[24] ), .B(\addr[23] ), .Z(n29097)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_adj_469.init = 16'heeee;
    LUT4 i1_2_lut_adj_470 (.A(\addr[18] ), .B(\addr[11] ), .Z(n29093)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_adj_470.init = 16'heeee;
    LUT4 i1_4_lut_adj_471 (.A(\addr[19] ), .B(\addr[21] ), .C(\addr[16] ), 
         .D(\addr[17] ), .Z(n29103)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_471.init = 16'hfffe;
    PFUMX mux_1877_i3 (.BLUT(n27524), .ALUT(n2618[2]), .C0(n2800), .Z(n2632[2]));
    L6MUX21 mux_1877_i2 (.D0(n2609[1]), .D1(n2618[1]), .SD(n2800), .Z(n2632[1]));
    PFUMX i8_adj_472 (.BLUT(n13456), .ALUT(n13458), .C0(clk_c_enable_41), 
          .Z(additional_mem_ops_2__N_749[2]));
    LUT4 n3340_bdd_3_lut_29026_4_lut (.A(\instr[31] ), .B(n32630), .C(n32539), 
         .D(n32026), .Z(n32027)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3340_bdd_3_lut_29026_4_lut.init = 16'hf808;
    PFUMX i10448 (.BLUT(n13151), .ALUT(n3410[3]), .C0(n4271), .Z(n13152));
    FD1P3IX pc_offset__i9 (.D(pc_23__N_911[6]), .SP(clk_c_enable_533), .CD(n32840), 
            .CK(clk_c), .Q(\pc[9] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i9.GSR = "DISABLED";
    PFUMX mux_1877_i1 (.BLUT(n2609[0]), .ALUT(n2618[0]), .C0(n2800), .Z(n2632[0]));
    FD1P3IX pc_offset__i8 (.D(pc_23__N_911[5]), .SP(clk_c_enable_533), .CD(n32840), 
            .CK(clk_c), .Q(\pc[8] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i8.GSR = "DISABLED";
    FD1P3IX pc_offset__i7 (.D(pc_23__N_911[4]), .SP(clk_c_enable_533), .CD(n32840), 
            .CK(clk_c), .Q(\pc[7] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i7.GSR = "DISABLED";
    L6MUX21 mux_2135_i5 (.D0(n3493[4]), .D1(n3446[4]), .SD(n32525), .Z(n3534[4]));
    LUT4 mux_1539_i11_3_lut (.A(n33[10]), .B(n34[10]), .C(n2130), .Z(n2202[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i11_3_lut.init = 16'hcaca;
    FD1P3IX pc_offset__i6 (.D(pc_23__N_911[3]), .SP(clk_c_enable_533), .CD(n32840), 
            .CK(clk_c), .Q(\pc[6] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i6.GSR = "DISABLED";
    L6MUX21 mux_2135_i8 (.D0(n3493[7]), .D1(n3446[7]), .SD(n32525), .Z(n3534[7]));
    FD1P3IX pc_offset__i5 (.D(pc_23__N_911[2]), .SP(clk_c_enable_533), .CD(n32840), 
            .CK(clk_c), .Q(\pc[5] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i5.GSR = "DISABLED";
    PFUMX mux_2135_i9 (.BLUT(n3410[8]), .ALUT(n3493[8]), .C0(n30032), 
          .Z(n3534[8]));
    LUT4 i15294_3_lut_4_lut (.A(n32595), .B(n32656), .C(n32639), .D(n32655), 
         .Z(n29_c)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (D)))) */ ;
    defparam i15294_3_lut_4_lut.init = 16'h001f;
    LUT4 i1_2_lut_rep_826 (.A(\instr_len[2] ), .B(\pc[2] ), .Z(n32841)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_2_lut_rep_826.init = 16'h6666;
    PFUMX mux_2135_i10 (.BLUT(n3410[9]), .ALUT(n3493[9]), .C0(n30032), 
          .Z(n3534[9]));
    LUT4 i1_2_lut_adj_473 (.A(\addr[22] ), .B(\addr[20] ), .Z(n29085)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_adj_473.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_474 (.A(\instr_len[2] ), .B(\pc[2] ), .C(instr_addr_23__N_318[1]), 
         .Z(n28971)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_2_lut_3_lut_adj_474.init = 16'h9696;
    LUT4 i28601_3_lut_rep_670_4_lut (.A(n32851), .B(addr[10]), .C(n7), 
         .D(n27178), .Z(n32685)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;
    defparam i28601_3_lut_rep_670_4_lut.init = 16'h0f0d;
    LUT4 i1536_3_lut_rep_719_4_lut_4_lut (.A(\instr_len[2] ), .B(\pc[2] ), 
         .C(n34285), .D(n32842), .Z(n32734)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C (D))+!B !(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1536_3_lut_rep_719_4_lut_4_lut.init = 16'h9c6c;
    LUT4 i4408_2_lut_rep_827 (.A(\pc[1] ), .B(instr_len[1]), .Z(n32842)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i4408_2_lut_rep_827.init = 16'h8888;
    LUT4 i2_2_lut_rep_751_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), .C(\pc[2] ), 
         .D(\instr_len[2] ), .Z(n32766)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i2_2_lut_rep_751_3_lut_4_lut.init = 16'h8778;
    PFUMX mux_2135_i11 (.BLUT(n3410[10]), .ALUT(n3493[10]), .C0(n30024), 
          .Z(n3534[10]));
    LUT4 i4406_2_lut_rep_828 (.A(\pc[1] ), .B(instr_len[1]), .Z(n32843)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i4406_2_lut_rep_828.init = 16'h6666;
    LUT4 i27127_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), .C(counter_hi[2]), 
         .D(\next_pc_for_core[5] ), .Z(n29836)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i27127_3_lut_4_lut.init = 16'hf606;
    LUT4 i1_4_lut_4_lut_adj_475 (.A(\pc[1] ), .B(instr_len[1]), .C(n34285), 
         .D(\instr_addr_23__N_318[0] ), .Z(n10253)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_4_lut_4_lut_adj_475.init = 16'h956a;
    LUT4 i4818_2_lut_rep_736_3_lut (.A(\pc[1] ), .B(instr_len[1]), .C(\instr_addr_23__N_318[0] ), 
         .Z(n32751)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i4818_2_lut_rep_736_3_lut.init = 16'hf9f9;
    LUT4 mux_347_i1_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), .C(n32544), 
         .D(return_addr[1]), .Z(n1768[0])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam mux_347_i1_3_lut_4_lut.init = 16'hf606;
    FD1P3IX pc_offset__i4 (.D(pc_23__N_911[1]), .SP(clk_c_enable_533), .CD(n32840), 
            .CK(clk_c), .Q(\pc[4] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i4.GSR = "DISABLED";
    PFUMX mux_2135_i12 (.BLUT(n3493[11]), .ALUT(n3446[11]), .C0(n32525), 
          .Z(n3534[11]));
    PFUMX mux_2135_i13 (.BLUT(n3493[12]), .ALUT(n3446[12]), .C0(n32525), 
          .Z(n3534[12]));
    PFUMX mux_2135_i14 (.BLUT(n3493[13]), .ALUT(n3446[13]), .C0(n32525), 
          .Z(n3534[13]));
    PFUMX mux_2135_i15 (.BLUT(n3493[14]), .ALUT(n3446[14]), .C0(n32525), 
          .Z(n3534[14]));
    LUT4 mux_1543_i11_3_lut (.A(n36[10]), .B(n31[10]), .C(n2150), .Z(n2222[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i11_3_lut.init = 16'hcaca;
    PFUMX i27546 (.BLUT(n30251), .ALUT(n30252), .C0(counter_hi[3]), .Z(n30255));
    PFUMX mux_2135_i16 (.BLUT(n3493[15]), .ALUT(n3446[15]), .C0(n32525), 
          .Z(n3534[15]));
    L6MUX21 mux_2135_i17 (.D0(n3493[16]), .D1(n3446[16]), .SD(n32525), 
            .Z(n3534[16]));
    LUT4 is_system_I_0_481_2_lut_rep_831 (.A(is_system), .B(n34285), .Z(n32846)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam is_system_I_0_481_2_lut_rep_831.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_476 (.A(rst_reg_n_adj_6), .B(clk_c_enable_41), 
         .C(n43), .D(n32630), .Z(n2122)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(35[19:36])
    defparam i1_3_lut_4_lut_adj_476.init = 16'h8880;
    LUT4 mux_2135_i3_3_lut (.A(n3493[2]), .B(n3446[2]), .C(n32525), .Z(n3534[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2135_i3_3_lut.init = 16'hcaca;
    LUT4 i28268_4_lut (.A(n32552), .B(rst_reg_n_adj_6), .C(n32544), .D(n28475), 
         .Z(clk_c_enable_309)) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;
    defparam i28268_4_lut.init = 16'h3733;
    FD1P3IX pc_offset__i3 (.D(pc_23__N_911[0]), .SP(clk_c_enable_533), .CD(n32840), 
            .CK(clk_c), .Q(\pc[3] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i3.GSR = "DISABLED";
    FD1P3IX pc_offset__i2 (.D(pc_2__N_932[1]), .SP(clk_c_enable_533), .CD(n32840), 
            .CK(clk_c), .Q(\pc[2] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i2.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_477 (.A(is_system), .B(debug_instr_valid), .C(\imm[6] ), 
         .D(n32847), .Z(n24384)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_3_lut_4_lut_adj_477.init = 16'h8000;
    PFUMX mux_2135_i28 (.BLUT(n5205[27]), .ALUT(n3446[27]), .C0(n29917), 
          .Z(n3534[27]));
    LUT4 i1_3_lut_rep_753_4_lut (.A(is_system), .B(n34285), .C(n32847), 
         .D(alu_op_in[2]), .Z(n32768)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_3_lut_rep_753_4_lut.init = 16'h0008;
    PFUMX mux_2135_i31 (.BLUT(n5205[30]), .ALUT(n3446[30]), .C0(n29917), 
          .Z(n3534[30]));
    LUT4 i15132_2_lut (.A(\pc[4] ), .B(counter_hi[2]), .Z(n149_adj_3198)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam i15132_2_lut.init = 16'h8888;
    PFUMX mux_1131_i4 (.BLUT(n27546), .ALUT(n1708[3]), .C0(n2122), .Z(n1734[3]));
    LUT4 i1_4_lut_adj_478 (.A(n19_adj_3201), .B(n28731), .C(n32623), .D(n672), 
         .Z(n28733)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A ((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_478.init = 16'h0c88;
    PFUMX mux_1131_i3 (.BLUT(n27541), .ALUT(n1708[2]), .C0(n2122), .Z(n1734[2]));
    PFUMX mux_1131_i2 (.BLUT(n27545), .ALUT(n1708[1]), .C0(n2122), .Z(n1734[1]));
    PFUMX mux_2111_i17 (.BLUT(n3328[16]), .ALUT(n5205[16]), .C0(n32540), 
          .Z(n3446[16]));
    LUT4 i15000_3_lut (.A(n32783), .B(rst_reg_n_adj_6), .C(n32547), .Z(data_continue_N_963)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i15000_3_lut.init = 16'ha8a8;
    PFUMX mux_2111_i5 (.BLUT(n3328[4]), .ALUT(n5205[4]), .C0(n32540), 
          .Z(n3446[4]));
    LUT4 i1_2_lut_rep_835 (.A(addr_c[26]), .B(addr_c[25]), .Z(n32850)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_835.init = 16'heeee;
    PFUMX mux_2126_i17 (.BLUT(n3259[16]), .ALUT(n3410[16]), .C0(n30007), 
          .Z(n3493[16]));
    LUT4 i1_rep_143_2_lut_3_lut (.A(addr_c[26]), .B(addr_c[25]), .C(addr[27]), 
         .Z(n30929)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_rep_143_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_rep_144_2_lut_3_lut (.A(addr_c[26]), .B(addr_c[25]), .C(addr[27]), 
         .Z(n30930)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_rep_144_2_lut_3_lut.init = 16'hfefe;
    LUT4 i15638_2_lut_rep_696_3_lut_4_lut (.A(addr_c[26]), .B(addr_c[25]), 
         .C(n21414), .D(addr[27]), .Z(n32711)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i15638_2_lut_rep_696_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_756_3_lut (.A(addr_c[26]), .B(addr_c[25]), .C(addr[27]), 
         .Z(n32771)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_756_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_722_3_lut_4_lut (.A(addr_c[26]), .B(addr_c[25]), .C(n21414), 
         .D(addr[27]), .Z(n32737)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_722_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i28571_2_lut_rep_720_3_lut_4_lut (.A(addr_c[26]), .B(addr_c[25]), 
         .C(counter_hi[4]), .D(addr[27]), .Z(n32735)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i28571_2_lut_rep_720_3_lut_4_lut.init = 16'hffef;
    PFUMX mux_2126_i8 (.BLUT(n3369[7]), .ALUT(n3410[7]), .C0(n4271), .Z(n3493[7]));
    LUT4 i28308_2_lut_rep_836 (.A(\addr[8] ), .B(\addr[9] ), .Z(n32851)) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i28308_2_lut_rep_836.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_adj_479 (.A(\addr[8] ), .B(\addr[9] ), .C(n32255), 
         .Z(\data_from_peri_31__N_2415[0] )) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_adj_479.init = 16'h1010;
    LUT4 i1_2_lut_rep_747_3_lut (.A(\addr[8] ), .B(\addr[9] ), .C(addr[10]), 
         .Z(n32762)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_747_3_lut.init = 16'hfefe;
    LUT4 i6_3_lut_3_lut_4_lut (.A(n32654), .B(n24900), .C(n32548), .D(n32227), 
         .Z(n13458)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D))+!B !(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i6_3_lut_3_lut_4_lut.init = 16'hb444;
    L6MUX21 mux_2126_i6 (.D0(n3369[5]), .D1(n3410[5]), .SD(n4271), .Z(n3493[5]));
    PFUMX mux_2126_i5 (.BLUT(n3369[4]), .ALUT(n3410[4]), .C0(n4271), .Z(n3493[4]));
    LUT4 i4337_2_lut_rep_838 (.A(rs2[0]), .B(mem_op_increment_reg), .Z(n32853)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i4337_2_lut_rep_838.init = 16'h8888;
    LUT4 fsm_state_0__bdd_4_lut_29703 (.A(fsm_state[0]), .B(n32778), .C(fsm_state[1]), 
         .D(fsm_state[2]), .Z(n31866)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (B+!(C (D)+!C !(D))))) */ ;
    defparam fsm_state_0__bdd_4_lut_29703.init = 16'h3203;
    LUT4 i28293_3_lut_4_lut (.A(n32693), .B(n32721), .C(rst_reg_n), .D(n10944), 
         .Z(clk_c_enable_50)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;
    defparam i28293_3_lut_4_lut.init = 16'h0f1f;
    L6MUX21 mux_2126_i3 (.D0(n3369[2]), .D1(n3410[2]), .SD(n4271), .Z(n3493[2]));
    PFUMX mux_1135_i4 (.BLUT(n1713[3]), .ALUT(n27657), .C0(n2124), .Z(n1742[3]));
    LUT4 i4345_2_lut_rep_758_3_lut (.A(rs2[0]), .B(mem_op_increment_reg), 
         .C(rs2[1]), .Z(n32773)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i4345_2_lut_rep_758_3_lut.init = 16'h8080;
    LUT4 i28419_3_lut_4_lut (.A(n32693), .B(n32721), .C(rst_reg_n), .D(n32818), 
         .Z(clk_c_enable_154)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;
    defparam i28419_3_lut_4_lut.init = 16'h0f1f;
    PFUMX mux_1135_i3 (.BLUT(n1713[2]), .ALUT(n27655), .C0(n2124), .Z(n1742[2]));
    LUT4 i28288_3_lut_4_lut (.A(n32693), .B(n32721), .C(rst_reg_n), .D(n32819), 
         .Z(clk_c_enable_283)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;
    defparam i28288_3_lut_4_lut.init = 16'h0f1f;
    PFUMX mux_1135_i2 (.BLUT(n1713[1]), .ALUT(n27656), .C0(n2124), .Z(n1742[1]));
    LUT4 i4352_2_lut_3_lut_4_lut (.A(rs2[0]), .B(mem_op_increment_reg), 
         .C(rs2[2]), .D(rs2[1]), .Z(n6634)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i4352_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i28263_3_lut_4_lut (.A(n32693), .B(n32721), .C(rst_reg_n), .D(n8854), 
         .Z(clk_c_enable_354)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !((D)+!C)))) */ ;
    defparam i28263_3_lut_4_lut.init = 16'h1f0f;
    LUT4 \gpio_out_func_sel_0[[2__bdd_3_lut_29665  (.A(\gpio_out_func_sel[0][2] ), 
         .B(addr[2]), .C(\gpio_out_func_sel[1][2] ), .Z(n31881)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam \gpio_out_func_sel_0[[2__bdd_3_lut_29665 .init = 16'he2e2;
    LUT4 \gpio_out_func_sel_0[[2__bdd_3_lut_28962  (.A(\gpio_out_func_sel[2][2] ), 
         .B(addr[2]), .C(\gpio_out_func_sel[3][2] ), .Z(n31880)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam \gpio_out_func_sel_0[[2__bdd_3_lut_28962 .init = 16'he2e2;
    LUT4 i15185_2_lut_4_lut_4_lut (.A(n7), .B(n32694), .C(n32756), .D(\addr[4] ), 
         .Z(n5169)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i15185_2_lut_4_lut_4_lut.init = 16'h5040;
    PFUMX mux_2098_i7 (.BLUT(n13165), .ALUT(n3183[6]), .C0(n30037), .Z(n3369[6]));
    PFUMX i27547 (.BLUT(n30253), .ALUT(n30254), .C0(counter_hi[3]), .Z(n30256));
    LUT4 i4787_2_lut (.A(\instr_addr_23__N_318[0] ), .B(\pc[1] ), .Z(n2_adj_3202)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i4787_2_lut.init = 16'hbbbb;
    LUT4 i1_3_lut_adj_480 (.A(next_pc_offset[3]), .B(n4_adj_3203), .C(\instr_write_offset[3] ), 
         .Z(n27804)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i1_3_lut_adj_480.init = 16'h9696;
    LUT4 i15300_2_lut_3_lut (.A(n32654), .B(n32655), .C(n32653), .Z(n17949)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i15300_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_481 (.A(debug_early_branch), .B(n32544), .C(n32551), 
         .D(n29618), .Z(start_instr)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_481.init = 16'h0010;
    PFUMX mux_1867_i2 (.BLUT(n11066), .ALUT(n2595[1]), .C0(n2798), .Z(n2618[1]));
    LUT4 i15796_4_lut_4_lut (.A(n7), .B(n32694), .C(n32825), .D(n29127), 
         .Z(n18458)) /* synthesis lut_function=(!(A+!(B+(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i15796_4_lut_4_lut.init = 16'h5444;
    L6MUX21 i10452 (.D0(n13155), .D1(n3410[1]), .SD(n4271), .Z(n13156));
    PFUMX mux_1575_i1 (.BLUT(n2291[0]), .ALUT(n2281[0]), .C0(n2559), .Z(n2302[0]));
    LUT4 n29834_bdd_3_lut_29686 (.A(\gpio_out_func_sel[4][2] ), .B(addr[3]), 
         .C(\gpio_out_func_sel[6][2] ), .Z(n31878)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n29834_bdd_3_lut_29686.init = 16'he2e2;
    PFUMX mux_1575_i2 (.BLUT(n2291[1]), .ALUT(n2281[1]), .C0(n2559), .Z(n2302[1]));
    PFUMX i27553 (.BLUT(n30258), .ALUT(n30259), .C0(counter_hi[3]), .Z(n30262));
    PFUMX mux_1575_i3 (.BLUT(n2291[2]), .ALUT(n2281[2]), .C0(n2559), .Z(n2302[2]));
    PFUMX mux_1575_i4 (.BLUT(n2291[3]), .ALUT(n2281[3]), .C0(n2559), .Z(n2302[3]));
    FD1P3IX instr_valid_392_rep_848 (.D(debug_instr_valid_N_436), .SP(clk_c_enable_545), 
            .CD(n32840), .CK(clk_c), .Q(n34285)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_valid_392_rep_848.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_482 (.A(n32545), .B(n8), .C(n32552), .D(n28873), 
         .Z(debug_early_branch)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_482.init = 16'h0200;
    LUT4 mux_2111_i23_3_lut_4_lut (.A(n32525), .B(n32540), .C(n3446[24]), 
         .D(n29710), .Z(n3446[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2111_i23_3_lut_4_lut.init = 16'hf870;
    PFUMX mux_2107_i7 (.BLUT(n3259[6]), .ALUT(n3292[6]), .C0(n4267), .Z(n3410[6]));
    LUT4 i14598_3_lut (.A(\uart_rx_buf_data[4] ), .B(\baud_divider[4] ), 
         .C(addr[3]), .Z(n15_adj_3188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i14598_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_483 (.A(n27003), .B(n27585), .C(instr_fetch_running_N_945), 
         .D(instr_fetch_stopped), .Z(clk_c_enable_367)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_483.init = 16'hfffd;
    PFUMX mux_2107_i6 (.BLUT(n3259[5]), .ALUT(n3292[5]), .C0(n4267), .Z(n3410[5]));
    LUT4 i14913_4_lut (.A(n16), .B(rst_reg_n_adj_6), .C(was_early_branch), 
         .D(n32552), .Z(n6396)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam i14913_4_lut.init = 16'hc088;
    LUT4 i1_3_lut_adj_484 (.A(is_jal_de), .B(n34287), .C(is_ret_de), .Z(n28685)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut_adj_484.init = 16'hc8c8;
    PFUMX mux_2107_i3 (.BLUT(n3259[2]), .ALUT(n3292[2]), .C0(n4267), .Z(n3410[2]));
    LUT4 i1_2_lut_adj_485 (.A(is_jal_de), .B(n34287), .Z(n28873)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_485.init = 16'h8888;
    PFUMX mux_2107_i2 (.BLUT(n3259[1]), .ALUT(n3292[1]), .C0(n4267), .Z(n3410[1]));
    PFUMX i27554 (.BLUT(n30260), .ALUT(n30261), .C0(counter_hi[3]), .Z(n30263));
    PFUMX mux_2126_i19 (.BLUT(n3259[17]), .ALUT(n3410[17]), .C0(n30197), 
          .Z(n3493[17]));
    PFUMX mux_2098_i6 (.BLUT(n3183[5]), .ALUT(n27483), .C0(n4265), .Z(n3369[5]));
    PFUMX mux_2098_i3 (.BLUT(n3183[2]), .ALUT(n27356), .C0(n4265), .Z(n3369[2]));
    PFUMX mux_2111_i1 (.BLUT(n27731), .ALUT(n5205[0]), .C0(n32540), .Z(n3446[0]));
    LUT4 i17356_4_lut (.A(data_to_write[3]), .B(instr_data[11]), .C(qspi_data_ready), 
         .D(n32826), .Z(\instr_data_7__N_1969[3] )) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i17356_4_lut.init = 16'h0aca;
    LUT4 mux_1520_i13_3_lut (.A(n31[12]), .B(n33[12]), .C(n2150), .Z(n2151[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1516_i13_3_lut (.A(n34[12]), .B(n36[12]), .C(n2130), .Z(n2131[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i13_3_lut.init = 16'hcaca;
    LUT4 i17350_4_lut (.A(data_to_write[1]), .B(instr_data[9]), .C(qspi_data_ready), 
         .D(n32826), .Z(\instr_data_7__N_1969[1] )) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i17350_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_adj_486 (.A(n32545), .B(n27003), .C(n8), .D(n28827), 
         .Z(n26962)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B))) */ ;
    defparam i1_4_lut_adj_486.init = 16'h3b33;
    LUT4 no_write_in_progress_I_42_4_lut (.A(n29173), .B(addr_out[27]), 
         .C(n32692), .D(n32575), .Z(no_write_in_progress_N_471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(279[18] 289[12])
    defparam no_write_in_progress_I_42_4_lut.init = 16'hcfca;
    PFUMX i10451 (.BLUT(n13154), .ALUT(n3222[1]), .C0(n4265), .Z(n13155));
    LUT4 pc_23__I_0_450_i157_3_lut (.A(\pc[8] ), .B(\pc[12] ), .C(counter_hi[2]), 
         .Z(n157_adj_3187)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam pc_23__I_0_450_i157_3_lut.init = 16'hcaca;
    LUT4 i28178_3_lut_4_lut (.A(n32530), .B(n32637), .C(n4265), .D(n27492), 
         .Z(n3369[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i28178_3_lut_4_lut.init = 16'hf808;
    PFUMX i32 (.BLUT(n27427), .ALUT(n29594), .C0(n32659), .Z(n13_adj_3170));
    LUT4 i4638_2_lut_3_lut (.A(n32707), .B(\instr_addr_23__N_318[0] ), .C(instr_addr_23__N_318[1]), 
         .Z(n6920)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i4638_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_2084_i15_3_lut_4_lut (.A(n32642), .B(n32608), .C(n4267), 
         .D(n29723), .Z(n3259[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2084_i15_3_lut_4_lut.init = 16'h8f80;
    LUT4 next_instr_write_offset_3__I_0_i2_2_lut_3_lut_4_lut (.A(n32707), 
         .B(\instr_addr_23__N_318[0] ), .C(\pc[2] ), .D(instr_addr_23__N_318[1]), 
         .Z(n2_c)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam next_instr_write_offset_3__I_0_i2_2_lut_3_lut_4_lut.init = 16'h8778;
    LUT4 next_instr_write_offset_3__I_0_i1_2_lut_3_lut (.A(n32707), .B(\instr_addr_23__N_318[0] ), 
         .C(\pc[1] ), .Z(n1_c)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam next_instr_write_offset_3__I_0_i1_2_lut_3_lut.init = 16'h9696;
    LUT4 mux_2084_i17_3_lut_4_lut (.A(n32642), .B(n32608), .C(n4267), 
         .D(n2970[16]), .Z(n3259[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2084_i17_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_346_i1_3_lut_4_lut (.A(n32707), .B(\instr_addr_23__N_318[0] ), 
         .C(n32544), .D(return_addr[1]), .Z(n1764[0])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam mux_346_i1_3_lut_4_lut.init = 16'hf606;
    LUT4 i1_4_lut_adj_487 (.A(n32549), .B(n27653), .C(n32546), .D(n28851), 
         .Z(clk_c_enable_545)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;
    defparam i1_4_lut_adj_487.init = 16'h3332;
    LUT4 mux_2084_i9_3_lut_4_lut (.A(n32642), .B(n32608), .C(n4267), .D(n2590[2]), 
         .Z(n3259[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2084_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2084_i10_3_lut_4_lut (.A(n32642), .B(n32608), .C(n4267), 
         .D(n2590[3]), .Z(n3259[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2084_i10_3_lut_4_lut.init = 16'h8f80;
    PFUMX mux_2111_i7 (.BLUT(n29725), .ALUT(n3328[6]), .C0(n30041), .Z(n3446[6]));
    PFUMX mux_2084_i8 (.BLUT(n5138[6]), .ALUT(n2970[7]), .C0(n4259), .Z(n3259[7]));
    LUT4 i1_2_lut_rep_515 (.A(n13140), .B(n4243), .Z(n32530)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_515.init = 16'heeee;
    LUT4 mux_2107_i19_3_lut_3_lut_4_lut (.A(n32642), .B(n32608), .C(n3369[11]), 
         .D(n4271), .Z(n3410[17])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2107_i19_3_lut_3_lut_4_lut.init = 16'h88f0;
    LUT4 i1_2_lut_4_lut_adj_488 (.A(n27178), .B(n7), .C(n32762), .D(gpio_out_sel[6]), 
         .Z(n14)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_2_lut_4_lut_adj_488.init = 16'hff32;
    LUT4 i1_2_lut_4_lut_adj_489 (.A(n27178), .B(n7), .C(n32762), .D(gpio_out_sel[7]), 
         .Z(n14_adj_8)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_2_lut_4_lut_adj_489.init = 16'hff32;
    LUT4 i24415_2_lut_4_lut (.A(n27178), .B(n7), .C(n32762), .D(\addr[4] ), 
         .Z(n26988)) /* synthesis lut_function=(A (B+(D))+!A (B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i24415_2_lut_4_lut.init = 16'hffcd;
    LUT4 i1_2_lut_4_lut_adj_490 (.A(n27178), .B(n7), .C(n32762), .D(n32728), 
         .Z(n29293)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B (D)+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_2_lut_4_lut_adj_490.init = 16'h00cd;
    PFUMX mux_2084_i5 (.BLUT(n5138[3]), .ALUT(n2970[4]), .C0(n4259), .Z(n3259[4]));
    PFUMX mux_2098_i10 (.BLUT(n27430), .ALUT(n27486), .C0(n4265), .Z(n3369[9]));
    LUT4 mux_1539_i10_3_lut (.A(n33[9]), .B(n34[9]), .C(n2130), .Z(n2202[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i10_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_491 (.A(n35), .B(n10772), .Z(n4265)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_491.init = 16'h8888;
    PFUMX mux_2098_i9 (.BLUT(n27428), .ALUT(n27495), .C0(n4265), .Z(n3369[8]));
    LUT4 i21713_2_lut (.A(counter_hi[3]), .B(counter_hi[2]), .Z(n39[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i21713_2_lut.init = 16'h6666;
    LUT4 i21734_4_lut (.A(n58), .B(n28963), .C(addr_offset[3]), .D(instr_complete_N_1647), 
         .Z(n38[1])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i21734_4_lut.init = 16'h6ca0;
    PFUMX i29383 (.BLUT(n32990), .ALUT(\data_from_read[6] ), .C0(n30930), 
          .Z(n32991));
    LUT4 i43_3_lut_4_lut (.A(n32628), .B(n32602), .C(n32653), .D(n23), 
         .Z(n26)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam i43_3_lut_4_lut.init = 16'h2f20;
    PFUMX mux_1862_i2 (.BLUT(n2577[1]), .ALUT(n2585[1]), .C0(n2796), .Z(n2609[1]));
    LUT4 pc_23__I_0_450_i269_3_lut (.A(n209_adj_3186), .B(data_rs1[0]), 
         .C(n32806), .Z(debug_branch_N_442[28])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam pc_23__I_0_450_i269_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_adj_492 (.A(n13140), .B(n4243), .C(n32651), .Z(n3183[2])) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_492.init = 16'he0e0;
    LUT4 i10450_1_lut_2_lut (.A(n13140), .B(n4243), .Z(n13154)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i10450_1_lut_2_lut.init = 16'h1111;
    LUT4 i28532_4_lut (.A(n32552), .B(n32546), .C(n10024), .D(is_ret_de), 
         .Z(debug_instr_valid_N_436)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i28532_4_lut.init = 16'h0001;
    LUT4 i6371_4_lut_4_lut (.A(n32654), .B(n155[3]), .C(n30), .D(n29119), 
         .Z(n9052)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i6371_4_lut_4_lut.init = 16'hd850;
    LUT4 i15345_2_lut_3_lut (.A(n13140), .B(n4243), .C(n32642), .Z(n3183[5])) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i15345_2_lut_3_lut.init = 16'he0e0;
    LUT4 n23_bdd_3_lut_3_lut (.A(n32654), .B(n32639), .C(n32656), .Z(n32487)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam n23_bdd_3_lut_3_lut.init = 16'h1414;
    LUT4 i10461_4_lut_4_lut (.A(n13140), .B(n4243), .C(n1_adj_3208), .D(n32638), 
         .Z(n13165)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B (C+(D)))) */ ;
    defparam i10461_4_lut_4_lut.init = 16'heec0;
    LUT4 mux_2111_i22_3_lut_4_lut (.A(n32525), .B(n32540), .C(n3446[24]), 
         .D(n29702), .Z(n3446[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2111_i22_3_lut_4_lut.init = 16'hf870;
    LUT4 is_store_I_0_469_2_lut_rep_677 (.A(is_store), .B(address_ready), 
         .Z(n32692)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(275[22:47])
    defparam is_store_I_0_469_2_lut_rep_677.init = 16'h8888;
    LUT4 i1_4_lut_rep_529 (.A(n32545), .B(n8), .C(n32552), .D(n28827), 
         .Z(n32544)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_rep_529.init = 16'h0200;
    LUT4 n32018_bdd_3_lut (.A(n32016), .B(\instr[31] ), .C(n4251), .Z(n32019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n32018_bdd_3_lut.init = 16'hcaca;
    LUT4 n32179_bdd_3_lut_3_lut (.A(n32654), .B(n32178), .C(n32179), .Z(n32180)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam n32179_bdd_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_4_lut_adj_493 (.A(n32671), .B(n32575), .C(data_ready_sync), 
         .D(clk_c_enable_285), .Z(clk_c_enable_513)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_493.init = 16'hfeee;
    LUT4 i1_4_lut_adj_494 (.A(n824), .B(n32549), .C(is_load), .D(mem_op[1]), 
         .Z(n27630)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_4_lut_adj_494.init = 16'hffef;
    LUT4 i1_2_lut_3_lut_4_lut_adj_495 (.A(is_store), .B(address_ready), 
         .C(mem_op[0]), .D(rst_reg_n_adj_6), .Z(data_write_n_1__N_369[0])) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(275[22:47])
    defparam i1_2_lut_3_lut_4_lut_adj_495.init = 16'hf7ff;
    LUT4 i1_2_lut_3_lut_4_lut_adj_496 (.A(is_store), .B(address_ready), 
         .C(mem_op[1]), .D(rst_reg_n_adj_6), .Z(data_write_n_1__N_369[1])) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(275[22:47])
    defparam i1_2_lut_3_lut_4_lut_adj_496.init = 16'hf7ff;
    PFUMX mux_2111_i8 (.BLUT(n3328[7]), .ALUT(n5205[7]), .C0(n32540), 
          .Z(n3446[7]));
    PFUMX mux_2111_i6 (.BLUT(n3328[5]), .ALUT(n5205[5]), .C0(n32540), 
          .Z(n3446[5]));
    LUT4 i2_2_lut_rep_657_3_lut (.A(addr[7]), .B(n32723), .C(n7), .Z(n32672)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i2_2_lut_rep_657_3_lut.init = 16'hfefe;
    PFUMX mux_833_i21 (.BLUT(n1742_adj_3219[20]), .ALUT(n1203[20]), .C0(n30928), 
          .Z(pc_23__N_911[20]));
    LUT4 i28576_2_lut_3_lut_4_lut (.A(addr[7]), .B(n32723), .C(\addr[4] ), 
         .D(n7), .Z(n4)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i28576_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i6177_3_lut_3_lut_4_lut (.A(addr[7]), .B(n32723), .C(n8854), 
         .D(n7), .Z(n19)) /* synthesis lut_function=(A (D)+!A (B (D)+!B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i6177_3_lut_3_lut_4_lut.init = 16'hff01;
    LUT4 i1_2_lut_3_lut_4_lut_adj_497 (.A(addr[7]), .B(n32723), .C(\addr[4] ), 
         .D(n7), .Z(n46)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_4_lut_adj_497.init = 16'h0010;
    PFUMX mux_833_i20 (.BLUT(n1742_adj_3219[19]), .ALUT(n1203[19]), .C0(n30928), 
          .Z(pc_23__N_911[19]));
    LUT4 connect_peripheral_3__I_1_i2_3_lut_3_lut_4_lut (.A(addr[7]), .B(n32723), 
         .C(addr[3]), .D(n7), .Z(\connect_peripheral[1] )) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam connect_peripheral_3__I_1_i2_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 connect_peripheral_3__I_1_i1_3_lut_3_lut_4_lut (.A(addr[7]), .B(n32723), 
         .C(addr[2]), .D(n7), .Z(\connect_peripheral[0] )) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam connect_peripheral_3__I_1_i1_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 connect_peripheral_3__I_1_i3_3_lut_rep_645_3_lut_4_lut (.A(addr[7]), 
         .B(n32723), .C(\addr[4] ), .D(n7), .Z(n32660)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam connect_peripheral_3__I_1_i3_3_lut_rep_645_3_lut_4_lut.init = 16'h00fe;
    LUT4 n2166_bdd_3_lut (.A(n2151[1]), .B(n32734), .C(n29745), .Z(n32016)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n2166_bdd_3_lut.init = 16'hb8b8;
    LUT4 n5568_bdd_3_lut_29221 (.A(counter_hi[2]), .B(\qspi_data_buf[9] ), 
         .C(\qspi_data_buf[13] ), .Z(n32383)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5568_bdd_3_lut_29221.init = 16'he4e4;
    LUT4 i1_4_lut_adj_498 (.A(addr_out[3]), .B(n32690), .C(addr_offset[3]), 
         .D(addr_offset[2]), .Z(n27823)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(121[15:26])
    defparam i1_4_lut_adj_498.init = 16'h965a;
    PFUMX mux_833_i19 (.BLUT(n1742_adj_3219[18]), .ALUT(n1203[18]), .C0(n30928), 
          .Z(pc_23__N_911[18]));
    PFUMX mux_833_i18 (.BLUT(n1742_adj_3219[17]), .ALUT(n1203[17]), .C0(n30928), 
          .Z(pc_23__N_911[17]));
    FD1S3IX counter_hi_3544__i3_rep_846 (.D(n39[1]), .CK(clk_c), .CD(n32840), 
            .Q(n34283));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3544__i3_rep_846.GSR = "DISABLED";
    LUT4 instr_addr_23__I_0_i2_3_lut (.A(instr_addr_23__N_318[1]), .B(\early_branch_addr[2] ), 
         .C(was_early_branch), .Z(\instr_addr[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[25:119])
    defparam instr_addr_23__I_0_i2_3_lut.init = 16'hcaca;
    PFUMX mux_833_i17 (.BLUT(n1742_adj_3219[16]), .ALUT(n1203[16]), .C0(n30927), 
          .Z(pc_23__N_911[16]));
    LUT4 i21726_3_lut (.A(n32548), .B(n58), .C(addr_offset[2]), .Z(n38[0])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i21726_3_lut.init = 16'h6a6a;
    LUT4 n3508_bdd_3_lut_29024 (.A(n3493[17]), .B(n32021), .C(n32525), 
         .Z(n32022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3508_bdd_3_lut_29024.init = 16'hcaca;
    LUT4 i1_4_lut_adj_499 (.A(n32546), .B(n32543), .C(n32548), .D(n10024), 
         .Z(n58)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_499.init = 16'hfffb;
    LUT4 n4251_bdd_3_lut_29036 (.A(n2151[2]), .B(n32734), .C(n29743), 
         .Z(n32025)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n4251_bdd_3_lut_29036.init = 16'hb8b8;
    PFUMX mux_833_i16 (.BLUT(n1742_adj_3219[15]), .ALUT(n1203[15]), .C0(n30927), 
          .Z(pc_23__N_911[15]));
    PFUMX mux_833_i15 (.BLUT(n1742_adj_3219[14]), .ALUT(n1203[14]), .C0(n30927), 
          .Z(pc_23__N_911[14]));
    PFUMX mux_833_i13 (.BLUT(n1742_adj_3219[12]), .ALUT(n1203[12]), .C0(n30927), 
          .Z(pc_23__N_911[12]));
    LUT4 i1_3_lut_4_lut_adj_500 (.A(n32774), .B(n32549), .C(n28685), .D(n8), 
         .Z(n27585)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[22:78])
    defparam i1_3_lut_4_lut_adj_500.init = 16'h00d0;
    PFUMX mux_833_i12 (.BLUT(n1742_adj_3219[11]), .ALUT(n1203[11]), .C0(n30926), 
          .Z(pc_23__N_911[11]));
    LUT4 i1_3_lut_adj_501 (.A(debug_early_branch_N_955), .B(n32548), .C(n10024), 
         .Z(n8)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_501.init = 16'hfefe;
    LUT4 i1_2_lut_adj_502 (.A(is_ret_de), .B(n34287), .Z(n28827)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_502.init = 16'h8888;
    PFUMX mux_833_i11 (.BLUT(n1742_adj_3219[10]), .ALUT(n1203[10]), .C0(n30926), 
          .Z(pc_23__N_911[10]));
    PFUMX mux_833_i10 (.BLUT(n1742_adj_3219[9]), .ALUT(n1203[9]), .C0(n30926), 
          .Z(pc_23__N_911[9]));
    LUT4 i1_4_lut_adj_503 (.A(addr[7]), .B(n32835), .C(addr[6]), .D(\addr[5] ), 
         .Z(n27178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_503.init = 16'hfffe;
    LUT4 n32025_bdd_3_lut (.A(n32025), .B(\instr[31] ), .C(n4251), .Z(n32026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n32025_bdd_3_lut.init = 16'hcaca;
    PFUMX mux_833_i9 (.BLUT(n1742_adj_3219[8]), .ALUT(n1203[8]), .C0(n30926), 
          .Z(pc_23__N_911[8]));
    PFUMX mux_833_i8 (.BLUT(n1742_adj_3219[7]), .ALUT(n1203[7]), .C0(n30925), 
          .Z(pc_23__N_911[7]));
    PFUMX mux_833_i7 (.BLUT(n1742_adj_3219[6]), .ALUT(n1203[6]), .C0(n30925), 
          .Z(pc_23__N_911[6]));
    PFUMX mux_833_i6 (.BLUT(n1742_adj_3219[5]), .ALUT(n1203[5]), .C0(n30925), 
          .Z(pc_23__N_911[5]));
    LUT4 i1_4_lut_adj_504 (.A(n28937), .B(n32609), .C(n28925), .D(n32656), 
         .Z(is_ret_de)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_504.init = 16'h0020;
    PFUMX mux_833_i5 (.BLUT(n1742_adj_3219[4]), .ALUT(n1203[4]), .C0(n30925), 
          .Z(pc_23__N_911[4]));
    LUT4 mux_1520_i10_3_lut (.A(n31[9]), .B(n33[9]), .C(n2150), .Z(n2151[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i10_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_505 (.A(n32617), .B(n29661), .C(n32655), .D(n28919), 
         .Z(n28937)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_505.init = 16'h0200;
    LUT4 n3340_bdd_3_lut_29021_4_lut (.A(\instr[31] ), .B(n32630), .C(n32539), 
         .D(n32019), .Z(n32020)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3340_bdd_3_lut_29021_4_lut.init = 16'hf808;
    LUT4 i1_4_lut_adj_506 (.A(n32640), .B(n32661), .C(n32639), .D(n32638), 
         .Z(n28925)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_506.init = 16'h1000;
    PFUMX mux_833_i4 (.BLUT(n1742_adj_3219[3]), .ALUT(n1203[3]), .C0(n30924), 
          .Z(pc_23__N_911[3]));
    LUT4 mux_2089_i14_3_lut_4_lut (.A(\instr[31] ), .B(n32630), .C(n32539), 
         .D(n4969[6]), .Z(n3328[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2089_i14_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_3151_i28_3_lut_3_lut_4_lut (.A(\instr[31] ), .B(n32630), .C(n29747), 
         .D(n32540), .Z(n5205[27])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3151_i28_3_lut_3_lut_4_lut.init = 16'hf088;
    PFUMX mux_833_i3 (.BLUT(n1742_adj_3219[2]), .ALUT(n1203[2]), .C0(n30924), 
          .Z(pc_23__N_911[2]));
    LUT4 i1_4_lut_4_lut_4_lut_adj_507 (.A(n32548), .B(n32543), .C(n28797), 
         .D(n32546), .Z(n27509)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_507.init = 16'h0040;
    LUT4 mux_2089_i15_3_lut_4_lut (.A(\instr[31] ), .B(n32630), .C(n32539), 
         .D(n4969[7]), .Z(n3328[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2089_i15_3_lut_4_lut.init = 16'hf808;
    PFUMX mux_833_i2 (.BLUT(n1742_adj_3219[1]), .ALUT(n1203[1]), .C0(n30924), 
          .Z(pc_23__N_911[1]));
    LUT4 mux_2089_i13_3_lut_4_lut (.A(\instr[31] ), .B(n32630), .C(n32539), 
         .D(n4969[5]), .Z(n3328[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2089_i13_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_1539_i9_3_lut (.A(n33[8]), .B(n34[8]), .C(n2130), .Z(n2202[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i9_3_lut.init = 16'hcaca;
    LUT4 n3508_bdd_3_lut_29029 (.A(n3493[17]), .B(n32028), .C(n32525), 
         .Z(n32029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3508_bdd_3_lut_29029.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_4_lut_adj_508 (.A(n32548), .B(n32543), .C(n28733), 
         .D(n32546), .Z(n2557)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_508.init = 16'h0040;
    LUT4 mux_1543_i9_3_lut (.A(n36[8]), .B(n31[8]), .C(n2150), .Z(n2222[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i9_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_4_lut_adj_509 (.A(n32548), .B(n32543), .C(n28647), 
         .D(n32546), .Z(n27483)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_509.init = 16'h0040;
    LUT4 n4263_bdd_3_lut (.A(n4251), .B(\instr[31] ), .C(instr[19]), .Z(n32031)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n4263_bdd_3_lut.init = 16'hd8d8;
    LUT4 mux_2089_i16_3_lut_4_lut (.A(\instr[31] ), .B(n32630), .C(n32539), 
         .D(n4969[8]), .Z(n3328[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2089_i16_3_lut_4_lut.init = 16'hf808;
    PFUMX mux_833_i1 (.BLUT(n1742_adj_3219[0]), .ALUT(n1203[0]), .C0(n30924), 
          .Z(pc_23__N_911[0]));
    LUT4 mux_1539_i13_3_lut (.A(n33[12]), .B(n34[12]), .C(n2130), .Z(n2202[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1543_i13_3_lut (.A(n36[12]), .B(n31[12]), .C(n2150), .Z(n2222[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i13_3_lut.init = 16'hcaca;
    LUT4 n4251_bdd_4_lut_29496 (.A(n32630), .B(n29714), .C(n29702), .D(n32734), 
         .Z(n32051)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n4251_bdd_4_lut_29496.init = 16'h88a0;
    LUT4 n32049_bdd_3_lut (.A(n32049), .B(n32643), .C(n4251), .Z(n32050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n32049_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_510 (.A(n32689), .B(n32537), .C(data_txn_len[1]), 
         .D(instr_active), .Z(txn_len[1])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(435[34:115])
    defparam i1_3_lut_4_lut_adj_510.init = 16'h00b0;
    LUT4 n3508_bdd_3_lut (.A(n3493[17]), .B(n32033), .C(n32525), .Z(n32034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3508_bdd_3_lut.init = 16'hcaca;
    LUT4 n3340_bdd_3_lut_29030_4_lut (.A(\instr[31] ), .B(n32630), .C(n32539), 
         .D(n32031), .Z(n32032)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3340_bdd_3_lut_29030_4_lut.init = 16'hf808;
    LUT4 mux_1516_i10_3_lut (.A(n34[9]), .B(n36[9]), .C(n2130), .Z(n2131[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i10_3_lut.init = 16'hcaca;
    LUT4 mux_2135_i32_3_lut_4_lut (.A(\instr[31] ), .B(n32630), .C(n32525), 
         .D(n3493[17]), .Z(n3446[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2135_i32_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_1543_i10_3_lut (.A(n36[9]), .B(n31[9]), .C(n2150), .Z(n2222[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i10_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_511 (.A(n32543), .B(n32546), .C(n32548), .D(n28575), 
         .Z(n10772)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_511.init = 16'h0200;
    LUT4 i8958_2_lut_rep_632_3_lut_4_lut (.A(alu_op[0]), .B(n32732), .C(data_rs1[3]), 
         .D(n32733), .Z(n32647)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i8958_2_lut_rep_632_3_lut_4_lut.init = 16'hf040;
    LUT4 i1_2_lut_adj_512 (.A(n26), .B(n10772), .Z(n4257)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_512.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_513 (.A(alu_op[0]), .B(n32732), .C(data_rs1[2]), 
         .D(n32733), .Z(n21665)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_3_lut_4_lut_adj_513.init = 16'hf040;
    LUT4 i1_3_lut_4_lut_adj_514 (.A(n32765), .B(rst_reg_n_adj_6), .C(data_ready_latch), 
         .D(address_ready), .Z(clk_c_enable_325)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_514.init = 16'hff7f;
    LUT4 mux_1520_i9_3_lut (.A(n31[8]), .B(n33[8]), .C(n2150), .Z(n2151[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i9_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_515 (.A(n32765), .B(rst_reg_n_adj_6), .C(data_ready_latch), 
         .D(n32575), .Z(n27854)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_515.init = 16'h0800;
    LUT4 mux_1516_i9_3_lut (.A(n34[8]), .B(n36[8]), .C(n2130), .Z(n2131[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_516 (.A(qspi_data_ready), .B(n32742), .C(instr_fetch_running), 
         .D(n32824), .Z(n28475)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_2_lut_4_lut_adj_516.init = 16'h8000;
    LUT4 mux_1520_i4_3_lut (.A(n31[3]), .B(n33[3]), .C(n2150), .Z(n2151[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1516_i4_3_lut (.A(n34[3]), .B(n36[3]), .C(n2130), .Z(n2131[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i4_3_lut.init = 16'hcaca;
    LUT4 mux_2089_i12_3_lut_4_lut (.A(n32540), .B(n32539), .C(n4969[4]), 
         .D(n29700), .Z(n3328[11])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2089_i12_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_1539_i16_3_lut (.A(n33[15]), .B(n34[15]), .C(n2130), .Z(n2202[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i16_3_lut.init = 16'hcaca;
    LUT4 i4629_2_lut_rep_667_4_lut (.A(qspi_data_ready), .B(n32742), .C(instr_fetch_running), 
         .D(\instr_addr_23__N_318[0] ), .Z(n32682)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i4629_2_lut_rep_667_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_517 (.A(qspi_data_ready), .B(n32742), .C(instr_fetch_running), 
         .D(n32798), .Z(n28699)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_2_lut_4_lut_adj_517.init = 16'hff7f;
    LUT4 mux_2107_i1_4_lut (.A(n28413), .B(n10024), .C(n4267), .D(n28585), 
         .Z(n29685)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2107_i1_4_lut.init = 16'h3a0a;
    LUT4 mux_1543_i16_3_lut (.A(n36[15]), .B(n31[15]), .C(n2150), .Z(n2222[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i16_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_518 (.A(qspi_data_ready), .B(n32742), .C(instr_fetch_running), 
         .D(n32797), .Z(n28705)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_2_lut_4_lut_adj_518.init = 16'hff7f;
    LUT4 i1_2_lut_4_lut_adj_519 (.A(qspi_data_ready), .B(n32742), .C(instr_fetch_running), 
         .D(n32796), .Z(n28719)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_2_lut_4_lut_adj_519.init = 16'hff7f;
    LUT4 i1_4_lut_4_lut_4_lut_adj_520 (.A(n32548), .B(n32543), .C(n28553), 
         .D(n32546), .Z(n27364)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_520.init = 16'h0040;
    LUT4 mux_2111_i21_3_lut_4_lut (.A(n32525), .B(n32540), .C(n3446[24]), 
         .D(n29700), .Z(n3446[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2111_i21_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_4_lut_4_lut_4_lut_adj_521 (.A(n32548), .B(n32543), .C(n28611), 
         .D(n32546), .Z(n27492)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_521.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_522 (.A(n32548), .B(n32543), .C(n28567), 
         .D(n32546), .Z(n27356)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_522.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_523 (.A(n32548), .B(n32543), .C(n28599), 
         .D(n32546), .Z(n27495)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_523.init = 16'h0040;
    LUT4 i1_2_lut_adj_524 (.A(n16_c), .B(n10772), .Z(n4267)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_524.init = 16'h8888;
    LUT4 i1_4_lut_adj_525 (.A(n32655), .B(n10772), .C(n32489), .D(n28), 
         .Z(n4271)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_525.init = 16'hc8c0;
    LUT4 i28368_4_lut (.A(n32552), .B(n32544), .C(n32707), .D(n28755), 
         .Z(clk_c_enable_232)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i28368_4_lut.init = 16'h0010;
    LUT4 i28343_4_lut (.A(n32552), .B(rst_reg_n_adj_6), .C(n32544), .D(n28699), 
         .Z(clk_c_enable_234)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i28343_4_lut.init = 16'h3337;
    LUT4 mux_1539_i8_3_lut (.A(n33[7]), .B(\instr_data[1][7] ), .C(n2130), 
         .Z(n2211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i8_3_lut.init = 16'hcaca;
    LUT4 i3063_4_lut_4_lut_4_lut (.A(n32548), .B(n32543), .C(n28577), 
         .D(n32546), .Z(n2577[1])) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i3063_4_lut_4_lut_4_lut.init = 16'hffbf;
    LUT4 mux_1520_i5_rep_93_3_lut (.A(n31[4]), .B(n33[4]), .C(n2150), 
         .Z(n29712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i5_rep_93_3_lut.init = 16'hcaca;
    LUT4 mux_1516_i5_rep_81_3_lut (.A(n34[4]), .B(n36[4]), .C(n2130), 
         .Z(n29700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i5_rep_81_3_lut.init = 16'hcaca;
    L6MUX21 shift_right_317_i272 (.D0(n29759), .D1(n11061), .SD(n30160), 
            .Z(debug_branch_N_840[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i28348_4_lut (.A(n32552), .B(n32544), .C(n32707), .D(n28747), 
         .Z(clk_c_enable_248)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i28348_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_4_lut_4_lut_adj_526 (.A(n32548), .B(n32543), .C(n28837), 
         .D(n32546), .Z(n27567)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_526.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_527 (.A(n32548), .B(rst_reg_n_adj_6), .C(n17949), 
         .D(n10024), .Z(n28429)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_527.init = 16'h0004;
    LUT4 i1_4_lut_4_lut_adj_528 (.A(n32548), .B(n28435), .C(n17949), .D(n10024), 
         .Z(n28441)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_528.init = 16'h0004;
    LUT4 i28340_4_lut (.A(n32552), .B(rst_reg_n_adj_6), .C(n32544), .D(n28705), 
         .Z(clk_c_enable_250)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i28340_4_lut.init = 16'h3337;
    LUT4 i1_4_lut_4_lut_4_lut_adj_529 (.A(n32548), .B(n32543), .C(n28635), 
         .D(n32546), .Z(n27486)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_529.init = 16'h0040;
    LUT4 mux_1520_i6_rep_95_3_lut (.A(n31[5]), .B(n33[5]), .C(n2150), 
         .Z(n29714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i6_rep_95_3_lut.init = 16'hcaca;
    LUT4 mux_1516_i6_rep_83_3_lut (.A(n34[5]), .B(n36[5]), .C(n2130), 
         .Z(n29702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i6_rep_83_3_lut.init = 16'hcaca;
    PFUMX i29_adj_530 (.BLUT(n29758), .ALUT(n29760), .C0(n32735), .Z(n11061));
    LUT4 mux_1520_i7_rep_97_3_lut (.A(n31[6]), .B(n33[6]), .C(n2150), 
         .Z(n29716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i7_rep_97_3_lut.init = 16'hcaca;
    LUT4 mux_1516_i7_rep_91_3_lut (.A(n34[6]), .B(n36[6]), .C(n2130), 
         .Z(n29710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i7_rep_91_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_531 (.A(n32654), .B(n24), .C(n32653), .D(n10772), 
         .Z(n1_adj_3208)) /* synthesis lut_function=(A (C (D))+!A !((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i1_2_lut_4_lut_adj_531.init = 16'ha400;
    LUT4 mux_2089_i17_3_lut_4_lut (.A(n32539), .B(n32568), .C(n4969[9]), 
         .D(n29741), .Z(n3328[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2089_i17_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_1520_i8_rep_99_3_lut (.A(\instr_data[3][7] ), .B(n33[7]), .C(n2150), 
         .Z(n29718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i8_rep_99_3_lut.init = 16'hcaca;
    LUT4 i28334_4_lut (.A(n32552), .B(n32544), .C(n32707), .D(n28739), 
         .Z(clk_c_enable_292)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i28334_4_lut.init = 16'h0010;
    LUT4 mux_1520_i11_3_lut (.A(n31[10]), .B(n33[10]), .C(n2150), .Z(n2151[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1516_i11_rep_108_3_lut (.A(n34[10]), .B(n36[10]), .C(n2130), 
         .Z(n29727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i11_rep_108_3_lut.init = 16'hcaca;
    LUT4 debug_branch_I_48_i4_3_lut (.A(debug_branch_N_840[31]), .B(timer_data[3]), 
         .C(is_timer_addr), .Z(debug_branch_N_450[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_48_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_4_lut_adj_532 (.A(n32548), .B(n32543), .C(n28673), 
         .D(n32546), .Z(n3369[11])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_532.init = 16'h0040;
    LUT4 mux_1539_i12_3_lut (.A(n33[11]), .B(n34[11]), .C(n2130), .Z(n2202[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1539_i12_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_533 (.A(n29), .B(\uart_rx_buf_data[7] ), .C(\baud_divider[7] ), 
         .D(addr[3]), .Z(n2)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_533.init = 16'ha088;
    PFUMX i27135 (.BLUT(n29843), .ALUT(n227), .C0(counter_hi[4]), .Z(n29844));
    LUT4 mux_1543_i12_3_lut (.A(n36[11]), .B(n31[11]), .C(n2150), .Z(n2222[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1543_i12_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_4_lut_adj_534 (.A(n32548), .B(n28413), .C(n32552), 
         .D(n32545), .Z(n28417)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_534.init = 16'h4440;
    LUT4 additional_mem_ops_2__N_1132_0__bdd_3_lut_29242 (.A(additional_mem_ops_2__N_1132[0]), 
         .B(n32656), .C(n32653), .Z(n32179)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam additional_mem_ops_2__N_1132_0__bdd_3_lut_29242.init = 16'h8080;
    LUT4 i28591_3_lut (.A(n32540), .B(n32533), .C(n32734), .Z(n30084)) /* synthesis lut_function=(A+!((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28591_3_lut.init = 16'haeae;
    L6MUX21 i27613 (.D0(n30320), .D1(n30321), .SD(counter_hi[3]), .Z(n30322));
    LUT4 i1_4_lut_adj_535 (.A(n22), .B(n10024), .C(n4_c), .D(n32571), 
         .Z(n28837)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_535.init = 16'h0200;
    LUT4 i1_4_lut_adj_536 (.A(n32614), .B(n32619), .C(n32613), .D(n32653), 
         .Z(n4_c)) /* synthesis lut_function=(!((B (C (D))+!B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_536.init = 16'h0a88;
    LUT4 mux_1526_i3_3_lut (.A(n29743), .B(n2151[2]), .C(n32734), .Z(instr[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i3_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_537 (.A(clk_c_enable_365), .B(n32630), .C(n32617), 
         .D(n32612), .Z(n2798)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_537.init = 16'ha888;
    LUT4 mux_1516_i3_rep_124_3_lut (.A(n34[2]), .B(n36[2]), .C(n2130), 
         .Z(n29743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i3_rep_124_3_lut.init = 16'hcaca;
    LUT4 mux_1520_i3_3_lut (.A(n31[2]), .B(n33[2]), .C(n2150), .Z(n2151[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i3_3_lut.init = 16'hcaca;
    PFUMX i48 (.BLUT(n12_adj_3192), .ALUT(n30_adj_3211), .C0(n30919), 
          .Z(n43));
    LUT4 i1_4_lut_adj_538 (.A(clk_c_enable_365), .B(n32630), .C(n20_adj_3181), 
         .D(n25), .Z(n2800)) /* synthesis lut_function=(A (B+!(C+(D)))) */ ;
    defparam i1_4_lut_adj_538.init = 16'h888a;
    LUT4 i1_2_lut_adj_539 (.A(mie[2]), .B(\next_fsm_state_3__N_3046[3] ), 
         .Z(n76)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(71[11:25])
    defparam i1_2_lut_adj_539.init = 16'h8888;
    LUT4 is_alu_imm_N_1367_bdd_3_lut_29261_4_lut (.A(n32642), .B(n32605), 
         .C(n32655), .D(n32639), .Z(n32268)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam is_alu_imm_N_1367_bdd_3_lut_29261_4_lut.init = 16'h0800;
    LUT4 i1_4_lut_adj_540 (.A(n32639), .B(n32642), .C(n32570), .D(n29681), 
         .Z(n26863)) /* synthesis lut_function=(!((B (C+(D))+!B !((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_540.init = 16'h220a;
    LUT4 i2_2_lut (.A(n22), .B(n10772), .Z(n2796)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_4_lut_4_lut_adj_541 (.A(n32548), .B(n32543), .C(n28659), 
         .D(n32546), .Z(n27480)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_541.init = 16'h0040;
    L6MUX21 i29736 (.D0(n33739), .D1(n33736), .SD(n2126), .Z(n33740));
    LUT4 mux_1526_i2_3_lut (.A(n29745), .B(n2151[1]), .C(n32734), .Z(instr[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i2_3_lut.init = 16'hcaca;
    PFUMX i29734 (.BLUT(n33738), .ALUT(n33737), .C0(n2122), .Z(n33739));
    LUT4 mux_1516_i2_rep_126_3_lut (.A(n34[1]), .B(n36[1]), .C(n2130), 
         .Z(n29745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i2_rep_126_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_4_lut_adj_542 (.A(n32548), .B(n32543), .C(n28285), 
         .D(n32546), .Z(n4243)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_542.init = 16'h0040;
    LUT4 mux_1520_i2_3_lut (.A(n31[1]), .B(n33[1]), .C(n2150), .Z(n2151[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i2_3_lut.init = 16'hcaca;
    L6MUX21 i27611 (.D0(n30316), .D1(n30317), .SD(counter_hi[2]), .Z(n30320));
    L6MUX21 i27612 (.D0(n30318), .D1(n30319), .SD(counter_hi[2]), .Z(n30321));
    LUT4 i15309_2_lut_3_lut_4_lut (.A(n32836), .B(n32835), .C(\ui_in_sync[5] ), 
         .D(n32818), .Z(data_from_user_peri_1__31__N_2455[5])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i15309_2_lut_3_lut_4_lut.init = 16'h0010;
    FD1S3IX counter_hi_3544__i4_rep_844 (.D(n39[2]), .CK(clk_c), .CD(n32840), 
            .Q(n34281));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3544__i4_rep_844.GSR = "DISABLED";
    L6MUX21 i27618 (.D0(n30323), .D1(n30324), .SD(counter_hi[2]), .Z(n30327));
    LUT4 i1_2_lut_3_lut_4_lut_adj_543 (.A(n32836), .B(n32835), .C(\ui_in_sync[6] ), 
         .D(n32818), .Z(n19_adj_3193)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_4_lut_adj_543.init = 16'h0010;
    LUT4 i1_4_lut_adj_544 (.A(n21414), .B(addr[10]), .C(addr[6]), .D(data_ready_r), 
         .Z(n29485)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_544.init = 16'hfffe;
    PFUMX i29731 (.BLUT(n33735), .ALUT(n32072), .C0(n2124), .Z(n33736));
    LUT4 i1_2_lut_rep_679_4_lut (.A(n32835), .B(n32762), .C(addr[6]), 
         .D(addr[7]), .Z(n32694)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_679_4_lut.init = 16'hfffe;
    LUT4 data_from_read_2__bdd_4_lut (.A(n32598), .B(data_txn_len[0]), .C(instr_data[10]), 
         .D(instr_data[2]), .Z(n32992)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam data_from_read_2__bdd_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_adj_545 (.A(n19_c), .B(n10772), .Z(n4259)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_545.init = 16'h8888;
    PFUMX i29307 (.BLUT(n32858), .ALUT(n32859), .C0(counter_hi[2]), .Z(n32860));
    LUT4 i11800_4_lut (.A(n32632), .B(n32637), .C(n32639), .D(n32602), 
         .Z(n7_adj_3212)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(47[17:22])
    defparam i11800_4_lut.init = 16'h0a3a;
    LUT4 i1_4_lut_adj_546 (.A(n32819), .B(n29614), .C(qv_data_write_n[1]), 
         .D(addr[10]), .Z(n29549)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_546.init = 16'h0100;
    L6MUX21 i27714 (.D0(n30419), .D1(n30420), .SD(counter_hi[2]), .Z(n30423));
    LUT4 i26972_2_lut (.A(\addr[4] ), .B(qv_data_write_n[0]), .Z(n29614)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26972_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_4_lut_4_lut_adj_547 (.A(n32548), .B(n32543), .C(n28811), 
         .D(n32546), .Z(n27502)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_547.init = 16'h0040;
    LUT4 i28609_2_lut (.A(n32525), .B(n4271), .Z(n30032)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28609_2_lut.init = 16'hbbbb;
    PFUMX i28802 (.BLUT(n31651), .ALUT(n31650), .C0(counter_hi[2]), .Z(n31652));
    PFUMX next_pc_for_core_23__I_0_i209 (.BLUT(n149), .ALUT(n225), .C0(counter_hi[4]), 
          .Z(n209)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i28271_4_lut (.A(n32552), .B(rst_reg_n_adj_6), .C(n32544), .D(n28719), 
         .Z(clk_c_enable_294)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i28271_4_lut.init = 16'h3337;
    PFUMX i38 (.BLUT(n17), .ALUT(n22_adj_3213), .C0(n32639), .Z(n24_adj_3199));
    LUT4 mux_2084_i11_4_lut (.A(n32643), .B(n32584), .C(n4267), .D(n32656), 
         .Z(n3259[10])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2084_i11_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_4_lut_4_lut_adj_548 (.A(n32548), .B(n32543), .C(n28783), 
         .D(n32546), .Z(n27516)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_548.init = 16'h0040;
    LUT4 n10904_bdd_4_lut_29273 (.A(n32577), .B(n32638), .C(n32654), .D(additional_mem_ops_2__N_1132[0]), 
         .Z(n32189)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam n10904_bdd_4_lut_29273.init = 16'hf808;
    LUT4 i1_3_lut_adj_549 (.A(n35), .B(n26), .C(n28669), .Z(n28673)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_549.init = 16'h8080;
    LUT4 i1_4_lut_adj_550 (.A(n32552), .B(n32544), .C(n32707), .D(n28821), 
         .Z(clk_c_enable_308)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(410[18] 430[16])
    defparam i1_4_lut_adj_550.init = 16'h1000;
    PFUMX i27749 (.BLUT(n30454), .ALUT(n30455), .C0(counter_hi[3]), .Z(n30458));
    LUT4 i15308_2_lut_3_lut_4_lut (.A(n32836), .B(n32835), .C(\ui_in_sync[7] ), 
         .D(n32818), .Z(\data_from_user_peri_1__31__N_2455[7] )) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i15308_2_lut_3_lut_4_lut.init = 16'h0010;
    PFUMX i27129 (.BLUT(n29837), .ALUT(n226), .C0(counter_hi[4]), .Z(n29838));
    PFUMX i27750 (.BLUT(n30456), .ALUT(n30457), .C0(counter_hi[3]), .Z(n30459));
    LUT4 i1_4_lut_adj_551 (.A(n2_c), .B(next_instr_write_offset[3]), .C(n1_c), 
         .D(n28511), .Z(n19867)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_551.init = 16'h0400;
    LUT4 i15544_2_lut_rep_569_3_lut (.A(n32653), .B(n32656), .C(n32642), 
         .Z(n32584)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15544_2_lut_rep_569_3_lut.init = 16'h4040;
    LUT4 i1_4_lut_adj_552 (.A(\uart_rx_buf_data[6] ), .B(n26856), .C(\baud_divider[6] ), 
         .D(addr[3]), .Z(n26858)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_4_lut_adj_552.init = 16'hc088;
    LUT4 mux_1526_i15_3_lut (.A(n29733), .B(n2151[14]), .C(n32734), .Z(instr[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1526_i15_3_lut.init = 16'hcaca;
    PFUMX i27756 (.BLUT(n30461), .ALUT(n30462), .C0(counter_hi[3]), .Z(n30465));
    LUT4 i1_4_lut_adj_553 (.A(\uart_rx_buf_data[5] ), .B(n26856), .C(\baud_divider[5] ), 
         .D(addr[3]), .Z(n26857)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_4_lut_adj_553.init = 16'hc088;
    LUT4 mux_1516_i15_rep_114_3_lut (.A(n34[14]), .B(n36[14]), .C(n2130), 
         .Z(n29733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i15_rep_114_3_lut.init = 16'hcaca;
    LUT4 mux_1520_i15_3_lut (.A(n31[14]), .B(n33[14]), .C(n2150), .Z(n2151[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i15_3_lut.init = 16'hcaca;
    LUT4 n8539_bdd_4_lut (.A(n32560), .B(n32601), .C(n32618), .D(n32654), 
         .Z(n32224)) /* synthesis lut_function=(!(A (B (C))+!A !(((D)+!C)+!B))) */ ;
    defparam n8539_bdd_4_lut.init = 16'h7f3f;
    PFUMX i27608 (.BLUT(\mem_data_from_read[4] ), .ALUT(\data_from_read[4] ), 
          .C0(n30930), .Z(n30317));
    LUT4 n32224_bdd_3_lut (.A(n32224), .B(n32223), .C(n30920), .Z(n32225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n32224_bdd_3_lut.init = 16'hcaca;
    PFUMX i27757 (.BLUT(n30463), .ALUT(n30464), .C0(counter_hi[3]), .Z(n30466));
    LUT4 i15677_2_lut_rep_678_4_lut (.A(addr[6]), .B(n32762), .C(addr[7]), 
         .D(n32728), .Z(n32693)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i15677_2_lut_rep_678_4_lut.init = 16'hfffd;
    LUT4 additional_mem_ops_1__bdd_2_lut_29432 (.A(additional_mem_ops[1]), 
         .B(additional_mem_ops[0]), .Z(n32226)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam additional_mem_ops_1__bdd_2_lut_29432.init = 16'h1111;
    PFUMX i27609 (.BLUT(\mem_data_from_read[8] ), .ALUT(\data_from_read[8] ), 
          .C0(n30929), .Z(n30318));
    LUT4 mux_3119_i12_3_lut (.A(n32642), .B(n32658), .C(n32656), .Z(n5138[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3119_i12_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_then_4_lut (.A(n8_c), .B(n2222[3]), .C(n28501), .D(n32658), 
         .Z(n32876)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h4010;
    LUT4 mux_3119_i13_3_lut (.A(n32642), .B(n32657), .C(n32656), .Z(n5138[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3119_i13_3_lut.init = 16'hcaca;
    LUT4 mux_3119_i14_3_lut (.A(n32642), .B(n32661), .C(n32656), .Z(n5138[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3119_i14_3_lut.init = 16'hcaca;
    PFUMX i27610 (.BLUT(\mem_data_from_read[12] ), .ALUT(\data_from_read[12] ), 
          .C0(n30929), .Z(n30319));
    PFUMX i27614 (.BLUT(\mem_data_from_read[1] ), .ALUT(\data_from_read[1] ), 
          .C0(n30929), .Z(n30323));
    LUT4 i6612_3_lut_4_lut (.A(n32630), .B(n32734), .C(n29748), .D(n2131[11]), 
         .Z(n3328[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i6612_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_3119_i15_3_lut (.A(n32642), .B(n32659), .C(n32656), .Z(n5138[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3119_i15_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_554 (.A(mie[14]), .B(n21665), .C(n8_adj_3200), .Z(n926)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_554.init = 16'hcece;
    LUT4 data_from_user_peri_1__31__N_2455_0__bdd_4_lut (.A(\data_from_user_peri_1__31__N_2455[0] ), 
         .B(n32720), .C(addr[6]), .D(\uo_out_from_user_peri[1][0] ), .Z(n32254)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(B+!(C (D)))) */ ;
    defparam data_from_user_peri_1__31__N_2455_0__bdd_4_lut.init = 16'hb080;
    PFUMX i27615 (.BLUT(\mem_data_from_read[5] ), .ALUT(\data_from_read[5] ), 
          .C0(n30929), .Z(n30324));
    LUT4 i1_4_lut_adj_555 (.A(n6920), .B(n28237), .C(\instr_write_offset[3] ), 
         .D(instr_complete_N_1647), .Z(next_instr_write_offset[3])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i1_4_lut_adj_555.init = 16'h965a;
    LUT4 i26959_4_lut_4_lut_4_lut (.A(n32548), .B(n32543), .C(n29685), 
         .D(n32546), .Z(n29600)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i26959_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_556 (.A(n32548), .B(n32607), .C(n17949), .D(n10024), 
         .Z(n28465)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_556.init = 16'h0004;
    LUT4 i1_4_lut_4_lut_4_lut_adj_557 (.A(n32548), .B(n32543), .C(n28769), 
         .D(n32546), .Z(n27523)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_557.init = 16'h0040;
    LUT4 n32360_bdd_2_lut_3_lut_3_lut_4_lut (.A(n32656), .B(n32655), .C(n32360), 
         .D(n32630), .Z(n32361)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;
    defparam n32360_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'hf010;
    LUT4 i1_4_lut_4_lut_adj_558 (.A(n32548), .B(n28269), .C(n17949), .D(n10024), 
         .Z(n28275)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_558.init = 16'h0004;
    LUT4 i15541_2_lut_3_lut (.A(n32653), .B(n32656), .C(n32657), .Z(n3292[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15541_2_lut_3_lut.init = 16'h4040;
    LUT4 mux_2084_i12_4_lut_4_lut_4_lut (.A(n32653), .B(n32656), .C(n4267), 
         .D(n32642), .Z(n3259[11])) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (C (D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2084_i12_4_lut_4_lut_4_lut.init = 16'h4300;
    LUT4 i1_4_lut_4_lut_adj_559 (.A(n32548), .B(n34287), .C(n32655), .D(n10024), 
         .Z(n28483)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_559.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_560 (.A(n32548), .B(n28447), .C(n17949), .D(n10024), 
         .Z(n28453)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_560.init = 16'h0004;
    LUT4 i28569_2_lut (.A(n34281), .B(n34283), .Z(n30179)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i28569_2_lut.init = 16'heeee;
    PFUMX i29290 (.BLUT(n32494), .ALUT(n32493), .C0(n32639), .Z(n22));
    LUT4 i1_4_lut_adj_561 (.A(no_write_in_progress), .B(data_ready_core), 
         .C(debug_instr_valid), .D(is_load), .Z(debug_rd_3__N_1575)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_4_lut_adj_561.init = 16'h8000;
    PFUMX i28782 (.BLUT(n31626), .ALUT(n31625), .C0(counter_hi[2]), .Z(n31627));
    LUT4 i1_3_lut_rep_691_4_lut (.A(n32771), .B(n21414), .C(data_out_hold), 
         .D(n12), .Z(n32706)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_3_lut_rep_691_4_lut.init = 16'h0200;
    LUT4 i1_3_lut_rep_566_4_lut (.A(n32656), .B(n32655), .C(n32654), .D(n32639), 
         .Z(n32581)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_3_lut_rep_566_4_lut.init = 16'hefff;
    LUT4 i1_2_lut_3_lut_4_lut_adj_562 (.A(n32656), .B(n32655), .C(n32605), 
         .D(n32642), .Z(n19_adj_3214)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_562.init = 16'h1101;
    LUT4 i1_4_lut_adj_563 (.A(was_early_branch), .B(n10253), .C(n16_adj_3168), 
         .D(n32630), .Z(n10024)) /* synthesis lut_function=(A+(B (C (D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[82:120])
    defparam i1_4_lut_adj_563.init = 16'hfaba;
    PFUMX i27710 (.BLUT(\mem_data_from_read[3] ), .ALUT(\data_from_read[3] ), 
          .C0(n30930), .Z(n30419));
    LUT4 i1_4_lut_4_lut_4_lut_adj_564 (.A(n32548), .B(n32543), .C(n28623), 
         .D(n32546), .Z(n27489)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_564.init = 16'h0040;
    PFUMX i29286 (.BLUT(n32488), .ALUT(n32487), .C0(n30919), .Z(n32489));
    PFUMX i29535 (.BLUT(n33404), .ALUT(n33403), .C0(n32548), .Z(additional_mem_ops_2__N_749[1]));
    LUT4 mux_1520_i12_3_lut (.A(n31[11]), .B(n33[11]), .C(n2150), .Z(n2151[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1520_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1516_i12_3_lut (.A(n34[11]), .B(n36[11]), .C(n2130), .Z(n2131[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i12_3_lut.init = 16'hcaca;
    PFUMX i27711 (.BLUT(\mem_data_from_read[7] ), .ALUT(\data_from_read[7] ), 
          .C0(n32771), .Z(n30420));
    PFUMX i28778 (.BLUT(n31621), .ALUT(n31620), .C0(counter_hi[2]), .Z(n31622));
    LUT4 i1_3_lut_rep_532 (.A(address_ready), .B(n32549), .C(is_load), 
         .Z(n32547)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(291[13:39])
    defparam i1_3_lut_rep_532.init = 16'h2020;
    LUT4 i1_4_lut_adj_565 (.A(n29), .B(\uart_rx_buf_data[3] ), .C(\baud_divider[3] ), 
         .D(addr[3]), .Z(n2_adj_9)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_565.init = 16'ha088;
    PFUMX i27607 (.BLUT(\mem_data_from_read[0] ), .ALUT(\data_from_read[0] ), 
          .C0(n30930), .Z(n30316));
    LUT4 i28356_3_lut_4_lut (.A(n4271), .B(n16_c), .C(n10772), .D(n19_c), 
         .Z(n30007)) /* synthesis lut_function=(!(A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i28356_3_lut_4_lut.init = 16'h5f7f;
    LUT4 i2_4_lut_rep_510 (.A(n32630), .B(clk_c_enable_365), .C(n32617), 
         .D(n32619), .Z(n32525)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;
    defparam i2_4_lut_rep_510.init = 16'hc888;
    PFUMX i32_adj_566 (.BLUT(n27896), .ALUT(n17_adj_3197), .C0(n32654), 
          .Z(n19_c));
    LUT4 i1_3_lut_rep_692_4_lut (.A(n32787), .B(instr_active), .C(instr_fetch_running), 
         .D(qspi_data_ready), .Z(n32707)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_3_lut_rep_692_4_lut.init = 16'h8000;
    LUT4 mux_1516_i1_rep_122_3_lut (.A(\instr_data[1][0] ), .B(\instr_data[2][0] ), 
         .C(n2130), .Z(n29741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1516_i1_rep_122_3_lut.init = 16'hcaca;
    PFUMX i54 (.BLUT(n37), .ALUT(n32), .C0(n30132), .Z(n35));
    LUT4 i1_2_lut_rep_580_3_lut (.A(n32641), .B(n32637), .C(n32642), .Z(n32595)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_580_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_567 (.A(n32605), .B(n32604), .C(n32580), .D(n32642), 
         .Z(n27959)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_567.init = 16'h5fdd;
    LUT4 i15099_2_lut_3_lut_4_lut (.A(n32641), .B(n32637), .C(n32654), 
         .D(n32642), .Z(n17747)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15099_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_568 (.A(n32641), .B(n32637), .C(n26937), .Z(alu_op_3__N_1337[2])) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_568.init = 16'hf7f7;
    LUT4 i1_3_lut_adj_569 (.A(mie[10]), .B(n21665), .C(n8_adj_3200), .Z(n893)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_569.init = 16'hcece;
    PFUMX i42 (.BLUT(n10), .ALUT(n29_c), .C0(n32654), .Z(n23));
    LUT4 i1_2_lut_4_lut_adj_570 (.A(address_ready), .B(n32549), .C(is_load), 
         .D(n32671), .Z(clk_c_enable_52)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(291[13:39])
    defparam i1_2_lut_4_lut_adj_570.init = 16'hff20;
    LUT4 i15828_3_lut_4_lut (.A(n34281), .B(n32854), .C(mem_op[0]), .D(n32759), 
         .Z(n18098)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i15828_3_lut_4_lut.init = 16'hbfb0;
    LUT4 mux_3119_i16_3_lut (.A(n32642), .B(n32651), .C(n32656), .Z(n5138[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3119_i16_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_571 (.A(n28971), .B(n27804), .C(n32751), .D(n32842), 
         .Z(n12_c)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !((C (D)+!C !(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[82:120])
    defparam i1_4_lut_adj_571.init = 16'h8448;
    LUT4 n13_bdd_3_lut_29178 (.A(\mem_data_from_read[18] ), .B(\mem_data_from_read[22] ), 
         .C(counter_hi[2]), .Z(n32313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n13_bdd_3_lut_29178.init = 16'hcaca;
    LUT4 i1_4_lut_adj_572 (.A(n32543), .B(n10024), .C(n32561), .D(n28489), 
         .Z(n28495)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_572.init = 16'h2000;
    LUT4 n32315_bdd_3_lut (.A(n32994), .B(n30365), .C(counter_hi[3]), 
         .Z(n32316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n32315_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_581_3_lut (.A(n32641), .B(n32637), .C(n32642), .Z(n32596)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_581_3_lut.init = 16'hf7f7;
    PFUMX i27155 (.BLUT(\mem_data_from_read[26] ), .ALUT(\mem_data_from_read[30] ), 
          .C0(counter_hi[2]), .Z(n29864));
    PFUMX i27131 (.BLUT(\mem_data_from_read[24] ), .ALUT(\mem_data_from_read[28] ), 
          .C0(counter_hi[2]), .Z(n29840));
    LUT4 mux_2126_i12_3_lut_4_lut (.A(n4271), .B(n32527), .C(n3410[11]), 
         .D(n29723), .Z(n3493[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2126_i12_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i1_4_lut_adj_573 (.A(\uart_rx_buf_data[2] ), .B(n26856), .C(\baud_divider[2] ), 
         .D(addr[3]), .Z(n26859)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_4_lut_adj_573.init = 16'hc088;
    PFUMX i27050 (.BLUT(\mem_data_from_read[27] ), .ALUT(\mem_data_from_read[31] ), 
          .C0(counter_hi[2]), .Z(n29759));
    PFUMX i29332 (.BLUT(n32899), .ALUT(n32900), .C0(counter_hi[2]), .Z(n32901));
    PFUMX i29330 (.BLUT(n32896), .ALUT(n32897), .C0(counter_hi[2]), .Z(n32898));
    PFUMX i29232 (.BLUT(n32407), .ALUT(n32406), .C0(n32578), .Z(n32408));
    LUT4 i4826_3_lut_4_lut (.A(\instr_addr_23__N_318[0] ), .B(n32843), .C(n32766), 
         .D(instr_addr_23__N_318[1]), .Z(n4_adj_3203)) /* synthesis lut_function=(A ((D)+!C)+!A !(B (C+!(D))+!B !((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i4826_3_lut_4_lut.init = 16'hbf0b;
    LUT4 i1_4_lut_4_lut_adj_574 (.A(\instr_write_offset[3] ), .B(instr_addr_23__N_318[1]), 
         .C(\pc[2] ), .D(n2_adj_3202), .Z(n9)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A !(B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam i1_4_lut_4_lut_adj_574.init = 16'h4124;
    PFUMX i27149 (.BLUT(\mem_data_from_read[25] ), .ALUT(\mem_data_from_read[29] ), 
          .C0(counter_hi[2]), .Z(n29858));
    PFUMX i29322 (.BLUT(n32884), .ALUT(n32885), .C0(n32734), .Z(\instr[31] ));
    LUT4 i1_3_lut_adj_575 (.A(mie[6]), .B(n21665), .C(n8_adj_3200), .Z(n860)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_575.init = 16'hcece;
    PFUMX i29316 (.BLUT(n32875), .ALUT(n32876), .C0(n32734), .Z(n32877));
    PFUMX i28757 (.BLUT(n31589), .ALUT(n31588), .C0(n4257), .Z(n31590));
    PFUMX i29223 (.BLUT(n32394), .ALUT(n32393), .C0(n32578), .Z(n32395));
    LUT4 i1_4_lut_adj_576 (.A(n10024), .B(n17949), .C(n32656), .D(rst_reg_n_adj_6), 
         .Z(n28285)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_576.init = 16'h1000;
    tinyQV_time i_timer (.clk_c(clk_c), .n32840(n32840), .time_pulse_r(time_pulse_r), 
            .clk_c_enable_363(clk_c_enable_363), .n32717(n32717), .\data_rs2[2] (data_rs2[2]), 
            .data_out_3__N_1385(data_out_3__N_1385), .timer_data_3__N_631(timer_data_3__N_631), 
            .\data_rs2[0] (data_rs2[0]), .\mtimecmp[7] (mtimecmp[7]), .\mtimecmp[5] (mtimecmp[5]), 
            .clk_c_enable_285(clk_c_enable_285), .mtimecmp_1__N_1941(mtimecmp_1__N_1941), 
            .mtime_out({Open_111, Open_112, Open_113, mtime_out[0]}), 
            .\addr[2] (addr[2]), .timer_data({timer_data}), .timer_interrupt(timer_interrupt), 
            .mtimecmp_3__N_1935(mtimecmp_3__N_1935), .n10737(n10737), .cy(cy), 
            .n32663(n32663), .n32680(n32680), .rst_reg_n(rst_reg_n_adj_6), 
            .is_timer_addr(is_timer_addr), .n32801(n32801), .n32653(n32653), 
            .n32654(n32654), .n32588(n32588), .no_write_in_progress(no_write_in_progress), 
            .is_store(is_store), .clk_c_enable_178(clk_c_enable_178), .mstatus_mie_N_1709(mstatus_mie_N_1709), 
            .n32670(n32670), .n32675(n32675), .mstatus_mie_N_1707(mstatus_mie_N_1707), 
            .n32765(n32765), .clk_c_enable_207(clk_c_enable_207), .n34287(n34287), 
            .n32758(n32758), .n32746(n32746), .n32759(n32759), .clk_c_enable_433(clk_c_enable_433), 
            .\instr_addr_23__N_318[1] (instr_addr_23__N_318[1]), .\instr_addr_23__N_318[0] (\instr_addr_23__N_318[0] ), 
            .n28739(n28739), .n32691(n32691), .n29317(n29317), .n32548(n32548), 
            .n32541(n32541), .clk_c_enable_338(clk_c_enable_338), .\reg_access[4][3] (\reg_access[4] [3]), 
            .clk_c_enable_182(clk_c_enable_182), .n32760(n32760), .clk_c_enable_191(clk_c_enable_191), 
            .address_ready(address_ready), .n32671(n32671), .n28747(n28747), 
            .\instr_data[1] (instr_data[1]), .\instr_data_0__15__N_638[49] (instr_data_0__15__N_638[49]), 
            .\reg_access[3][2] (\reg_access[3] [2]), .clk_c_enable_200(clk_c_enable_200), 
            .n28755(n28755), .\instr_data[0] (instr_data[0]), .\instr_data_0__15__N_638[0] (instr_data_0__15__N_638[0]), 
            .\cycle_count_wide[3] (cycle_count_wide[3]), .n32652(n32652), 
            .clk_c_enable_276(clk_c_enable_276), .clk_c_enable_204(clk_c_enable_204), 
            .n32611(n32611), .n10024(n10024), .n32630(n32630), .n28391(n28391), 
            .n32697(n32697), .is_double_fault_r(is_double_fault_r), .mstatus_mte(mstatus_mte), 
            .n32650(n32650), .clk_c_enable_99(clk_c_enable_99), .clk_c_enable_174(clk_c_enable_174), 
            .n32668(n32668), .n32664(n32664), .\data_out_slice[0] (data_out_slice[0]), 
            .n32644(n32644), .\data_out_slice[2] (data_out_slice[2])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(450[17] 461[6])
    tinyqv_decoder i_decoder (.n32361(n32361), .n32623(n32623), .n32362(n32362), 
            .is_jal_N_1374(is_jal_N_1374), .n32630(n32630), .is_jal_de(is_jal_de), 
            .n7(n7_adj_3212), .n22(n22_adj_3179), .n32653(n32653), .n32566(n32566), 
            .n32340(n32340), .n32634(n32634), .n32637(n32637), .n32641(n32641), 
            .n32651(n32651), .n29039(n29039), .\additional_mem_ops_2__N_1132[0] (additional_mem_ops_2__N_1132[0]), 
            .n32654(n32654), .n32599(n32599), .n32659(n32659), .n32658(n32658), 
            .n32661(n32661), .n32657(n32657), .n32638(n32638), .n32640(n32640), 
            .n32582(n32582), .n32643(n32643), .n32576(n32576), .n7_adj_1(n7_adj_3196), 
            .n9(n9_adj_3180), .n8330(n8330), .n8(n8_c), .n29119(n29119), 
            .n32642(n32642), .n32655(n32655), .n32656(n32656), .n32639(n32639), 
            .n10(n10), .n24(n24), .n32594(n32594), .n2225(n2222[13]), 
            .n2156(n2151[11]), .n29748(n29748), .n34287(n34287), .n28501(n28501), 
            .\instr[16] (\instr[16] ), .n2598(n2595[1]), .n29605(n29605), 
            .n32565(n32565), .\instr[20] (instr[20]), .n32539(n32539), 
            .n27731(n27731), .n28489(n28489), .rst_reg_n(rst_reg_n_adj_6), 
            .n10024(n10024), .n28575(n28575), .n29681(n29681), .is_load_de(is_load_de), 
            .\instr[25] (instr[25]), .n3355(n3328[5]), .n672(n672), .mem_op_increment_reg_de(mem_op_increment_reg_de), 
            .n32571(n32571), .n2157(n2151[10]), .n29725(n29725), .n32540(n32540), 
            .n32734(n32734), .n30041(n30041), .n32573(n32573), .n4251(n4251), 
            .n32533(n32533), .\alu_op_3__N_1170[1] (alu_op_3__N_1170[1]), 
            .n26937(n26937), .n27(n27), .\instr[30] (instr[30]), .n3(n3_adj_3194), 
            .n156(n155[3]), .n32563(n32563), .n41(n41), .n30(n30_adj_3211), 
            .n22_adj_2(n22_adj_3213), .n32629(n32629), .\alu_op_3__N_1337[2] (alu_op_3__N_1337[2]), 
            .n32585(n32585), .n32(n32), .n4257(n4257), .n3253(n3222[1]), 
            .n32176(n32176), .n32609(n32609), .n4259(n4259), .n3286(n3259[5]), 
            .n3288(n3259[3]), .n32577(n32577), .n3290(n3259[1]), .n3289(n3259[2]), 
            .n29025(n29025), .n28577(n28577), .n32615(n32615), .n32597(n32597), 
            .n32222(n32222), .n9394(n9394), .\instr[29] (instr[29]), .\instr[31] (\instr[31] ), 
            .n5207(n5205[29]), .\instr[24] (instr[24]), .n5212(n5205[24]), 
            .n5222(n5205[14]), .\instr[19] (instr[19]), .n32030(n32030), 
            .n5221(n5205[15]), .n2205(n2202[13]), .n5224(n5205[12]), .n29716(n29716), 
            .n29705(n29705), .n32025(n32025), .n32024(n32024), .n29712(n29712), 
            .n29695(n29695), .\instr[28] (instr[28]), .n5208(n5205[28]), 
            .n5220(n5205[16]), .n5211(n5205[25]), .n29714(n29714), .n29697(n29697), 
            .n32016(n32016), .n32017(n32017), .n29726(n29726), .n29718(n29718), 
            .n29703(n29703), .n5223(n5205[13]), .n29747(n29747), .n2153(n2151[14]), 
            .n29732(n29732), .n32583(n32583), .is_auipc_de(is_auipc_de), 
            .n5231(n5205[5]), .n32559(n32559), .n5236(n5205[0]), .n5232(n5205[4]), 
            .n32569(n32569), .n32617(n32617), .n32618(n32618), .is_system_de(is_system_de), 
            .n29211(n29211), .is_store_de(is_store_de), .\instr[26] (instr[26]), 
            .n32627(n32627), .is_alu_imm_de(is_alu_imm_de), .n32581(n32581), 
            .n29031(n29031), .n32603(n32603), .n2986(n2970[16]), .n331(n328[1]), 
            .n32602(n32602), .n32596(n32596), .n11066(n11066), .n29723(n29723), 
            .n32570(n32570), .n28919(n28919), .\instr[23] (instr[23]), 
            .n28791(n28791), .\instr[22] (instr[22]), .n28763(n28763), 
            .\instr[21] (instr[21]), .n28805(n28805), .n28777(n28777), 
            .n31698(n31698), .n32619(n32619), .n32633(n32633), .is_branch_de(is_branch_de), 
            .n32589(n32589), .\mem_op_de[2] (mem_op_de[2]), .n28617(n28617), 
            .n26(n26), .n28623(n28623), .n28593(n28593), .n28599(n28599), 
            .n4(n4_c), .n28539(n28539), .n28653(n28653), .n28659(n28659), 
            .n2798(n2798), .\instr[17] (instr[17]), .n2592(n2590[2]), 
            .n2620(n2618[2]), .n28561(n28561), .n28567(n28567), .n28641(n28641), 
            .n28647(n28647), .n28547(n28547), .n28553(n28553), .n28605(n28605), 
            .n28611(n28611), .n12(n12_adj_3169), .n28527(n28527), .n28407(n28407), 
            .n19(n19_c), .n28413(n28413), .n26879(n26879), .n28669(n28669), 
            .n19_adj_3(n19_adj_3201), .n27959(n27959), .alu_op_de({alu_op_de}), 
            .n32613(n32613), .n28363(n28363), .n27788(n27788), .n9048(n9048), 
            .n30919(n30919), .n32610(n32610), .n9052(n9052), .n30920(n30920), 
            .n32612(n32612), .n32190(n32190), .n32541(n32541), .n17665(n17665), 
            .n4_adj_4(n4_adj_3177), .n32580(n32580), .n2994(n2970[8]), 
            .is_alu_reg_de(is_alu_reg_de), .n2136(n2131[11]), .n32360(n32360), 
            .is_jalr_de(is_jalr_de), .is_lui_N_1365(is_lui_N_1365), .is_lui_de(is_lui_de), 
            .n32427(n32427), .n26863(n26863), .n19_adj_5(n19_adj_3214), 
            .n24898(n24898), .n24900(n24900)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    tinyqv_core i_core (.\imm[6] (\imm[6] ), .clk_c(clk_c), .n32840(n32840), 
            .mip_reg({Open_114, mip_reg[16]}), .clk_c_enable_342(clk_c_enable_342), 
            .n32650(n32650), .n32351(n32351), .counter_hi({counter_hi}), 
            .\imm[10] (\imm[10] ), .\imm[0] (imm_c[0]), .n32759(n32759), 
            .\imm[2] (\imm[2] ), .\debug_branch_N_450[1] (debug_branch_N_450[1]), 
            .n5660(n5658[2]), .n5661(n5658[1]), .n30329(n30329), .n32309(n32309), 
            .instr_complete_N_1647(instr_complete_N_1647), .clk_c_enable_285(clk_c_enable_285), 
            .cycle({cycle[1], \cycle[0] }), .\alu_op[0] (alu_op[0]), .\alu_op[1] (alu_op[1]), 
            .is_system(is_system), .debug_instr_valid(debug_instr_valid), 
            .n32702(n32702), .n32733(n32733), .n32704(n32704), .n32746(n32746), 
            .\ui_in_sync[1] (\ui_in_sync[1] ), .n24384(n24384), .stall_core(stall_core), 
            .n32774(n32774), .n32545(n32545), .is_load(is_load), .n829(n829), 
            .n26962(n26962), .clk_c_enable_533(clk_c_enable_533), .\alu_op_in[2] (alu_op_in[2]), 
            .\ui_in_sync[0] (\ui_in_sync[0] ), .debug_rd({debug_rd}), .\mie[10] (mie[10]), 
            .\mie[14] (mie[14]), .\mie[2] (mie[2]), .\mie[6] (mie[6]), 
            .n27294(n27294), .n5017({n5017}), .n1766(n1764[1]), .\instr_write_offset_3__N_934[1] (instr_write_offset_3__N_934[1]), 
            .n1767(n1764[0]), .\instr_write_offset_3__N_934[0] (instr_write_offset_3__N_934[0]), 
            .n1768({n1768}), .pc_2__N_932({pc_2__N_932}), .\next_pc_for_core[15] (\next_pc_for_core[15] ), 
            .\next_pc_for_core[11] (\next_pc_for_core[11] ), .n32846(n32846), 
            .n32847(n32847), .\imm[7] (\imm[7] ), .n9058(n9058), .n29689(n29689), 
            .n32691(n32691), .n32549(n32549), .n32543(n32543), .instr_fetch_running(instr_fetch_running), 
            .was_early_branch(was_early_branch), .n32550(n32550), .n32564(n32564), 
            .data_ready_sync(data_ready_sync), .data_ready_core(data_ready_core), 
            .n131(n131), .n32768(n32768), .n32849(n32849), .n32697(n32697), 
            .clk_c_enable_538(clk_c_enable_538), .\imm[1] (\imm[1] ), .n32838(n32838), 
            .n29866(n29866), .clk_c_enable_433(clk_c_enable_433), .n32854(n32854), 
            .interrupt_core(interrupt_core), .rst_reg_n(rst_reg_n_adj_6), 
            .n17920(n17920), .n28685(n28685), .n28687(n28687), .n34285(n34285), 
            .is_lui(is_lui), .is_jal(is_jal), .is_branch(is_branch), .is_jalr(is_jalr), 
            .is_auipc(is_auipc), .n34281(n34281), .n32551(n32551), .mstatus_mte(mstatus_mte), 
            .n92({n92}), .n34287(n34287), .n27003(n27003), .n32821(n32821), 
            .mem_op({mem_op}), .n32741(n32741), .\alu_op[3] (alu_op[3]), 
            .accum({accum}), .d_3__N_1868({d_3__N_1868}), .data_out_3__N_1385(data_out_3__N_1385), 
            .is_timer_addr(is_timer_addr), .n30160(n30160), .n32784(n32784), 
            .n32677(n32677), .debug_rd_3__N_1575(debug_rd_3__N_1575), .\imm[11] (\imm[11] ), 
            .clk_c_enable_276(clk_c_enable_276), .fsm_state({fsm_state_adj_14}), 
            .n32791(n32791), .n32763(n32763), .n32730(n32730), .timer_interrupt(timer_interrupt), 
            .n32765(n32765), .n5642(n5640[2]), .n926(n926), .n33057(n33057), 
            .\timer_data[0] (timer_data[0]), .clk_c_enable_321(clk_c_enable_321), 
            .n893(n893), .load_done(load_done), .clk_c_enable_363(clk_c_enable_363), 
            .n8228(n8228), .n32317(n32317), .\timer_data[2] (timer_data[2]), 
            .data_rs1({Open_115, data_rs1[2], Open_116, Open_117}), 
            .n860(n860), .n793(n793), .n32546(n32546), .n28417(n28417), 
            .n32580(n32580), .n32642(n32642), .n3274(n3259[17]), .n28429(n28429), 
            .n4(n4_adj_3177), .n27546(n27546), .n28465(n28465), .n27541(n27541), 
            .\debug_branch_N_450[3] (debug_branch_N_450[3]), .load_top_bit(load_top_bit), 
            .n32806(n32806), .n32808(n32808), .instr_complete_N_1651(instr_complete_N_1651), 
            .instr_complete_N_1652(instr_complete_N_1652), .is_double_fault_r(is_double_fault_r), 
            .n28441(n28441), .n27545(n27545), .n32732(n32732), .n8(n8_adj_3200), 
            .n5659(n5658[3]), .debug_rd_3__N_413(debug_rd_3__N_413), .n28275(n28275), 
            .n1(n1_adj_3208), .n27427(n27427), .\imm[4] (\imm[4] ), .n5607(n5605[2]), 
            .\cycle_count_wide[3] (cycle_count_wide[3]), .n28343(n28343), 
            .n32559(n32559), .n32539(n32539), .data_rs2({data_rs2}), .\data_out_slice[0] (data_out_slice[0]), 
            .n32644(n32644), .n34283(n34283), .timer_data_3__N_631(timer_data_3__N_631), 
            .\mtimecmp[7] (mtimecmp[7]), .mtimecmp_3__N_1935(mtimecmp_3__N_1935), 
            .\data_rs1[3] (data_rs1[3]), .mstatus_mie_N_1709(mstatus_mie_N_1709), 
            .\data_rs1[0] (data_rs1[0]), .\imm[9] (\imm[9] ), .\imm[8] (\imm[8] ), 
            .\addr_out[27] (addr_out[27]), .\addr_out[24] (addr_out[24]), 
            .\addr_out[25] (addr_out[25]), .\addr_out[26] (addr_out[26]), 
            .n32829(n32829), .\imm[5] (\imm[5] ), .\imm[3] (\imm[3] ), 
            .n27656(n27656), .n28909(n28909), .n27655(n27655), .n29838(n29838), 
            .n30172(n30172), .n27657(n27657), .n28533(n28533), .n32548(n32548), 
            .clk_c_enable_524(clk_c_enable_524), .n2559(n2559), .n32834(n32834), 
            .n32760(n32760), .n32758(n32758), .clk_c_enable_187(clk_c_enable_187), 
            .n28363(n28363), .n28483(n28483), .n32538(n32538), .n32828(n32828), 
            .address_ready(address_ready), .is_store(is_store), .mstatus_mie_N_1707(mstatus_mie_N_1707), 
            .n32710(n32710), .n30425(n30425), .n13(n13_adj_3173), .n29760(n29760), 
            .n32668(n32668), .\mtimecmp[5] (mtimecmp[5]), .mtimecmp_1__N_1941(mtimecmp_1__N_1941), 
            .\debug_rd_3__N_405[28] (debug_rd_3__N_405[28]), .n32848(n32848), 
            .n29844(n29844), .n32678(n32678), .n32675(n32675), .is_alu_imm(is_alu_imm), 
            .is_alu_reg(is_alu_reg), .n28889(n28889), .n27653(n27653), 
            .n31351(n31351), .n29864(n29864), .clk_c_enable_195(clk_c_enable_195), 
            .n18(n39[2]), .n29317(n29317), .n32647(n32647), .n32670(n32670), 
            .clk_c_enable_28(clk_c_enable_28), .n32552(n32552), .n32783(n32783), 
            .n30928(n30928), .n30927(n30927), .n30926(n30926), .n30925(n30925), 
            .n30924(n30924), .n32769(n32769), .\debug_branch_N_442[31] (debug_branch_N_442[31]), 
            .\debug_branch_N_442[30] (debug_branch_N_442[30]), .\debug_rd_3__N_405[30] (debug_rd_3__N_405[30]), 
            .\debug_branch_N_442[29] (debug_branch_N_442[29]), .\addr_offset[2] (addr_offset[2]), 
            .n28963(n28963), .\debug_rd_3__N_405[29] (debug_rd_3__N_405[29]), 
            .n157(n157_adj_3187), .\debug_branch_N_442[28] (debug_branch_N_442[28]), 
            .n28495(n28495), .n2124(n2124), .\debug_rd_3__N_405[31] (debug_rd_3__N_405[31]), 
            .n701(n699[0]), .\data_out_slice[2] (data_out_slice[2]), .debug_early_branch_N_955(debug_early_branch_N_955), 
            .no_write_in_progress(no_write_in_progress), .n1152(n1152), 
            .\next_pc_offset[3] (next_pc_offset[3]), .n28237(n28237), .\debug_branch_N_450[0] (debug_branch_N_450[0]), 
            .n18098(n18098), .\debug_branch_N_446[28] (debug_branch_N_446[28]), 
            .n238(n234[0]), .n30070(n30070), .n76(n76), .\mtime_out[0] (mtime_out[0]), 
            .n32717(n32717), .cy(cy), .n32663(n32663), .n9620(n9620), 
            .time_pulse_r(time_pulse_r), .n10737(n10737), .n32680(n32680), 
            .\next_pc_for_core[7] (\next_pc_for_core[7] ), .\next_pc_for_core[3] (\next_pc_for_core[3] ), 
            .\next_pc_for_core[23] (\next_pc_for_core[23] ), .\next_pc_for_core[19] (\next_pc_for_core[19] ), 
            .\addr_out[1] (addr_out[1]), .\addr_out[0] (addr_out[0]), .n32690(n32690), 
            .\addr_out[23] (addr_out[23]), .\addr_out[22] (addr_out[22]), 
            .\addr_out[21] (addr_out[21]), .\addr_out[20] (addr_out[20]), 
            .\addr_out[19] (addr_out[19]), .\addr_out[18] (addr_out[18]), 
            .\addr_out[17] (addr_out[17]), .\addr_out[16] (addr_out[16]), 
            .\addr_out[15] (addr_out[15]), .\addr_out[14] (addr_out[14]), 
            .\addr_out[13] (addr_out[13]), .\addr_out[12] (addr_out[12]), 
            .\addr_out[11] (addr_out[11]), .\addr_out[10] (addr_out[10]), 
            .\addr_out[9] (addr_out[9]), .\addr_out[8] (addr_out[8]), .\addr_out[7] (addr_out[7]), 
            .\addr_out[6] (addr_out[6]), .\addr_out[5] (addr_out[5]), .\addr_out[4] (addr_out[4]), 
            .\addr_out[3] (addr_out[3]), .\mem_data_from_read[17] (\mem_data_from_read[17] ), 
            .\mem_data_from_read[21] (\mem_data_from_read[21] ), .n32308(n32308), 
            .\timer_data[1] (timer_data[1]), .\mul_out[3] (\mul_out[3] ), 
            .\mul_out[2] (\mul_out[2] ), .rd({rd_c[3:1], rd[0]}), .n32776(n32776), 
            .\mul_out[1] (\mul_out[1] ), .\debug_branch_N_446[31] (debug_branch_N_446[31]), 
            .n30175(n30175), .n29842(n29842), .\debug_branch_N_446[30] (debug_branch_N_446[30]), 
            .\csr_read_3__N_1447[2] (\csr_read_3__N_1447[2] ), .n29836(n29836), 
            .\debug_branch_N_446[29] (debug_branch_N_446[29]), .n32767(n32767), 
            .\next_accum[5] (\next_accum[5] ), .GND_net(GND_net), .VCC_net(VCC_net), 
            .\next_accum[16] (\next_accum[16] ), .\next_accum[17] (\next_accum[17] ), 
            .\next_accum[18] (\next_accum[18] ), .\next_accum[19] (\next_accum[19] ), 
            .\next_accum[6] (\next_accum[6] ), .\next_accum[7] (\next_accum[7] ), 
            .\next_accum[8] (\next_accum[8] ), .\next_accum[9] (\next_accum[9] ), 
            .\next_accum[10] (\next_accum[10] ), .\next_accum[11] (\next_accum[11] ), 
            .\next_accum[12] (\next_accum[12] ), .\next_accum[13] (\next_accum[13] ), 
            .\next_accum[14] (\next_accum[14] ), .\next_accum[15] (\next_accum[15] ), 
            .\next_accum[4] (\next_accum[4] ), .n21667(n21667), .rs1({rs1}), 
            .rs2({rs2}), .\reg_access[3][2] (\reg_access[3] [2]), .return_addr({return_addr[23:17], 
            \return_addr[16] , return_addr[15:1]}), .\reg_access[4][3] (\reg_access[4] [3]), 
            .n32652(n32652)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(322[72] 368[6])
    
endmodule
//
// Verilog Description of module tinyQV_time
//

module tinyQV_time (clk_c, n32840, time_pulse_r, clk_c_enable_363, n32717, 
            \data_rs2[2] , data_out_3__N_1385, timer_data_3__N_631, \data_rs2[0] , 
            \mtimecmp[7] , \mtimecmp[5] , clk_c_enable_285, mtimecmp_1__N_1941, 
            mtime_out, \addr[2] , timer_data, timer_interrupt, mtimecmp_3__N_1935, 
            n10737, cy, n32663, n32680, rst_reg_n, is_timer_addr, 
            n32801, n32653, n32654, n32588, no_write_in_progress, 
            is_store, clk_c_enable_178, mstatus_mie_N_1709, n32670, 
            n32675, mstatus_mie_N_1707, n32765, clk_c_enable_207, n34287, 
            n32758, n32746, n32759, clk_c_enable_433, \instr_addr_23__N_318[1] , 
            \instr_addr_23__N_318[0] , n28739, n32691, n29317, n32548, 
            n32541, clk_c_enable_338, \reg_access[4][3] , clk_c_enable_182, 
            n32760, clk_c_enable_191, address_ready, n32671, n28747, 
            \instr_data[1] , \instr_data_0__15__N_638[49] , \reg_access[3][2] , 
            clk_c_enable_200, n28755, \instr_data[0] , \instr_data_0__15__N_638[0] , 
            \cycle_count_wide[3] , n32652, clk_c_enable_276, clk_c_enable_204, 
            n32611, n10024, n32630, n28391, n32697, is_double_fault_r, 
            mstatus_mte, n32650, clk_c_enable_99, clk_c_enable_174, 
            n32668, n32664, \data_out_slice[0] , n32644, \data_out_slice[2] ) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output n32840;
    output time_pulse_r;
    input clk_c_enable_363;
    output n32717;
    input \data_rs2[2] ;
    input data_out_3__N_1385;
    input timer_data_3__N_631;
    input \data_rs2[0] ;
    output \mtimecmp[7] ;
    output \mtimecmp[5] ;
    input clk_c_enable_285;
    input mtimecmp_1__N_1941;
    output [3:0]mtime_out;
    input \addr[2] ;
    output [3:0]timer_data;
    output timer_interrupt;
    input mtimecmp_3__N_1935;
    input n10737;
    output cy;
    input n32663;
    input n32680;
    input rst_reg_n;
    input is_timer_addr;
    input n32801;
    input n32653;
    input n32654;
    output n32588;
    input no_write_in_progress;
    input is_store;
    output clk_c_enable_178;
    input mstatus_mie_N_1709;
    input n32670;
    input n32675;
    output mstatus_mie_N_1707;
    input n32765;
    output clk_c_enable_207;
    input n34287;
    output n32758;
    input n32746;
    input n32759;
    output clk_c_enable_433;
    input \instr_addr_23__N_318[1] ;
    input \instr_addr_23__N_318[0] ;
    output n28739;
    input n32691;
    output n29317;
    input n32548;
    input n32541;
    output clk_c_enable_338;
    input \reg_access[4][3] ;
    output clk_c_enable_182;
    input n32760;
    output clk_c_enable_191;
    input address_ready;
    output n32671;
    output n28747;
    input \instr_data[1] ;
    output \instr_data_0__15__N_638[49] ;
    input \reg_access[3][2] ;
    output clk_c_enable_200;
    output n28755;
    input \instr_data[0] ;
    output \instr_data_0__15__N_638[0] ;
    input \cycle_count_wide[3] ;
    input n32652;
    output clk_c_enable_276;
    output clk_c_enable_204;
    input n32611;
    input n10024;
    input n32630;
    output n28391;
    input n32697;
    input is_double_fault_r;
    input mstatus_mte;
    output n32650;
    output clk_c_enable_99;
    output clk_c_enable_174;
    input n32668;
    input n32664;
    input \data_out_slice[0] ;
    input n32644;
    input \data_out_slice[2] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [31:0]mtimecmp;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(30[16:24])
    
    wire mtimecmp_0__N_1943, mtimecmp_2__N_1939, cy_c;
    wire [4:0]comparison;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[16:26])
    wire [3:0]mtime_out_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(29[16:25])
    
    wire timer_interrupt_N_1954, n4, n32867, n32866, n6, n2;
    
    FD1S3IX mtimecmp_0__92 (.D(mtimecmp_0__N_1943), .CK(clk_c), .CD(n32840), 
            .Q(mtimecmp[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_0__92.GSR = "DISABLED";
    FD1S3IX time_pulse_r_95 (.D(n32717), .CK(clk_c), .CD(clk_c_enable_363), 
            .Q(time_pulse_r)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(82[12] 85[8])
    defparam time_pulse_r_95.GSR = "DISABLED";
    LUT4 mtimecmp_6__I_0_3_lut_4_lut (.A(mtimecmp[6]), .B(\data_rs2[2] ), 
         .C(data_out_3__N_1385), .D(timer_data_3__N_631), .Z(mtimecmp_2__N_1939)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(67[18:49])
    defparam mtimecmp_6__I_0_3_lut_4_lut.init = 16'h0caa;
    LUT4 mtimecmp_4__I_0_3_lut_4_lut (.A(mtimecmp[4]), .B(\data_rs2[0] ), 
         .C(data_out_3__N_1385), .D(timer_data_3__N_631), .Z(mtimecmp_0__N_1943)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(67[18:49])
    defparam mtimecmp_4__I_0_3_lut_4_lut.init = 16'h0caa;
    FD1S3AX mtimecmp_30__62 (.D(mtimecmp[2]), .CK(clk_c), .Q(mtimecmp[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_30__62.GSR = "DISABLED";
    FD1S3AX mtimecmp_29__63 (.D(mtimecmp[1]), .CK(clk_c), .Q(mtimecmp[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_29__63.GSR = "DISABLED";
    FD1S3AX mtimecmp_28__64 (.D(mtimecmp[0]), .CK(clk_c), .Q(mtimecmp[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_28__64.GSR = "DISABLED";
    FD1S3AX mtimecmp_27__65 (.D(mtimecmp[31]), .CK(clk_c), .Q(mtimecmp[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_27__65.GSR = "DISABLED";
    FD1S3AX mtimecmp_26__66 (.D(mtimecmp[30]), .CK(clk_c), .Q(mtimecmp[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_26__66.GSR = "DISABLED";
    FD1S3AX mtimecmp_25__67 (.D(mtimecmp[29]), .CK(clk_c), .Q(mtimecmp[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_25__67.GSR = "DISABLED";
    FD1S3AX mtimecmp_24__68 (.D(mtimecmp[28]), .CK(clk_c), .Q(mtimecmp[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_24__68.GSR = "DISABLED";
    FD1S3AX mtimecmp_23__69 (.D(mtimecmp[27]), .CK(clk_c), .Q(mtimecmp[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_23__69.GSR = "DISABLED";
    FD1S3AX mtimecmp_22__70 (.D(mtimecmp[26]), .CK(clk_c), .Q(mtimecmp[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_22__70.GSR = "DISABLED";
    FD1S3AX mtimecmp_21__71 (.D(mtimecmp[25]), .CK(clk_c), .Q(mtimecmp[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_21__71.GSR = "DISABLED";
    FD1S3AX mtimecmp_20__72 (.D(mtimecmp[24]), .CK(clk_c), .Q(mtimecmp[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_20__72.GSR = "DISABLED";
    FD1S3AX mtimecmp_19__73 (.D(mtimecmp[23]), .CK(clk_c), .Q(mtimecmp[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_19__73.GSR = "DISABLED";
    FD1S3AX mtimecmp_18__74 (.D(mtimecmp[22]), .CK(clk_c), .Q(mtimecmp[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_18__74.GSR = "DISABLED";
    FD1S3AX mtimecmp_17__75 (.D(mtimecmp[21]), .CK(clk_c), .Q(mtimecmp[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_17__75.GSR = "DISABLED";
    FD1S3AX mtimecmp_16__76 (.D(mtimecmp[20]), .CK(clk_c), .Q(mtimecmp[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_16__76.GSR = "DISABLED";
    FD1S3AX mtimecmp_15__77 (.D(mtimecmp[19]), .CK(clk_c), .Q(mtimecmp[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_15__77.GSR = "DISABLED";
    FD1S3AX mtimecmp_14__78 (.D(mtimecmp[18]), .CK(clk_c), .Q(mtimecmp[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_14__78.GSR = "DISABLED";
    FD1S3AX mtimecmp_13__79 (.D(mtimecmp[17]), .CK(clk_c), .Q(mtimecmp[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_13__79.GSR = "DISABLED";
    FD1S3AX mtimecmp_12__80 (.D(mtimecmp[16]), .CK(clk_c), .Q(mtimecmp[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_12__80.GSR = "DISABLED";
    FD1S3AX mtimecmp_11__81 (.D(mtimecmp[15]), .CK(clk_c), .Q(mtimecmp[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_11__81.GSR = "DISABLED";
    FD1S3AX mtimecmp_10__82 (.D(mtimecmp[14]), .CK(clk_c), .Q(mtimecmp[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_10__82.GSR = "DISABLED";
    FD1S3AX mtimecmp_9__83 (.D(mtimecmp[13]), .CK(clk_c), .Q(mtimecmp[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_9__83.GSR = "DISABLED";
    FD1S3AX mtimecmp_8__84 (.D(mtimecmp[12]), .CK(clk_c), .Q(mtimecmp[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_8__84.GSR = "DISABLED";
    FD1S3AX mtimecmp_7__85 (.D(mtimecmp[11]), .CK(clk_c), .Q(\mtimecmp[7] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_7__85.GSR = "DISABLED";
    FD1S3AX mtimecmp_6__86 (.D(mtimecmp[10]), .CK(clk_c), .Q(mtimecmp[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_6__86.GSR = "DISABLED";
    FD1S3AX mtimecmp_5__87 (.D(mtimecmp[9]), .CK(clk_c), .Q(\mtimecmp[5] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_5__87.GSR = "DISABLED";
    FD1S3AX mtimecmp_4__88 (.D(mtimecmp[8]), .CK(clk_c), .Q(mtimecmp[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_4__88.GSR = "DISABLED";
    FD1S3JX cy_93 (.D(comparison[4]), .CK(clk_c), .PD(clk_c_enable_285), 
            .Q(cy_c)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(74[12] 76[8])
    defparam cy_93.GSR = "DISABLED";
    FD1S3IX mtimecmp_1__91 (.D(mtimecmp_1__N_1941), .CK(clk_c), .CD(n32840), 
            .Q(mtimecmp[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_1__91.GSR = "DISABLED";
    FD1S3AX mtimecmp_31__61 (.D(mtimecmp[3]), .CK(clk_c), .Q(mtimecmp[31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_31__61.GSR = "DISABLED";
    LUT4 mtime_out_3__I_0_96_i1_3_lut (.A(mtime_out[0]), .B(mtimecmp[4]), 
         .C(\addr[2] ), .Z(timer_data[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i1_3_lut.init = 16'hcaca;
    LUT4 mtime_out_3__I_0_96_i2_3_lut (.A(mtime_out_c[1]), .B(\mtimecmp[5] ), 
         .C(\addr[2] ), .Z(timer_data[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i2_3_lut.init = 16'hcaca;
    LUT4 mtime_out_3__I_0_96_i3_3_lut (.A(mtime_out_c[2]), .B(mtimecmp[6]), 
         .C(\addr[2] ), .Z(timer_data[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i3_3_lut.init = 16'hcaca;
    FD1P3AX timer_interrupt_94 (.D(timer_interrupt_N_1954), .SP(clk_c_enable_285), 
            .CK(clk_c), .Q(timer_interrupt)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(78[12] 80[8])
    defparam timer_interrupt_94.GSR = "DISABLED";
    FD1S3IX mtimecmp_3__89 (.D(mtimecmp_3__N_1935), .CK(clk_c), .CD(n32840), 
            .Q(mtimecmp[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_3__89.GSR = "DISABLED";
    FD1S3IX mtimecmp_2__90 (.D(mtimecmp_2__N_1939), .CK(clk_c), .CD(n32840), 
            .Q(mtimecmp[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_2__90.GSR = "DISABLED";
    LUT4 i15198_4_lut_then_4_lut (.A(mtime_out_c[3]), .B(n4), .C(mtimecmp[6]), 
         .D(\mtimecmp[7] ), .Z(n32867)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;
    defparam i15198_4_lut_then_4_lut.init = 16'h8241;
    LUT4 i15198_4_lut_else_4_lut (.A(mtime_out_c[3]), .B(n4), .C(mtimecmp[6]), 
         .D(\mtimecmp[7] ), .Z(n32866)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A (B (C+(D))+!B !(C (D))))) */ ;
    defparam i15198_4_lut_else_4_lut.init = 16'h1824;
    PFUMX i29311 (.BLUT(n32866), .ALUT(n32867), .C0(mtime_out_c[2]), .Z(timer_interrupt_N_1954));
    LUT4 i4575_3_lut (.A(mtime_out_c[3]), .B(\mtimecmp[7] ), .C(n6), .Z(comparison[4])) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i4575_3_lut.init = 16'hb2b2;
    LUT4 mtime_out_3__I_0_96_i4_3_lut (.A(mtime_out_c[3]), .B(\mtimecmp[7] ), 
         .C(\addr[2] ), .Z(timer_data[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i4_3_lut.init = 16'hcaca;
    LUT4 i4568_3_lut (.A(mtime_out_c[2]), .B(mtimecmp[6]), .C(n4), .Z(n6)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i4568_3_lut.init = 16'hb2b2;
    LUT4 i4561_3_lut (.A(mtime_out_c[1]), .B(\mtimecmp[5] ), .C(n2), .Z(n4)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i4561_3_lut.init = 16'hb2b2;
    LUT4 time_pulse_I_0_2_lut_rep_702 (.A(n10737), .B(time_pulse_r), .Z(n32717)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(37[14:39])
    defparam time_pulse_I_0_2_lut_rep_702.init = 16'hdddd;
    LUT4 i4554_3_lut (.A(mtime_out[0]), .B(mtimecmp[4]), .C(cy_c), .Z(n2)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i4554_3_lut.init = 16'hb2b2;
    tinyqv_counter i_mtime (.clk_c(clk_c), .n32840(n32840), .cy(cy), .mtime_out({mtime_out_c[3:1], 
            mtime_out[0]}), .n32663(n32663), .n32680(n32680), .rst_reg_n(rst_reg_n), 
            .is_timer_addr(is_timer_addr), .n32801(n32801), .\addr[2] (\addr[2] ), 
            .n32653(n32653), .n32654(n32654), .n32588(n32588), .clk_c_enable_285(clk_c_enable_285), 
            .no_write_in_progress(no_write_in_progress), .is_store(is_store), 
            .clk_c_enable_178(clk_c_enable_178), .mstatus_mie_N_1709(mstatus_mie_N_1709), 
            .n32670(n32670), .n32675(n32675), .mstatus_mie_N_1707(mstatus_mie_N_1707), 
            .n32765(n32765), .clk_c_enable_207(clk_c_enable_207), .n34287(n34287), 
            .n32758(n32758), .n32746(n32746), .n32759(n32759), .clk_c_enable_433(clk_c_enable_433), 
            .\instr_addr_23__N_318[1] (\instr_addr_23__N_318[1] ), .\instr_addr_23__N_318[0] (\instr_addr_23__N_318[0] ), 
            .n28739(n28739), .n32691(n32691), .n29317(n29317), .n32548(n32548), 
            .n32541(n32541), .clk_c_enable_338(clk_c_enable_338), .\reg_access[4][3] (\reg_access[4][3] ), 
            .clk_c_enable_182(clk_c_enable_182), .n32760(n32760), .clk_c_enable_191(clk_c_enable_191), 
            .address_ready(address_ready), .n32671(n32671), .n28747(n28747), 
            .\instr_data[1] (\instr_data[1] ), .\instr_data_0__15__N_638[49] (\instr_data_0__15__N_638[49] ), 
            .\reg_access[3][2] (\reg_access[3][2] ), .clk_c_enable_200(clk_c_enable_200), 
            .n28755(n28755), .\instr_data[0] (\instr_data[0] ), .\instr_data_0__15__N_638[0] (\instr_data_0__15__N_638[0] ), 
            .\cycle_count_wide[3] (\cycle_count_wide[3] ), .n32652(n32652), 
            .clk_c_enable_276(clk_c_enable_276), .clk_c_enable_204(clk_c_enable_204), 
            .n32611(n32611), .n10024(n10024), .n32630(n32630), .n28391(n28391), 
            .n32697(n32697), .is_double_fault_r(is_double_fault_r), .mstatus_mte(mstatus_mte), 
            .n32650(n32650), .clk_c_enable_99(clk_c_enable_99), .clk_c_enable_174(clk_c_enable_174), 
            .n32668(n32668), .n32664(n32664), .\data_out_slice[0] (\data_out_slice[0] ), 
            .n32644(n32644), .\data_out_slice[2] (\data_out_slice[2] )) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(34[20] 42[6])
    
endmodule
//
// Verilog Description of module tinyqv_counter
//

module tinyqv_counter (clk_c, n32840, cy, mtime_out, n32663, n32680, 
            rst_reg_n, is_timer_addr, n32801, \addr[2] , n32653, n32654, 
            n32588, clk_c_enable_285, no_write_in_progress, is_store, 
            clk_c_enable_178, mstatus_mie_N_1709, n32670, n32675, mstatus_mie_N_1707, 
            n32765, clk_c_enable_207, n34287, n32758, n32746, n32759, 
            clk_c_enable_433, \instr_addr_23__N_318[1] , \instr_addr_23__N_318[0] , 
            n28739, n32691, n29317, n32548, n32541, clk_c_enable_338, 
            \reg_access[4][3] , clk_c_enable_182, n32760, clk_c_enable_191, 
            address_ready, n32671, n28747, \instr_data[1] , \instr_data_0__15__N_638[49] , 
            \reg_access[3][2] , clk_c_enable_200, n28755, \instr_data[0] , 
            \instr_data_0__15__N_638[0] , \cycle_count_wide[3] , n32652, 
            clk_c_enable_276, clk_c_enable_204, n32611, n10024, n32630, 
            n28391, n32697, is_double_fault_r, mstatus_mte, n32650, 
            clk_c_enable_99, clk_c_enable_174, n32668, n32664, \data_out_slice[0] , 
            n32644, \data_out_slice[2] ) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output n32840;
    output cy;
    output [3:0]mtime_out;
    input n32663;
    input n32680;
    input rst_reg_n;
    input is_timer_addr;
    input n32801;
    input \addr[2] ;
    input n32653;
    input n32654;
    output n32588;
    input clk_c_enable_285;
    input no_write_in_progress;
    input is_store;
    output clk_c_enable_178;
    input mstatus_mie_N_1709;
    input n32670;
    input n32675;
    output mstatus_mie_N_1707;
    input n32765;
    output clk_c_enable_207;
    input n34287;
    output n32758;
    input n32746;
    input n32759;
    output clk_c_enable_433;
    input \instr_addr_23__N_318[1] ;
    input \instr_addr_23__N_318[0] ;
    output n28739;
    input n32691;
    output n29317;
    input n32548;
    input n32541;
    output clk_c_enable_338;
    input \reg_access[4][3] ;
    output clk_c_enable_182;
    input n32760;
    output clk_c_enable_191;
    input address_ready;
    output n32671;
    output n28747;
    input \instr_data[1] ;
    output \instr_data_0__15__N_638[49] ;
    input \reg_access[3][2] ;
    output clk_c_enable_200;
    output n28755;
    input \instr_data[0] ;
    output \instr_data_0__15__N_638[0] ;
    input \cycle_count_wide[3] ;
    input n32652;
    output clk_c_enable_276;
    output clk_c_enable_204;
    input n32611;
    input n10024;
    input n32630;
    output n28391;
    input n32697;
    input is_double_fault_r;
    input mstatus_mte;
    output n32650;
    output clk_c_enable_99;
    output clk_c_enable_174;
    input n32668;
    input n32664;
    input \data_out_slice[0] ;
    input n32644;
    input \data_out_slice[2] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    wire [4:0]increment_result;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[16:32])
    
    wire n9391;
    wire [4:0]increment_result_3__N_1925;
    
    wire n32635, n32606;
    
    FD1S3IX register_2__48 (.D(increment_result[2]), .CK(clk_c), .CD(n32840), 
            .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result[1]), .CK(clk_c), .CD(n32840), 
            .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(increment_result[0]), .CK(clk_c), .CD(n32840), 
            .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3IX cy_51 (.D(increment_result_3__N_1925[4]), .CK(clk_c), .CD(n9391), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(register[10])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(register[9])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(register[8])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(mtime_out[3])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(register[10]), .CK(clk_c), .Q(mtime_out[2])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(register[9]), .CK(clk_c), .Q(mtime_out[1])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(register[8]), .CK(clk_c), .Q(mtime_out[0])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result[3]), .CK(clk_c), .CD(n32840), 
            .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 i4858_2_lut_3_lut_4_lut (.A(mtime_out[1]), .B(n32663), .C(mtime_out[3]), 
         .D(mtime_out[2]), .Z(increment_result_3__N_1925[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4858_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4844_2_lut_rep_620_3_lut (.A(mtime_out[0]), .B(n32680), .C(mtime_out[1]), 
         .Z(n32635)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4844_2_lut_rep_620_3_lut.init = 16'h8080;
    LUT4 i4851_2_lut_rep_591_3_lut_4_lut (.A(mtime_out[0]), .B(n32680), 
         .C(mtime_out[2]), .D(mtime_out[1]), .Z(n32606)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4851_2_lut_rep_591_3_lut_4_lut.init = 16'h8000;
    LUT4 rstn_I_0_1_lut_rep_825 (.A(rst_reg_n), .Z(n32840)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam rstn_I_0_1_lut_rep_825.init = 16'h5555;
    LUT4 i6710_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(is_timer_addr), 
         .C(n32801), .D(\addr[2] ), .Z(n9391)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i6710_2_lut_3_lut_4_lut_4_lut.init = 16'h555d;
    LUT4 i15119_2_lut_rep_573_3_lut_3_lut (.A(rst_reg_n), .B(n32653), .C(n32654), 
         .Z(n32588)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i15119_2_lut_rep_573_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i15791_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(clk_c_enable_285), 
         .C(no_write_in_progress), .D(is_store), .Z(clk_c_enable_178)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i15791_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i15082_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(mstatus_mie_N_1709), 
         .C(n32670), .D(n32675), .Z(mstatus_mie_N_1707)) /* synthesis lut_function=((B ((D)+!C)+!B (D))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i15082_3_lut_4_lut_4_lut.init = 16'hff5d;
    LUT4 i28301_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n32765), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_207)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i28301_2_lut_4_lut_4_lut.init = 16'h3111;
    LUT4 i3802_3_lut_rep_743_3_lut (.A(n34287), .B(no_write_in_progress), 
         .C(is_store), .Z(n32758)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3802_3_lut_rep_743_3_lut.init = 16'hd5d5;
    LUT4 i1_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(n32746), .C(n32759), 
         .D(n32675), .Z(clk_c_enable_433)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_3_lut (.A(n34287), .B(\instr_addr_23__N_318[1] ), 
         .C(\instr_addr_23__N_318[0] ), .Z(n28739)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n34287), .B(n32675), .C(n32691), 
         .D(n32765), .Z(n29317)) /* synthesis lut_function=((B+!((D)+!C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hddfd;
    LUT4 i1_2_lut_3_lut_3_lut_adj_389 (.A(rst_reg_n), .B(n32548), .C(n32541), 
         .Z(clk_c_enable_338)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_3_lut_adj_389.init = 16'h7575;
    LUT4 i28431_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(\reg_access[4][3] ), 
         .C(no_write_in_progress), .D(is_store), .Z(clk_c_enable_182)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i28431_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i28406_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n32760), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_191)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i28406_2_lut_4_lut_4_lut.init = 16'h3111;
    LUT4 i1_2_lut_rep_656_3_lut_3_lut (.A(rst_reg_n), .B(address_ready), 
         .C(is_store), .Z(n32671)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_rep_656_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i1_2_lut_3_lut_3_lut_adj_390 (.A(n34287), .B(\instr_addr_23__N_318[1] ), 
         .C(\instr_addr_23__N_318[0] ), .Z(n28747)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_3_lut_adj_390.init = 16'hdfdf;
    LUT4 i15021_2_lut_2_lut (.A(rst_reg_n), .B(\instr_data[1] ), .Z(\instr_data_0__15__N_638[49] )) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i15021_2_lut_2_lut.init = 16'hdddd;
    LUT4 i28377_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(\reg_access[3][2] ), 
         .C(no_write_in_progress), .D(is_store), .Z(clk_c_enable_200)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i28377_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i1_2_lut_3_lut_3_lut_adj_391 (.A(n34287), .B(\instr_addr_23__N_318[0] ), 
         .C(\instr_addr_23__N_318[1] ), .Z(n28755)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_3_lut_adj_391.init = 16'hfdfd;
    LUT4 i14912_2_lut_2_lut (.A(rst_reg_n), .B(\instr_data[0] ), .Z(\instr_data_0__15__N_638[0] )) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i14912_2_lut_2_lut.init = 16'hdddd;
    LUT4 i3831_4_lut_4_lut (.A(n34287), .B(\cycle_count_wide[3] ), .C(n32652), 
         .D(clk_c_enable_285), .Z(clk_c_enable_276)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3831_4_lut_4_lut.init = 16'hd555;
    LUT4 i28376_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n32759), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_204)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i28376_2_lut_4_lut_4_lut.init = 16'h3111;
    LUT4 i1_3_lut_4_lut_4_lut_adj_392 (.A(rst_reg_n), .B(n32611), .C(n10024), 
         .D(n32630), .Z(n28391)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_3_lut_4_lut_4_lut_adj_392.init = 16'hfff7;
    LUT4 rstn_N_1579_I_0_2_lut_rep_635_4_lut_4_lut (.A(rst_reg_n), .B(n32697), 
         .C(is_double_fault_r), .D(mstatus_mte), .Z(n32650)) /* synthesis lut_function=((B (C+!(D))+!B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam rstn_N_1579_I_0_2_lut_rep_635_4_lut_4_lut.init = 16'hf5fd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_393 (.A(rst_reg_n), .B(clk_c_enable_285), 
         .C(address_ready), .D(is_store), .Z(clk_c_enable_99)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_393.init = 16'hfddd;
    LUT4 i3799_2_lut_2_lut (.A(rst_reg_n), .B(address_ready), .Z(clk_c_enable_174)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3799_2_lut_2_lut.init = 16'hdddd;
    LUT4 increment_result_3__I_168_i2_4_lut (.A(mtime_out[1]), .B(n32668), 
         .C(n32664), .D(n32663), .Z(increment_result[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i2_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_168_i1_4_lut (.A(mtime_out[0]), .B(\data_out_slice[0] ), 
         .C(n32664), .D(n32680), .Z(increment_result[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i1_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_168_i4_4_lut (.A(mtime_out[3]), .B(n32644), 
         .C(n32664), .D(n32606), .Z(increment_result[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i4_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_168_i3_4_lut (.A(mtime_out[2]), .B(\data_out_slice[2] ), 
         .C(n32664), .D(n32635), .Z(increment_result[2])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i3_4_lut.init = 16'hc5ca;
    
endmodule
//
// Verilog Description of module tinyqv_decoder
//

module tinyqv_decoder (n32361, n32623, n32362, is_jal_N_1374, n32630, 
            is_jal_de, n7, n22, n32653, n32566, n32340, n32634, 
            n32637, n32641, n32651, n29039, \additional_mem_ops_2__N_1132[0] , 
            n32654, n32599, n32659, n32658, n32661, n32657, n32638, 
            n32640, n32582, n32643, n32576, n7_adj_1, n9, n8330, 
            n8, n29119, n32642, n32655, n32656, n32639, n10, n24, 
            n32594, n2225, n2156, n29748, n34287, n28501, \instr[16] , 
            n2598, n29605, n32565, \instr[20] , n32539, n27731, 
            n28489, rst_reg_n, n10024, n28575, n29681, is_load_de, 
            \instr[25] , n3355, n672, mem_op_increment_reg_de, n32571, 
            n2157, n29725, n32540, n32734, n30041, n32573, n4251, 
            n32533, \alu_op_3__N_1170[1] , n26937, n27, \instr[30] , 
            n3, n156, n32563, n41, n30, n22_adj_2, n32629, \alu_op_3__N_1337[2] , 
            n32585, n32, n4257, n3253, n32176, n32609, n4259, 
            n3286, n3288, n32577, n3290, n3289, n29025, n28577, 
            n32615, n32597, n32222, n9394, \instr[29] , \instr[31] , 
            n5207, \instr[24] , n5212, n5222, \instr[19] , n32030, 
            n5221, n2205, n5224, n29716, n29705, n32025, n32024, 
            n29712, n29695, \instr[28] , n5208, n5220, n5211, n29714, 
            n29697, n32016, n32017, n29726, n29718, n29703, n5223, 
            n29747, n2153, n29732, n32583, is_auipc_de, n5231, n32559, 
            n5236, n5232, n32569, n32617, n32618, is_system_de, 
            n29211, is_store_de, \instr[26] , n32627, is_alu_imm_de, 
            n32581, n29031, n32603, n2986, n331, n32602, n32596, 
            n11066, n29723, n32570, n28919, \instr[23] , n28791, 
            \instr[22] , n28763, \instr[21] , n28805, n28777, n31698, 
            n32619, n32633, is_branch_de, n32589, \mem_op_de[2] , 
            n28617, n26, n28623, n28593, n28599, n4, n28539, n28653, 
            n28659, n2798, \instr[17] , n2592, n2620, n28561, n28567, 
            n28641, n28647, n28547, n28553, n28605, n28611, n12, 
            n28527, n28407, n19, n28413, n26879, n28669, n19_adj_3, 
            n27959, alu_op_de, n32613, n28363, n27788, n9048, n30919, 
            n32610, n9052, n30920, n32612, n32190, n32541, n17665, 
            n4_adj_4, n32580, n2994, is_alu_reg_de, n2136, n32360, 
            is_jalr_de, is_lui_N_1365, is_lui_de, n32427, n26863, 
            n19_adj_5, n24898, n24900) /* synthesis syn_module_defined=1 */ ;
    input n32361;
    input n32623;
    output n32362;
    input is_jal_N_1374;
    input n32630;
    output is_jal_de;
    input n7;
    input n22;
    input n32653;
    output n32566;
    output n32340;
    input n32634;
    input n32637;
    input n32641;
    input n32651;
    input n29039;
    output \additional_mem_ops_2__N_1132[0] ;
    input n32654;
    input n32599;
    input n32659;
    input n32658;
    input n32661;
    input n32657;
    input n32638;
    input n32640;
    output n32582;
    input n32643;
    output n32576;
    input n7_adj_1;
    output n9;
    output n8330;
    output n8;
    output n29119;
    input n32642;
    input n32655;
    input n32656;
    input n32639;
    output n10;
    output n24;
    input n32594;
    input n2225;
    input n2156;
    output n29748;
    input n34287;
    output n28501;
    input \instr[16] ;
    output n2598;
    output n29605;
    output n32565;
    input \instr[20] ;
    input n32539;
    output n27731;
    output n28489;
    input rst_reg_n;
    input n10024;
    output n28575;
    output n29681;
    output is_load_de;
    input \instr[25] ;
    output n3355;
    output n672;
    output mem_op_increment_reg_de;
    output n32571;
    input n2157;
    output n29725;
    input n32540;
    input n32734;
    output n30041;
    output n32573;
    output n4251;
    output n32533;
    output \alu_op_3__N_1170[1] ;
    output n26937;
    output n27;
    input \instr[30] ;
    input n3;
    output n156;
    output n32563;
    input n41;
    output n30;
    output n22_adj_2;
    input n32629;
    input \alu_op_3__N_1337[2] ;
    input n32585;
    output n32;
    input n4257;
    output n3253;
    output n32176;
    input n32609;
    input n4259;
    output n3286;
    output n3288;
    output n32577;
    output n3290;
    output n3289;
    input n29025;
    output n28577;
    input n32615;
    input n32597;
    output n32222;
    output n9394;
    input \instr[29] ;
    input \instr[31] ;
    output n5207;
    input \instr[24] ;
    output n5212;
    output n5222;
    input \instr[19] ;
    output n32030;
    output n5221;
    input n2205;
    output n5224;
    input n29716;
    output n29705;
    input n32025;
    output n32024;
    input n29712;
    output n29695;
    input \instr[28] ;
    output n5208;
    output n5220;
    output n5211;
    input n29714;
    output n29697;
    input n32016;
    output n32017;
    output n29726;
    input n29718;
    output n29703;
    output n5223;
    output n29747;
    input n2153;
    output n29732;
    input n32583;
    output is_auipc_de;
    output n5231;
    output n32559;
    output n5236;
    output n5232;
    input n32569;
    input n32617;
    input n32618;
    output is_system_de;
    input n29211;
    output is_store_de;
    input \instr[26] ;
    input n32627;
    output is_alu_imm_de;
    input n32581;
    input n29031;
    input n32603;
    output n2986;
    output n331;
    input n32602;
    input n32596;
    output n11066;
    output n29723;
    output n32570;
    output n28919;
    input \instr[23] ;
    output n28791;
    input \instr[22] ;
    output n28763;
    input \instr[21] ;
    output n28805;
    output n28777;
    input n31698;
    input n32619;
    input n32633;
    output is_branch_de;
    input n32589;
    output \mem_op_de[2] ;
    input n28617;
    input n26;
    output n28623;
    input n28593;
    output n28599;
    input n4;
    output n28539;
    input n28653;
    output n28659;
    input n2798;
    input \instr[17] ;
    input n2592;
    output n2620;
    input n28561;
    output n28567;
    input n28641;
    output n28647;
    input n28547;
    output n28553;
    input n28605;
    output n28611;
    output n12;
    output n28527;
    input n28407;
    input n19;
    output n28413;
    input n26879;
    output n28669;
    output n19_adj_3;
    input n27959;
    output [3:0]alu_op_de;
    input n32613;
    output n28363;
    input n27788;
    input n9048;
    input n30919;
    input n32610;
    input n9052;
    input n30920;
    input n32612;
    output n32190;
    input n32541;
    input n17665;
    output n4_adj_4;
    output n32580;
    output n2994;
    output is_alu_reg_de;
    input n2136;
    output n32360;
    output is_jalr_de;
    input is_lui_N_1365;
    output is_lui_de;
    input n32427;
    input n26863;
    input n19_adj_5;
    input n24898;
    output n24900;
    
    
    wire n32359, alu_op_3__N_1181, n8246, n32339, n32334, n32303, 
        n32586;
    wire [3:0]alu_op_3__N_1170;
    
    wire n32426, mem_op_2__N_1384, n32593, n19_c, n32600, n18321, 
        n32512, n32511, n32587, n8528;
    wire [3:0]alu_op_3__N_1107;
    
    wire n31699, n27874, n32863, n30_c, n32579, n32567, alu_op_3__N_1180, 
        imm_31__N_1169, n32_c, n27915, n15, n24899, n24_adj_3158, 
        n15_adj_3159, n32862, is_jalr_N_1370, n32590, n31700, n18306, 
        n29746, n43, n24_adj_3160, n27_adj_3161, n29189, n27753, 
        n15_adj_3162, n32864, n32428, n8537;
    
    PFUMX i29207 (.BLUT(n32361), .ALUT(n32359), .C0(n32623), .Z(n32362));
    PFUMX is_jal_I_0 (.BLUT(is_jal_N_1374), .ALUT(alu_op_3__N_1181), .C0(n32630), 
          .Z(is_jal_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    PFUMX i5586 (.BLUT(n7), .ALUT(n22), .C0(n32653), .Z(n8246));
    PFUMX i29190 (.BLUT(n32339), .ALUT(n32334), .C0(n32566), .Z(n32340));
    PFUMX i29169 (.BLUT(n32634), .ALUT(n32303), .C0(n32586), .Z(alu_op_3__N_1170[2]));
    LUT4 additional_mem_ops_2__N_1132_0__bdd_3_lut (.A(n32637), .B(n32641), 
         .C(n32651), .Z(n32426)) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam additional_mem_ops_2__N_1132_0__bdd_3_lut.init = 16'h1515;
    LUT4 i585_4_lut (.A(n32651), .B(mem_op_2__N_1384), .C(n32593), .D(n29039), 
         .Z(\additional_mem_ops_2__N_1132[0] )) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(93[13] 98[16])
    defparam i585_4_lut.init = 16'h3733;
    LUT4 i15663_4_lut (.A(n19_c), .B(n32600), .C(n32654), .D(n32599), 
         .Z(n18321)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i15663_4_lut.init = 16'hcac0;
    LUT4 instr_5__bdd_4_lut (.A(n32659), .B(n32658), .C(n32661), .D(n32657), 
         .Z(n32512)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B ((D)+!C)+!B (C+(D)))) */ ;
    defparam instr_5__bdd_4_lut.init = 16'hffbc;
    LUT4 instr_5__bdd_3_lut (.A(n32659), .B(n32658), .C(n32661), .Z(n32511)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam instr_5__bdd_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_567_3_lut (.A(n32638), .B(n32640), .C(n32641), .Z(n32582)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_rep_567_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_561_3_lut_4_lut (.A(n32638), .B(n32640), .C(n32643), 
         .D(n32641), .Z(n32576)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_rep_561_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_3_lut_rep_572_4_lut (.A(n32638), .B(n32640), .C(n32637), .D(n32641), 
         .Z(n32587)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_3_lut_rep_572_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_578_3_lut (.A(n32658), .B(n32657), .C(n32661), .Z(n32593)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(72[27:51])
    defparam i1_2_lut_rep_578_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32658), .B(n32657), .C(n7_adj_1), .D(n32661), 
         .Z(n9)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(72[27:51])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_360 (.A(n32658), .B(n32657), .C(n8330), 
         .D(n8), .Z(n29119)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(72[27:51])
    defparam i1_2_lut_3_lut_4_lut_adj_360.init = 16'hf0e0;
    LUT4 i15037_4_lut (.A(n32642), .B(n8330), .C(n32655), .D(n8528), 
         .Z(alu_op_3__N_1107[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[18] 85[91])
    defparam i15037_4_lut.init = 16'hc088;
    LUT4 i28260_3_lut_rep_585_4_lut (.A(n32658), .B(n32657), .C(n7_adj_1), 
         .D(n32661), .Z(n32600)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(72[27:51])
    defparam i28260_3_lut_rep_585_4_lut.init = 16'h0100;
    LUT4 instr_6__I_0_157_i9_2_lut_rep_571_3_lut (.A(n32658), .B(n32657), 
         .C(n8), .Z(n32586)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(72[27:51])
    defparam instr_6__I_0_157_i9_2_lut_rep_571_3_lut.init = 16'hfefe;
    LUT4 is_jalr_N_1372_bdd_2_lut_29267_3_lut (.A(n32656), .B(n32639), .C(n32655), 
         .Z(n31699)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam is_jalr_N_1372_bdd_2_lut_29267_3_lut.init = 16'h7070;
    LUT4 n8208_bdd_2_lut_3_lut_3_lut_4_lut (.A(n32656), .B(n32639), .C(n32655), 
         .D(n32630), .Z(n32359)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n8208_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i2_2_lut_3_lut (.A(n32656), .B(n32639), .C(n32655), .Z(n10)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h8080;
    LUT4 i37_3_lut_3_lut (.A(n32656), .B(n32639), .C(n32655), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;
    defparam i37_3_lut_3_lut.init = 16'h7a7a;
    LUT4 i1_3_lut (.A(n8330), .B(alu_op_3__N_1170[2]), .C(n32654), .Z(n27874)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i29188_then_4_lut (.A(n32656), .B(n32594), .C(n2225), .D(\additional_mem_ops_2__N_1132[0] ), 
         .Z(n32863)) /* synthesis lut_function=(A (B (C)+!B !(C+(D)))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam i29188_then_4_lut.init = 16'hc0c7;
    LUT4 i15622_2_lut_3_lut_4_lut (.A(n32639), .B(n32655), .C(n32656), 
         .D(n32654), .Z(n30_c)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i15622_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 mux_1526_i12_rep_129_3_lut_3_lut_4_lut (.A(n32654), .B(n32653), 
         .C(n2156), .D(n32643), .Z(n29748)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1526_i12_rep_129_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut (.A(n32654), .B(n32653), .C(n34287), .Z(n28501)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_361 (.A(n32654), .B(n32653), .C(\instr[16] ), 
         .Z(n2598)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_361.init = 16'h8080;
    LUT4 i26964_2_lut_3_lut (.A(n32654), .B(n32653), .C(n32656), .Z(n29605)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i26964_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i169_2_lut_rep_550_2_lut_3_lut (.A(n32654), .B(n32653), .C(n32655), 
         .Z(n32565)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i169_2_lut_rep_550_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_3_lut_3_lut_4_lut (.A(n32654), .B(n32653), .C(\instr[20] ), 
         .D(n32539), .Z(n27731)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n32654), .B(n32653), .C(n32643), 
         .D(n32587), .Z(n28489)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h7770;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_adj_362 (.A(n32654), .B(n32653), .C(rst_reg_n), 
         .D(n10024), .Z(n28575)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut_adj_362.init = 16'h0070;
    LUT4 is_load_I_0_4_lut_4_lut (.A(n32654), .B(n32653), .C(n29681), 
         .D(n8246), .Z(is_load_de)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(D))) */ ;
    defparam is_load_I_0_4_lut_4_lut.init = 16'h5d08;
    LUT4 i6608_3_lut_4_lut (.A(n32654), .B(n32653), .C(\instr[25] ), .D(n32642), 
         .Z(n3355)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i6608_3_lut_4_lut.init = 16'hf780;
    LUT4 n8208_bdd_2_lut_29206_2_lut_3_lut (.A(n32654), .B(n32653), .C(n32656), 
         .Z(n32334)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam n8208_bdd_2_lut_29206_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i1_2_lut_2_lut_3_lut (.A(n32654), .B(n32653), .C(n32656), .Z(n672)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'h7070;
    LUT4 i15045_2_lut_2_lut_3_lut (.A(n32654), .B(n32653), .C(mem_op_2__N_1384), 
         .Z(mem_op_increment_reg_de)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i15045_2_lut_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_556_2_lut_3_lut (.A(n32654), .B(n32653), .C(n34287), 
         .Z(n32571)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_rep_556_2_lut_3_lut.init = 16'h7070;
    LUT4 mux_1526_i11_rep_106_3_lut_3_lut_4_lut (.A(n32654), .B(n32653), 
         .C(n2157), .D(n32638), .Z(n29725)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1526_i11_rep_106_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 i28602_2_lut_3_lut_4_lut (.A(n32654), .B(n32653), .C(n32540), 
         .D(n32734), .Z(n30041)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;
    defparam i28602_2_lut_3_lut_4_lut.init = 16'hf0f8;
    LUT4 i5548_2_lut_rep_558_2_lut_3_lut_4_lut (.A(n32654), .B(n32653), 
         .C(n32655), .D(n32656), .Z(n32573)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;
    defparam i5548_2_lut_rep_558_2_lut_3_lut_4_lut.init = 16'h7770;
    LUT4 i6606_rep_518_4_lut (.A(n32654), .B(n32653), .C(n32539), .D(n4251), 
         .Z(n32533)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam i6606_rep_518_4_lut.init = 16'h08f8;
    LUT4 mux_29_i2_4_lut (.A(n32656), .B(n32579), .C(n32586), .D(n32655), 
         .Z(\alu_op_3__N_1170[1] )) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[18] 85[91])
    defparam mux_29_i2_4_lut.init = 16'hfaca;
    LUT4 i167_2_lut_rep_551_2_lut_3_lut (.A(n32654), .B(n32653), .C(n32639), 
         .Z(n32566)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i167_2_lut_rep_551_2_lut_3_lut.init = 16'h7070;
    LUT4 instr_6__I_0_142_i10_2_lut_3_lut (.A(n32657), .B(n32658), .C(n8), 
         .Z(alu_op_3__N_1181)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam instr_6__I_0_142_i10_2_lut_3_lut.init = 16'h0808;
    LUT4 i1_3_lut_adj_363 (.A(n32651), .B(n32642), .C(n32659), .Z(n26937)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam i1_3_lut_adj_363.init = 16'hfefe;
    LUT4 i42_4_lut_4_lut_4_lut (.A(n32655), .B(n32656), .C(n32654), .D(n32653), 
         .Z(n27)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i42_4_lut_4_lut_4_lut.init = 16'h404a;
    LUT4 i14978_4_lut (.A(\instr[30] ), .B(n32579), .C(n32659), .D(n3), 
         .Z(n156)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(85[18:91])
    defparam i14978_4_lut.init = 16'hecee;
    LUT4 i24422_2_lut_rep_548_3_lut_4_lut_4_lut (.A(n32658), .B(n32661), 
         .C(n32651), .D(n32657), .Z(n32563)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam i24422_2_lut_rep_548_3_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_rep_552_3_lut_3_lut (.A(n32658), .B(n32661), .C(n32657), 
         .Z(n32567)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam i1_2_lut_rep_552_3_lut_3_lut.init = 16'hf7f7;
    LUT4 instr_6__I_0_130_i10_2_lut_3_lut_3_lut (.A(n32658), .B(n8), .C(n32657), 
         .Z(alu_op_3__N_1180)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam instr_6__I_0_130_i10_2_lut_3_lut_3_lut.init = 16'h0202;
    LUT4 instr_6__I_0_127_i10_2_lut_3_lut_4_lut_4_lut (.A(n32658), .B(n32661), 
         .C(n7_adj_1), .D(n32657), .Z(imm_31__N_1169)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam instr_6__I_0_127_i10_2_lut_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n32655), .B(n41), .C(n32_c), .D(n32654), 
         .Z(n30)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h00dc;
    LUT4 i1_4_lut_4_lut_4_lut_adj_364 (.A(n32655), .B(n27915), .C(n32654), 
         .D(n32653), .Z(n22_adj_2)) /* synthesis lut_function=(!(A+(B (C (D))+!B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i1_4_lut_4_lut_4_lut_adj_364.init = 16'h0454;
    LUT4 i15528_4_lut_4_lut (.A(n32655), .B(n32656), .C(n32629), .D(\alu_op_3__N_1337[2] ), 
         .Z(n15)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i15528_4_lut_4_lut.init = 16'hd0c0;
    LUT4 i53_4_lut_4_lut (.A(n32655), .B(n32653), .C(n32585), .D(n32654), 
         .Z(n32)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i53_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_2079_i2_4_lut_4_lut (.A(n32655), .B(n4257), .C(n32657), .D(n32659), 
         .Z(n3253)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam mux_2079_i2_4_lut_4_lut.init = 16'h7340;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n32656), .B(n32655), .C(n32640), 
         .D(n32639), .Z(n24899)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam i1_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 n10904_bdd_2_lut_29106_3_lut_4_lut_4_lut_4_lut (.A(n32656), .B(n32655), 
         .C(n32643), .D(n32639), .Z(n32176)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam n10904_bdd_2_lut_29106_3_lut_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(n32656), .B(n32609), .C(n32593), 
         .D(n32639), .Z(n32_c)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h54ff;
    LUT4 mux_2084_i6_4_lut_4_lut (.A(n32656), .B(n4259), .C(n32639), .D(n32658), 
         .Z(n3286)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam mux_2084_i6_4_lut_4_lut.init = 16'hddc0;
    LUT4 mux_2084_i4_4_lut_4_lut (.A(n32656), .B(n4259), .C(n32639), .D(n32659), 
         .Z(n3288)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam mux_2084_i4_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i1_2_lut_rep_562_3_lut_3_lut_3_lut (.A(n32656), .B(n32655), .C(n32639), 
         .Z(n32577)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam i1_2_lut_rep_562_3_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 mux_2084_i2_4_lut_4_lut (.A(n32656), .B(n4259), .C(n32639), .D(n32657), 
         .Z(n3290)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam mux_2084_i2_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_2084_i3_4_lut_4_lut (.A(n32656), .B(n4259), .C(n32639), .D(n32661), 
         .Z(n3289)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam mux_2084_i3_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i1_4_lut_4_lut (.A(n32656), .B(n24_adj_3158), .C(n28575), .D(n29025), 
         .Z(n28577)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam i1_4_lut_4_lut.init = 16'hf040;
    LUT4 i15_2_lut_3_lut_4_lut_4_lut (.A(n32656), .B(n32643), .C(n32641), 
         .D(n32615), .Z(n15_adj_3159)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam i15_2_lut_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 n8539_bdd_3_lut_4_lut_4_lut (.A(n32656), .B(n32638), .C(n32643), 
         .D(n32597), .Z(n32222)) /* synthesis lut_function=(A+!(B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[49:59])
    defparam n8539_bdd_3_lut_4_lut_4_lut.init = 16'habff;
    LUT4 i6713_3_lut_4_lut (.A(n32567), .B(n32651), .C(n32540), .D(n32630), 
         .Z(n9394)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i6713_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_3151_i30_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[29] ), 
         .D(\instr[31] ), .Z(n5207)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_3151_i30_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_3151_i25_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[24] ), 
         .D(\instr[31] ), .Z(n5212)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_3151_i25_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_3151_i15_3_lut_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n32656), .Z(n5222)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3151_i15_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n4263_bdd_3_lut_29025_4_lut (.A(n32567), .B(n32651), .C(\instr[19] ), 
         .D(\instr[31] ), .Z(n32030)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam n4263_bdd_3_lut_29025_4_lut.init = 16'hfe10;
    LUT4 mux_3151_i16_3_lut_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n32639), .Z(n5221)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3151_i16_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i29188_else_4_lut (.A(n2205), .B(n32656), .C(n32594), .D(\additional_mem_ops_2__N_1132[0] ), 
         .Z(n32862)) /* synthesis lut_function=(A (C)+!A !(B (C+(D))+!B (D))) */ ;
    defparam i29188_else_4_lut.init = 16'ha0b5;
    LUT4 mux_3151_i13_3_lut_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n32642), .Z(n5224)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3151_i13_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1526_i7_rep_86_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n29716), .Z(n29705)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1526_i7_rep_86_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32023_bdd_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n32025), .Z(n32024)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam n32023_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1526_i5_rep_76_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n29712), .Z(n29695)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1526_i5_rep_76_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_3151_i29_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[28] ), 
         .D(\instr[31] ), .Z(n5208)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_3151_i29_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_3151_i17_3_lut_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(\instr[16] ), .Z(n5220)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3151_i17_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_3151_i26_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[25] ), 
         .D(\instr[31] ), .Z(n5211)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_3151_i26_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_1526_i6_rep_78_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n29714), .Z(n29697)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1526_i6_rep_78_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n32016_bdd_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n32016), .Z(n32017)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam n32016_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1526_i11_rep_107_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n2157), .Z(n29726)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1526_i11_rep_107_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1526_i8_rep_84_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n29718), .Z(n29703)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1526_i8_rep_84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_3151_i14_3_lut_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n32655), .Z(n5223)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3151_i14_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_365 (.A(n32651), .B(n32659), .C(n32661), .Z(n8)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_adj_365.init = 16'hf7f7;
    LUT4 mux_1526_i12_rep_128_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n2156), .Z(n29747)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1526_i12_rep_128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1526_i15_rep_113_3_lut_4_lut (.A(n32567), .B(n32651), .C(\instr[31] ), 
         .D(n2153), .Z(n29732)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1526_i15_rep_113_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut (.A(n32661), .B(n32583), .C(n32630), .D(n32609), 
         .Z(is_auipc_de)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i1_3_lut_4_lut.init = 16'h0020;
    LUT4 i15483_2_lut_3_lut_4_lut (.A(n32661), .B(n32583), .C(\instr[25] ), 
         .D(n32651), .Z(n5231)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i15483_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i15104_2_lut_rep_544_3_lut_4_lut (.A(n32661), .B(n32583), .C(n9), 
         .D(n32651), .Z(n32559)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i15104_2_lut_rep_544_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i15249_2_lut_3_lut_4_lut (.A(n32661), .B(n32583), .C(n32638), 
         .D(n32651), .Z(n5236)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i15249_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i15482_2_lut_3_lut_4_lut (.A(n32661), .B(n32583), .C(n32637), 
         .D(n32651), .Z(n5232)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i15482_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i1_3_lut_4_lut_adj_366 (.A(n32643), .B(n32587), .C(n32653), .D(n29681), 
         .Z(n27915)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_3_lut_4_lut_adj_366.init = 16'h00e0;
    LUT4 i1_3_lut_4_lut_adj_367 (.A(n32643), .B(n32587), .C(n32569), .D(n32617), 
         .Z(is_jalr_N_1370)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_3_lut_4_lut_adj_367.init = 16'he000;
    LUT4 n31700_bdd_3_lut_4_lut (.A(n32590), .B(n32618), .C(n32654), .D(n31700), 
         .Z(is_system_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam n31700_bdd_3_lut_4_lut.init = 16'h2f20;
    LUT4 is_store_I_0_4_lut (.A(n29211), .B(n9), .C(n32630), .D(n18306), 
         .Z(is_store_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam is_store_I_0_4_lut.init = 16'h3a30;
    LUT4 i15651_4_lut (.A(n32653), .B(n32656), .C(n32655), .D(n32637), 
         .Z(n18306)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i15651_4_lut.init = 16'hcdcc;
    LUT4 mux_1526_i12_rep_127_3_lut_4_lut (.A(\instr[26] ), .B(n32600), 
         .C(n32656), .D(n2156), .Z(n29746)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[22:45])
    defparam mux_1526_i12_rep_127_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_4_lut (.A(n32627), .B(n32654), .C(n43), .D(n24_adj_3160), 
         .Z(is_alu_imm_de)) /* synthesis lut_function=(A (B (D))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i1_4_lut.init = 16'hcd05;
    LUT4 i44_3_lut (.A(n32656), .B(n32653), .C(n32654), .Z(n43)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i44_3_lut.init = 16'hcaca;
    LUT4 i45_4_lut (.A(n27_adj_3161), .B(n29189), .C(n32653), .D(n32618), 
         .Z(n24_adj_3160)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i45_4_lut.init = 16'h0aca;
    LUT4 i1_4_lut_4_lut_adj_368 (.A(n32581), .B(n32637), .C(n32641), .D(n26937), 
         .Z(n27753)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i1_4_lut_4_lut_adj_368.init = 16'h1050;
    LUT4 i1_4_lut_adj_369 (.A(n32655), .B(n7_adj_1), .C(n32656), .D(n29031), 
         .Z(mem_op_2__N_1384)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_369.init = 16'hffdf;
    LUT4 mux_2051_i17_3_lut_4_lut (.A(n32657), .B(n32603), .C(n32639), 
         .D(n32642), .Z(n2986)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_2051_i17_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_61_i2_3_lut_4_lut (.A(n32657), .B(n32603), .C(n32642), .D(n32651), 
         .Z(n331)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_61_i2_3_lut_4_lut.init = 16'hbfb0;
    LUT4 i15637_2_lut_4_lut (.A(n32639), .B(n32654), .C(n32602), .D(n32596), 
         .Z(n15_adj_3162)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i15637_2_lut_4_lut.init = 16'h0008;
    LUT4 i8365_3_lut_4_lut (.A(n32615), .B(n32641), .C(n32643), .D(n32656), 
         .Z(n11066)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i8365_3_lut_4_lut.init = 16'h10f0;
    PFUMX i29309 (.BLUT(n32862), .ALUT(n32863), .C0(n32734), .Z(n32864));
    LUT4 mux_2051_i16_rep_103_3_lut_4_lut (.A(n32657), .B(n32603), .C(n32639), 
         .D(n32642), .Z(n29723)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(205[25] 214[32])
    defparam mux_2051_i16_rep_103_3_lut_4_lut.init = 16'hefe0;
    LUT4 i5866_2_lut_3_lut_4_lut (.A(n32618), .B(n8), .C(n32600), .D(\instr[26] ), 
         .Z(n8528)) /* synthesis lut_function=(A (C (D))+!A ((C (D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam i5866_2_lut_3_lut_4_lut.init = 16'hf111;
    LUT4 i1_2_lut_rep_555_4_lut (.A(n32641), .B(n32615), .C(n32637), .D(n32643), 
         .Z(n32570)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_rep_555_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(n32641), .B(n32615), .C(n32637), .D(n32643), 
         .Z(n28919)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_4_lut.init = 16'h00fe;
    LUT4 i1_3_lut_4_lut_adj_370 (.A(n32617), .B(n32623), .C(n34287), .D(\instr[23] ), 
         .Z(n28791)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_370.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_adj_371 (.A(n32617), .B(n32623), .C(rst_reg_n), 
         .D(\instr[22] ), .Z(n28763)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_371.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_adj_372 (.A(n32617), .B(n32623), .C(n34287), .D(\instr[21] ), 
         .Z(n28805)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_372.init = 16'h1000;
    LUT4 i1_3_lut_4_lut_adj_373 (.A(n32617), .B(n32623), .C(n34287), .D(\instr[20] ), 
         .Z(n28777)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_373.init = 16'h1000;
    PFUMX i28840 (.BLUT(n31699), .ALUT(n31698), .C0(n32653), .Z(n31700));
    LUT4 is_branch_I_0_4_lut (.A(n32619), .B(n32586), .C(n32630), .D(n32633), 
         .Z(is_branch_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam is_branch_I_0_4_lut.init = 16'h3a30;
    LUT4 i14954_2_lut_3_lut_4_lut (.A(n32661), .B(n32618), .C(n32655), 
         .D(n32609), .Z(n19_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam i14954_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n32630), .B(n32428), .C(n32589), .D(n32602), 
         .Z(\mem_op_de[2] )) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C+(D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h080c;
    LUT4 i1_4_lut_4_lut_adj_374 (.A(n32630), .B(n28617), .C(n10024), .D(n26), 
         .Z(n28623)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_374.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_375 (.A(n32630), .B(n28593), .C(n10024), .D(n26), 
         .Z(n28599)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_375.init = 16'h0400;
    LUT4 i1_3_lut_4_lut_4_lut_adj_376 (.A(n32630), .B(n10024), .C(n4), 
         .D(n34287), .Z(n28539)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_376.init = 16'h1000;
    LUT4 n32338_bdd_3_lut_3_lut_4_lut_4_lut (.A(n32630), .B(n32617), .C(n32864), 
         .D(n32602), .Z(n32339)) /* synthesis lut_function=(A (B+(C))+!A !(B (D)+!B !(C))) */ ;
    defparam n32338_bdd_3_lut_3_lut_4_lut_4_lut.init = 16'hb8fc;
    LUT4 i1_4_lut_4_lut_adj_377 (.A(n32630), .B(n28653), .C(n10024), .D(n26), 
         .Z(n28659)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_377.init = 16'h0400;
    LUT4 mux_1867_i3_4_lut_4_lut (.A(n32630), .B(n2798), .C(\instr[17] ), 
         .D(n2592), .Z(n2620)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;
    defparam mux_1867_i3_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i1_4_lut_4_lut_adj_378 (.A(n32630), .B(n28561), .C(n10024), .D(n26), 
         .Z(n28567)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_378.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_379 (.A(n32630), .B(n28641), .C(n10024), .D(n26), 
         .Z(n28647)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_379.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_380 (.A(n32630), .B(n28547), .C(n10024), .D(n26), 
         .Z(n28553)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_380.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_381 (.A(n32630), .B(n28605), .C(n10024), .D(n26), 
         .Z(n28611)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_381.init = 16'h0400;
    LUT4 i2_2_lut_3_lut_4_lut_4_lut (.A(n32630), .B(n32602), .C(n32593), 
         .D(n32609), .Z(n12)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i2_2_lut_3_lut_4_lut_4_lut.init = 16'hfff4;
    LUT4 i1_3_lut_4_lut_4_lut_adj_382 (.A(n32630), .B(n32623), .C(n32617), 
         .D(n32639), .Z(n28527)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_382.init = 16'h1000;
    LUT4 i1_4_lut_4_lut_adj_383 (.A(n32630), .B(n28407), .C(n10024), .D(n19), 
         .Z(n28413)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_383.init = 16'h0400;
    LUT4 instr_2__bdd_4_lut (.A(n32658), .B(n26879), .C(n32651), .D(n32657), 
         .Z(n4251)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam instr_2__bdd_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_384 (.A(n32630), .B(n34287), .C(n32642), .D(n10024), 
         .Z(n28669)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_384.init = 16'h0040;
    LUT4 i1_3_lut_4_lut_4_lut_adj_385 (.A(n32630), .B(n32623), .C(n32637), 
         .D(n32655), .Z(n19_adj_3)) /* synthesis lut_function=(A (B+(C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_385.init = 16'ha8fc;
    LUT4 i5876_4_lut (.A(n27959), .B(n8537), .C(n32653), .D(n32581), 
         .Z(alu_op_de[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i5876_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_4_lut_adj_386 (.A(n32630), .B(n32613), .C(n32633), .D(n10024), 
         .Z(n28363)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_4_lut_adj_386.init = 16'h0010;
    PFUMX i6368 (.BLUT(n27788), .ALUT(n9048), .C0(n32653), .Z(alu_op_de[1]));
    PFUMX i6370 (.BLUT(n15), .ALUT(n27874), .C0(n30919), .Z(alu_op_de[2]));
    PFUMX i5875 (.BLUT(alu_op_3__N_1107[0]), .ALUT(n30_c), .C0(n32610), 
          .Z(n8537));
    PFUMX i6372 (.BLUT(n27753), .ALUT(n9052), .C0(n30920), .Z(alu_op_de[3]));
    LUT4 i25_2_lut_rep_564_4_lut (.A(n32661), .B(n7_adj_1), .C(n32618), 
         .D(\instr[26] ), .Z(n32579)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(67[27:51])
    defparam i25_2_lut_rep_564_4_lut.init = 16'h0200;
    PFUMX i29303 (.BLUT(n32512), .ALUT(n32511), .C0(n32651), .Z(n8330));
    LUT4 n10904_bdd_3_lut_4_lut (.A(n32639), .B(n32612), .C(n32654), .D(n32658), 
         .Z(n32190)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam n10904_bdd_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_4_lut_adj_387 (.A(n32630), .B(n32541), .C(n17665), .D(n32639), 
         .Z(n4_adj_4)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_4_lut_adj_387.init = 16'h0444;
    LUT4 i28430_2_lut_rep_565_3_lut (.A(n32661), .B(n32658), .C(n32657), 
         .Z(n32580)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i28430_2_lut_rep_565_3_lut.init = 16'h0808;
    LUT4 mux_2051_i9_3_lut_4_lut_4_lut (.A(n32661), .B(n32658), .C(n32639), 
         .D(n32657), .Z(n2994)) /* synthesis lut_function=(A (B+((D)+!C))+!A (C (D))) */ ;
    defparam mux_2051_i9_3_lut_4_lut_4_lut.init = 16'hfa8a;
    PFUMX i15664 (.BLUT(n15_adj_3162), .ALUT(n18321), .C0(n30919), .Z(is_alu_reg_de));
    LUT4 i1_3_lut_rep_575_4_lut (.A(n32659), .B(n32651), .C(n32661), .D(n32653), 
         .Z(n32590)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(218[25] 223[32])
    defparam i1_3_lut_rep_575_4_lut.init = 16'h8000;
    LUT4 n2136_bdd_4_lut (.A(n2136), .B(n32734), .C(n32579), .D(n29746), 
         .Z(n32303)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam n2136_bdd_4_lut.init = 16'hef20;
    LUT4 n8208_bdd_4_lut_29246 (.A(\additional_mem_ops_2__N_1132[0] ), .B(n32566), 
         .C(n32642), .D(n32641), .Z(n32360)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam n8208_bdd_4_lut_29246.init = 16'hdc10;
    LUT4 i27036_3_lut_4_lut (.A(n32659), .B(n32651), .C(n32661), .D(n32618), 
         .Z(n29681)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam i27036_3_lut_4_lut.init = 16'hfffe;
    PFUMX is_jalr_I_0 (.BLUT(is_jalr_N_1370), .ALUT(alu_op_3__N_1180), .C0(n32630), 
          .Z(is_jalr_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    PFUMX is_lui_I_0 (.BLUT(is_lui_N_1365), .ALUT(imm_31__N_1169), .C0(n32630), 
          .Z(is_lui_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 i1_2_lut_3_lut_adj_388 (.A(n32659), .B(n32651), .C(n32661), .Z(n29189)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam i1_2_lut_3_lut_adj_388.init = 16'h1010;
    PFUMX i29244 (.BLUT(n32427), .ALUT(n32426), .C0(n32566), .Z(n32428));
    LUT4 i43_4_lut_3_lut (.A(n32653), .B(n26863), .C(n32655), .Z(n24_adj_3158)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i43_4_lut_3_lut.init = 16'h5858;
    PFUMX i43 (.BLUT(n15_adj_3159), .ALUT(n19_adj_5), .C0(n32639), .Z(n27_adj_3161));
    PFUMX i22327 (.BLUT(n24898), .ALUT(n24899), .C0(n30920), .Z(n24900));
    
endmodule
//
// Verilog Description of module tinyqv_core
//

module tinyqv_core (\imm[6] , clk_c, n32840, mip_reg, clk_c_enable_342, 
            n32650, n32351, counter_hi, \imm[10] , \imm[0] , n32759, 
            \imm[2] , \debug_branch_N_450[1] , n5660, n5661, n30329, 
            n32309, instr_complete_N_1647, clk_c_enable_285, cycle, 
            \alu_op[0] , \alu_op[1] , is_system, debug_instr_valid, 
            n32702, n32733, n32704, n32746, \ui_in_sync[1] , n24384, 
            stall_core, n32774, n32545, is_load, n829, n26962, clk_c_enable_533, 
            \alu_op_in[2] , \ui_in_sync[0] , debug_rd, \mie[10] , \mie[14] , 
            \mie[2] , \mie[6] , n27294, n5017, n1766, \instr_write_offset_3__N_934[1] , 
            n1767, \instr_write_offset_3__N_934[0] , n1768, pc_2__N_932, 
            \next_pc_for_core[15] , \next_pc_for_core[11] , n32846, n32847, 
            \imm[7] , n9058, n29689, n32691, n32549, n32543, instr_fetch_running, 
            was_early_branch, n32550, n32564, data_ready_sync, data_ready_core, 
            n131, n32768, n32849, n32697, clk_c_enable_538, \imm[1] , 
            n32838, n29866, clk_c_enable_433, n32854, interrupt_core, 
            rst_reg_n, n17920, n28685, n28687, n34285, is_lui, is_jal, 
            is_branch, is_jalr, is_auipc, n34281, n32551, mstatus_mte, 
            n92, n34287, n27003, n32821, mem_op, n32741, \alu_op[3] , 
            accum, d_3__N_1868, data_out_3__N_1385, is_timer_addr, n30160, 
            n32784, n32677, debug_rd_3__N_1575, \imm[11] , clk_c_enable_276, 
            fsm_state, n32791, n32763, n32730, timer_interrupt, n32765, 
            n5642, n926, n33057, \timer_data[0] , clk_c_enable_321, 
            n893, load_done, clk_c_enable_363, n8228, n32317, \timer_data[2] , 
            data_rs1, n860, n793, n32546, n28417, n32580, n32642, 
            n3274, n28429, n4, n27546, n28465, n27541, \debug_branch_N_450[3] , 
            load_top_bit, n32806, n32808, instr_complete_N_1651, instr_complete_N_1652, 
            is_double_fault_r, n28441, n27545, n32732, n8, n5659, 
            debug_rd_3__N_413, n28275, n1, n27427, \imm[4] , n5607, 
            \cycle_count_wide[3] , n28343, n32559, n32539, data_rs2, 
            \data_out_slice[0] , n32644, n34283, timer_data_3__N_631, 
            \mtimecmp[7] , mtimecmp_3__N_1935, \data_rs1[3] , mstatus_mie_N_1709, 
            \data_rs1[0] , \imm[9] , \imm[8] , \addr_out[27] , \addr_out[24] , 
            \addr_out[25] , \addr_out[26] , n32829, \imm[5] , \imm[3] , 
            n27656, n28909, n27655, n29838, n30172, n27657, n28533, 
            n32548, clk_c_enable_524, n2559, n32834, n32760, n32758, 
            clk_c_enable_187, n28363, n28483, n32538, n32828, address_ready, 
            is_store, mstatus_mie_N_1707, n32710, n30425, n13, n29760, 
            n32668, \mtimecmp[5] , mtimecmp_1__N_1941, \debug_rd_3__N_405[28] , 
            n32848, n29844, n32678, n32675, is_alu_imm, is_alu_reg, 
            n28889, n27653, n31351, n29864, clk_c_enable_195, n18, 
            n29317, n32647, n32670, clk_c_enable_28, n32552, n32783, 
            n30928, n30927, n30926, n30925, n30924, n32769, \debug_branch_N_442[31] , 
            \debug_branch_N_442[30] , \debug_rd_3__N_405[30] , \debug_branch_N_442[29] , 
            \addr_offset[2] , n28963, \debug_rd_3__N_405[29] , n157, 
            \debug_branch_N_442[28] , n28495, n2124, \debug_rd_3__N_405[31] , 
            n701, \data_out_slice[2] , debug_early_branch_N_955, no_write_in_progress, 
            n1152, \next_pc_offset[3] , n28237, \debug_branch_N_450[0] , 
            n18098, \debug_branch_N_446[28] , n238, n30070, n76, \mtime_out[0] , 
            n32717, cy, n32663, n9620, time_pulse_r, n10737, n32680, 
            \next_pc_for_core[7] , \next_pc_for_core[3] , \next_pc_for_core[23] , 
            \next_pc_for_core[19] , \addr_out[1] , \addr_out[0] , n32690, 
            \addr_out[23] , \addr_out[22] , \addr_out[21] , \addr_out[20] , 
            \addr_out[19] , \addr_out[18] , \addr_out[17] , \addr_out[16] , 
            \addr_out[15] , \addr_out[14] , \addr_out[13] , \addr_out[12] , 
            \addr_out[11] , \addr_out[10] , \addr_out[9] , \addr_out[8] , 
            \addr_out[7] , \addr_out[6] , \addr_out[5] , \addr_out[4] , 
            \addr_out[3] , \mem_data_from_read[17] , \mem_data_from_read[21] , 
            n32308, \timer_data[1] , \mul_out[3] , \mul_out[2] , rd, 
            n32776, \mul_out[1] , \debug_branch_N_446[31] , n30175, 
            n29842, \debug_branch_N_446[30] , \csr_read_3__N_1447[2] , 
            n29836, \debug_branch_N_446[29] , n32767, \next_accum[5] , 
            GND_net, VCC_net, \next_accum[16] , \next_accum[17] , \next_accum[18] , 
            \next_accum[19] , \next_accum[6] , \next_accum[7] , \next_accum[8] , 
            \next_accum[9] , \next_accum[10] , \next_accum[11] , \next_accum[12] , 
            \next_accum[13] , \next_accum[14] , \next_accum[15] , \next_accum[4] , 
            n21667, rs1, rs2, \reg_access[3][2] , return_addr, \reg_access[4][3] , 
            n32652) /* synthesis syn_module_defined=1 */ ;
    input \imm[6] ;
    input clk_c;
    input n32840;
    output [17:16]mip_reg;
    input clk_c_enable_342;
    input n32650;
    output n32351;
    input [4:2]counter_hi;
    input \imm[10] ;
    input \imm[0] ;
    output n32759;
    input \imm[2] ;
    input \debug_branch_N_450[1] ;
    output n5660;
    output n5661;
    input n30329;
    input n32309;
    output instr_complete_N_1647;
    output clk_c_enable_285;
    output [1:0]cycle;
    input \alu_op[0] ;
    input \alu_op[1] ;
    input is_system;
    input debug_instr_valid;
    output n32702;
    output n32733;
    output n32704;
    output n32746;
    input \ui_in_sync[1] ;
    input n24384;
    input stall_core;
    output n32774;
    output n32545;
    input is_load;
    output n829;
    input n26962;
    output clk_c_enable_533;
    input \alu_op_in[2] ;
    input \ui_in_sync[0] ;
    output [3:0]debug_rd;
    output \mie[10] ;
    output \mie[14] ;
    output \mie[2] ;
    output \mie[6] ;
    output n27294;
    input [1:0]n5017;
    input n1766;
    output \instr_write_offset_3__N_934[1] ;
    input n1767;
    output \instr_write_offset_3__N_934[0] ;
    input [1:0]n1768;
    output [1:0]pc_2__N_932;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[11] ;
    input n32846;
    output n32847;
    input \imm[7] ;
    output n9058;
    input n29689;
    output n32691;
    output n32549;
    output n32543;
    input instr_fetch_running;
    input was_early_branch;
    output n32550;
    input n32564;
    input data_ready_sync;
    output data_ready_core;
    input n131;
    input n32768;
    output n32849;
    output n32697;
    output clk_c_enable_538;
    input \imm[1] ;
    input n32838;
    input n29866;
    input clk_c_enable_433;
    output n32854;
    input interrupt_core;
    input rst_reg_n;
    output n17920;
    input n28685;
    output n28687;
    input n34285;
    input is_lui;
    input is_jal;
    input is_branch;
    input is_jalr;
    input is_auipc;
    input n34281;
    output n32551;
    output mstatus_mte;
    input [3:0]n92;
    input n34287;
    output n27003;
    input n32821;
    input [2:0]mem_op;
    output n32741;
    input \alu_op[3] ;
    output [15:0]accum;
    output [19:0]d_3__N_1868;
    output data_out_3__N_1385;
    input is_timer_addr;
    input n30160;
    output n32784;
    output n32677;
    input debug_rd_3__N_1575;
    input \imm[11] ;
    input clk_c_enable_276;
    input [3:0]fsm_state;
    output n32791;
    output n32763;
    output n32730;
    input timer_interrupt;
    output n32765;
    input n5642;
    input n926;
    input n33057;
    input \timer_data[0] ;
    input clk_c_enable_321;
    input n893;
    output load_done;
    output clk_c_enable_363;
    input n8228;
    input n32317;
    input \timer_data[2] ;
    output [3:0]data_rs1;
    input n860;
    input n793;
    output n32546;
    input n28417;
    input n32580;
    input n32642;
    output n3274;
    input n28429;
    input n4;
    output n27546;
    input n28465;
    output n27541;
    input \debug_branch_N_450[3] ;
    output load_top_bit;
    output n32806;
    input n32808;
    input instr_complete_N_1651;
    input instr_complete_N_1652;
    output is_double_fault_r;
    input n28441;
    output n27545;
    output n32732;
    output n8;
    output n5659;
    input debug_rd_3__N_413;
    input n28275;
    input n1;
    output n27427;
    input \imm[4] ;
    output n5607;
    output \cycle_count_wide[3] ;
    input n28343;
    input n32559;
    output n32539;
    output [3:0]data_rs2;
    output \data_out_slice[0] ;
    output n32644;
    input n34283;
    input timer_data_3__N_631;
    input \mtimecmp[7] ;
    output mtimecmp_3__N_1935;
    output \data_rs1[3] ;
    output mstatus_mie_N_1709;
    output \data_rs1[0] ;
    input \imm[9] ;
    input \imm[8] ;
    output \addr_out[27] ;
    output \addr_out[24] ;
    output \addr_out[25] ;
    output \addr_out[26] ;
    output n32829;
    input \imm[5] ;
    input \imm[3] ;
    output n27656;
    input n28909;
    output n27655;
    input n29838;
    input n30172;
    output n27657;
    input n28533;
    output n32548;
    input clk_c_enable_524;
    output n2559;
    output n32834;
    output n32760;
    input n32758;
    output clk_c_enable_187;
    input n28363;
    input n28483;
    output n32538;
    input n32828;
    output address_ready;
    input is_store;
    input mstatus_mie_N_1707;
    output n32710;
    input n30425;
    input n13;
    output n29760;
    output n32668;
    input \mtimecmp[5] ;
    output mtimecmp_1__N_1941;
    input \debug_rd_3__N_405[28] ;
    output n32848;
    input n29844;
    input n32678;
    output n32675;
    input is_alu_imm;
    input is_alu_reg;
    input n28889;
    output n27653;
    input n31351;
    input n29864;
    output clk_c_enable_195;
    output n18;
    input n29317;
    input n32647;
    output n32670;
    output clk_c_enable_28;
    output n32552;
    input n32783;
    output n30928;
    output n30927;
    output n30926;
    output n30925;
    output n30924;
    input n32769;
    input \debug_branch_N_442[31] ;
    input \debug_branch_N_442[30] ;
    input \debug_rd_3__N_405[30] ;
    input \debug_branch_N_442[29] ;
    input \addr_offset[2] ;
    output n28963;
    input \debug_rd_3__N_405[29] ;
    input n157;
    input \debug_branch_N_442[28] ;
    input n28495;
    output n2124;
    input \debug_rd_3__N_405[31] ;
    output n701;
    output \data_out_slice[2] ;
    output debug_early_branch_N_955;
    input no_write_in_progress;
    output n1152;
    input \next_pc_offset[3] ;
    output n28237;
    input \debug_branch_N_450[0] ;
    input n18098;
    input \debug_branch_N_446[28] ;
    input n238;
    input n30070;
    input n76;
    input \mtime_out[0] ;
    input n32717;
    input cy;
    output n32663;
    output n9620;
    input time_pulse_r;
    input n10737;
    output n32680;
    input \next_pc_for_core[7] ;
    input \next_pc_for_core[3] ;
    input \next_pc_for_core[23] ;
    input \next_pc_for_core[19] ;
    output \addr_out[1] ;
    output \addr_out[0] ;
    output n32690;
    output \addr_out[23] ;
    output \addr_out[22] ;
    output \addr_out[21] ;
    output \addr_out[20] ;
    output \addr_out[19] ;
    output \addr_out[18] ;
    output \addr_out[17] ;
    output \addr_out[16] ;
    output \addr_out[15] ;
    output \addr_out[14] ;
    output \addr_out[13] ;
    output \addr_out[12] ;
    output \addr_out[11] ;
    output \addr_out[10] ;
    output \addr_out[9] ;
    output \addr_out[8] ;
    output \addr_out[7] ;
    output \addr_out[6] ;
    output \addr_out[5] ;
    output \addr_out[4] ;
    output \addr_out[3] ;
    input \mem_data_from_read[17] ;
    input \mem_data_from_read[21] ;
    output n32308;
    input \timer_data[1] ;
    input \mul_out[3] ;
    input \mul_out[2] ;
    input [3:0]rd;
    input n32776;
    input \mul_out[1] ;
    input \debug_branch_N_446[31] ;
    input n30175;
    input n29842;
    input \debug_branch_N_446[30] ;
    output \csr_read_3__N_1447[2] ;
    input n29836;
    input \debug_branch_N_446[29] ;
    input n32767;
    input \next_accum[5] ;
    input GND_net;
    input VCC_net;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[4] ;
    input n21667;
    input [3:0]rs1;
    input [3:0]rs2;
    output \reg_access[3][2] ;
    output [23:1]return_addr;
    output \reg_access[4][3] ;
    output n32652;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n10660, n32703;
    wire [5:0]mcause;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(325[15:21])
    
    wire clk_c_enable_347;
    wire [5:0]n611;
    wire [1:0]n979;
    wire [16:0]mie;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(323[16:19])
    
    wire clk_c_enable_335, n31293;
    wire [2:0]time_hi;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(292[15:22])
    wire [2:0]n12;
    
    wire n32354, n32352, n32772, debug_reg_wen, n32350, n32348, 
        n5651, n4862;
    wire [3:0]n5632;
    
    wire n32349, n32347, n31441, mstatus_mpie, clk_c_enable_55, n6299, 
        clk_c_enable_310, n32311, n30171;
    wire [3:0]debug_rd_3__N_1571;
    wire [3:0]n5652;
    
    wire n29868;
    wire [3:0]n5646;
    
    wire n32310, n29671, n25410;
    wire [17:16]mip_reg_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(321[17:24])
    wire [1:0]last_interrupt_req;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(417[15:33])
    wire [1:0]n948;
    wire [1:0]n812;
    
    wire n27929, n32518, n31540, n31545, n32708;
    wire [65:0]dr_3__N_1864;
    
    wire n32402;
    wire [3:0]debug_rd_3__N_1392;
    wire [3:0]debug_rd_3__N_1396;
    
    wire n32882, n32881, n32894, n32893, n33040, n46;
    wire [3:0]n653;
    wire [3:0]n658;
    
    wire n32839, n29245, n32645, clk_c_enable_520, cmp, cmp_out;
    wire [3:0]instrret_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(301[16:30])
    
    wire n31616;
    wire [31:0]tmp_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(88[16:24])
    
    wire clk_c_enable_540, cy_c, instr_retired, n32683;
    wire [23:0]mepc;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(68[16:20])
    
    wire n31617, cy_adj_3149, n32748, n32688, n29882;
    wire [6:0]cycle_count_wide;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(279[16:32])
    
    wire cy_adj_3150, n32701;
    wire [4:0]increment_result_3__N_1911;
    
    wire n32805, n15, n32807, n30243, n32827, n32724, n29867, 
        n32736;
    wire [3:0]n196;
    wire [3:0]n191;
    wire [3:0]debug_rd_3__N_1559;
    
    wire n18087;
    wire [3:0]time_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(299[16:26])
    
    wire clk_c_enable_348, n29009, n11035, cy_out, clk_c_enable_115, 
        mstatus_mte_N_1703;
    wire [5:0]shift_amt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[16:25])
    
    wire clk_c_enable_436, n28179, n32804, n29411;
    wire [3:0]shift_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(132[16:25])
    
    wire n31407, n29851, n29852, n29853;
    wire [2:0]n5080;
    
    wire n27861;
    wire [3:0]alu_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(110[16:23])
    
    wire n32747, n31542, n31541, n32750;
    wire [3:0]csr_read_3__N_1439;
    wire [3:0]csr_read_3__N_1455;
    
    wire n17982, n34004, n34002, n34003, n27933, n27987;
    wire [2:0]n498;
    
    wire n32790, n34005, n34278, n34006, n30231, n32792, n40, 
        n29647, n32793, n101, n32794, n29011, n25980, clk_c_enable_316, 
        n25984;
    wire [59:0]debug_branch_N_840;
    
    wire n927, n928, n31408, n25986, n894, n895, clk_c_enable_332, 
        n25978;
    wire [3:0]tmp_data_in_3__N_1514;
    
    wire n861, n34277, n862, n25982, n794, n27994, n26364, instr_complete_N_1656, 
        instr_complete_N_1654, n32404, n31406, n31419, n30051, debug_rd_3__N_1401, 
        instr_complete_N_1650, n34276, n6086, n32738;
    wire [3:0]alu_b_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[16:24])
    
    wire n32624, n34007, n30073, n32625, n32626, n32646, n32749;
    wire [3:0]data_rs1_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(83[16:24])
    wire [1:0]n809;
    wire [3:0]tmp_data_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(242[15:26])
    
    wire n26850, n11722;
    wire [3:0]csr_read_3__N_1451;
    
    wire n31618, n29875, n32816;
    wire [4:0]shift_amt_adj_3153;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(124[15:24])
    
    wire clk_c_enable_437, n27962;
    wire [3:0]n5605;
    
    wire n32676, n14, n31292, n10687, n31428, n31425, n29445, 
        n29443, n31426, n31427, n32831, n29669, n28903;
    wire [3:0]n234;
    
    wire n31410, n28897, n31409, n9909, n29683, mstatus_mie;
    wire [3:0]csr_read_3__N_1637;
    
    wire n29881, load_top_bit_next_N_1731, n18385, clk_c_enable_522, 
        n31420, n32731, n34292, n10675, n26807, n31423, instr_complete_N_1648, 
        n17772, n32705, n11720;
    wire [3:0]csr_read_3__N_1443;
    
    wire n29227;
    wire [3:0]mul_out_3__N_1510;
    
    wire n29425, n652;
    wire [3:0]alu_a_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[16:24])
    
    wire alu_b_in_3__N_1504, n32883, n32699, instr_complete_N_1649;
    wire [3:0]tmp_data_in_3__N_1582;
    
    wire n30193, n27960;
    wire [3:0]debug_rd_3__N_1567;
    
    wire n27723;
    wire [4:0]increment_result_3__N_1925;
    
    wire n29121, n32665, interrupt_pending_N_1671, n28225, n10727, 
        n32592, n32353, n33042, n33039, n7739, n17891, n57;
    wire [3:0]n4826;
    
    wire n5721, n32401, n31758, n31760;
    wire [3:0]n4901;
    
    wire n33043, n33041, n32403;
    wire [1:0]n822;
    
    LUT4 i1_2_lut_rep_688 (.A(\imm[6] ), .B(n10660), .Z(n32703)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_2_lut_rep_688.init = 16'heeee;
    FD1P3IX mcause__i0 (.D(n611[0]), .SP(clk_c_enable_347), .CD(n32840), 
            .CK(clk_c), .Q(mcause[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i0.GSR = "DISABLED";
    FD1P3IX mip_reg__i16 (.D(n979[0]), .SP(clk_c_enable_342), .CD(n32650), 
            .CK(clk_c), .Q(mip_reg[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mip_reg__i16.GSR = "DISABLED";
    FD1P3IX mie__i0 (.D(n31293), .SP(clk_c_enable_335), .CD(n32650), .CK(clk_c), 
            .Q(mie[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i0.GSR = "DISABLED";
    FD1S3IX time_hi__i0 (.D(n12[0]), .CK(clk_c), .CD(n32840), .Q(time_hi[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i0.GSR = "DISABLED";
    PFUMX i29202 (.BLUT(n32354), .ALUT(n32352), .C0(n32772), .Z(debug_reg_wen));
    L6MUX21 i29199 (.D0(n32350), .D1(n32348), .SD(n5651), .Z(n32351));
    LUT4 i1_3_lut (.A(counter_hi[4]), .B(counter_hi[2]), .C(counter_hi[3]), 
         .Z(n4862)) /* synthesis lut_function=(A+!((C)+!B)) */ ;
    defparam i1_3_lut.init = 16'haeae;
    PFUMX i29197 (.BLUT(n5632[0]), .ALUT(n32349), .C0(\imm[10] ), .Z(n32350));
    PFUMX i29195 (.BLUT(n32347), .ALUT(n31441), .C0(\imm[0] ), .Z(n32348));
    FD1P3AX mstatus_mpie_525 (.D(n6299), .SP(clk_c_enable_55), .CK(clk_c), 
            .Q(mstatus_mpie)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam mstatus_mpie_525.GSR = "DISABLED";
    LUT4 i28486_2_lut_3_lut_4_lut (.A(\imm[6] ), .B(n10660), .C(n32759), 
         .D(\imm[2] ), .Z(clk_c_enable_310)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i28486_2_lut_3_lut_4_lut.init = 16'h0100;
    PFUMX i29173 (.BLUT(n32311), .ALUT(\debug_branch_N_450[1] ), .C0(n30171), 
          .Z(debug_rd_3__N_1571[1]));
    L6MUX21 mux_3507_i3 (.D0(n5652[2]), .D1(n29868), .SD(n5651), .Z(n5660));
    PFUMX mux_3507_i2 (.BLUT(n5652[1]), .ALUT(n5646[1]), .C0(n5651), .Z(n5661));
    PFUMX i29171 (.BLUT(n30329), .ALUT(n32309), .C0(counter_hi[4]), .Z(n32310));
    LUT4 i27027_3_lut_4_lut (.A(\imm[6] ), .B(n10660), .C(\imm[2] ), .D(n32759), 
         .Z(n29671)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i27027_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut (.A(instr_complete_N_1647), .B(clk_c_enable_285), 
         .C(cycle[1]), .D(cycle[0]), .Z(n25410)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_4_lut.init = 16'h0770;
    LUT4 i1_2_lut_rep_687_3_lut_4_lut_3_lut_4_lut (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .C(is_system), .D(debug_instr_valid), .Z(n32702)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_2_lut_rep_687_3_lut_4_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 is_csr_I_0_573_2_lut_rep_718_3_lut_4_lut_3_lut_4_lut (.A(\alu_op[0] ), 
         .B(\alu_op[1] ), .C(is_system), .D(debug_instr_valid), .Z(n32733)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam is_csr_I_0_573_2_lut_rep_718_3_lut_4_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_689_3_lut_4_lut_3_lut_4_lut (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .C(is_system), .D(debug_instr_valid), .Z(n32704)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_2_lut_rep_689_3_lut_4_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut (.A(n32746), .B(mip_reg_c[17]), .C(\ui_in_sync[1] ), 
         .D(last_interrupt_req[1]), .Z(n948[1])) /* synthesis lut_function=(A (B+!((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(482[33:47])
    defparam i1_4_lut.init = 16'h88a8;
    LUT4 i1_4_lut_adj_300 (.A(n10660), .B(n812[1]), .C(n24384), .D(\imm[2] ), 
         .Z(n27929)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_300.init = 16'h4000;
    PFUMX i28728 (.BLUT(n32518), .ALUT(n31540), .C0(\imm[6] ), .Z(n31545));
    LUT4 interrupt_core_I_32_2_lut_rep_530_4_lut (.A(stall_core), .B(instr_complete_N_1647), 
         .C(n32708), .D(n32774), .Z(n32545)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam interrupt_core_I_32_2_lut_rep_530_4_lut.init = 16'h80ff;
    LUT4 i1_2_lut_4_lut (.A(stall_core), .B(instr_complete_N_1647), .C(n32708), 
         .D(is_load), .Z(n829)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_4_lut.init = 16'h80ff;
    LUT4 i1_2_lut_4_lut_adj_301 (.A(stall_core), .B(instr_complete_N_1647), 
         .C(n32708), .D(n26962), .Z(clk_c_enable_533)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_4_lut_adj_301.init = 16'hff80;
    LUT4 dr_3__N_1864_31__bdd_3_lut_29288 (.A(dr_3__N_1864[31]), .B(dr_3__N_1864[34]), 
         .C(\alu_op_in[2] ), .Z(n32402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam dr_3__N_1864_31__bdd_3_lut_29288.init = 16'hcaca;
    LUT4 i1_4_lut_adj_302 (.A(n32746), .B(mip_reg[16]), .C(\ui_in_sync[0] ), 
         .D(last_interrupt_req[0]), .Z(n948[0])) /* synthesis lut_function=(A (B+!((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(482[33:47])
    defparam i1_4_lut_adj_302.init = 16'h88a8;
    LUT4 n14411_bdd_2_lut_3_lut_4_lut_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .D(mip_reg_c[17]), .Z(n31540)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam n14411_bdd_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 debug_rd_3__I_0_i1_3_lut (.A(debug_rd_3__N_1392[0]), .B(debug_rd_3__N_1396[0]), 
         .C(n32772), .Z(debug_rd[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(176[18] 194[12])
    defparam debug_rd_3__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 n30235_bdd_4_lut_28805_then_4_lut (.A(mie[12]), .B(mie[4]), .C(counter_hi[4]), 
         .D(counter_hi[3]), .Z(n32882)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(((D)+!C)+!B)) */ ;
    defparam n30235_bdd_4_lut_28805_then_4_lut.init = 16'ha0c0;
    LUT4 n30235_bdd_4_lut_28805_else_4_lut (.A(mie[0]), .B(counter_hi[4]), 
         .C(counter_hi[3]), .D(mie[8]), .Z(n32881)) /* synthesis lut_function=(A (B ((D)+!C))+!A (B (C (D)))) */ ;
    defparam n30235_bdd_4_lut_28805_else_4_lut.init = 16'hc808;
    LUT4 n31548_bdd_4_lut_then_4_lut (.A(\mie[10] ), .B(\mie[14] ), .C(counter_hi[2]), 
         .D(counter_hi[4]), .Z(n32894)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n31548_bdd_4_lut_then_4_lut.init = 16'hca00;
    LUT4 n31548_bdd_4_lut_else_4_lut (.A(\mie[2] ), .B(\mie[6] ), .C(counter_hi[2]), 
         .D(counter_hi[4]), .Z(n32893)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n31548_bdd_4_lut_else_4_lut.init = 16'hca00;
    LUT4 mux_351_i2_3_lut_4_lut (.A(clk_c_enable_285), .B(n27294), .C(n5017[1]), 
         .D(n1766), .Z(\instr_write_offset_3__N_934[1] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_351_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_351_i1_3_lut_4_lut (.A(clk_c_enable_285), .B(n27294), .C(n5017[0]), 
         .D(n1767), .Z(\instr_write_offset_3__N_934[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_351_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_352_i1_3_lut_4_lut (.A(clk_c_enable_285), .B(n27294), .C(n5017[0]), 
         .D(n1768[0]), .Z(pc_2__N_932[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_352_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 next_pc_for_core_23__bdd_3_lut (.A(\next_pc_for_core[15] ), .B(\next_pc_for_core[11] ), 
         .C(counter_hi[2]), .Z(n33040)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam next_pc_for_core_23__bdd_3_lut.init = 16'hacac;
    LUT4 i1_3_lut_4_lut_adj_303 (.A(n32846), .B(n32847), .C(\imm[7] ), 
         .D(n46), .Z(n9058)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(75[19:52])
    defparam i1_3_lut_4_lut_adj_303.init = 16'h0800;
    PFUMX mux_252_i1 (.BLUT(n653[0]), .ALUT(n29689), .C0(n32691), .Z(n658[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 interrupt_core_I_31_2_lut_rep_528_3_lut_4_lut (.A(clk_c_enable_285), 
         .B(n27294), .C(n32549), .D(n32774), .Z(n32543)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (C+!(D))) */ ;
    defparam interrupt_core_I_31_2_lut_rep_528_3_lut_4_lut.init = 16'hf8ff;
    LUT4 mux_352_i2_3_lut_4_lut (.A(clk_c_enable_285), .B(n27294), .C(n5017[1]), 
         .D(n1768[1]), .Z(pc_2__N_932[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_352_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_535_3_lut_4_lut (.A(clk_c_enable_285), .B(n27294), 
         .C(instr_fetch_running), .D(was_early_branch), .Z(n32550)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (C))) */ ;
    defparam i1_2_lut_rep_535_3_lut_4_lut.init = 16'h0f07;
    LUT4 data_ready_sync_I_0_3_lut_4_lut (.A(n32839), .B(counter_hi[2]), 
         .C(n32564), .D(data_ready_sync), .Z(data_ready_core)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam data_ready_sync_I_0_3_lut_4_lut.init = 16'hfe10;
    LUT4 i28324_4_lut (.A(n32650), .B(n29245), .C(n32645), .D(n131), 
         .Z(clk_c_enable_520)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i28324_4_lut.init = 16'hfbfa;
    LUT4 i1_2_lut_rep_682_3_lut_4_lut (.A(n32839), .B(counter_hi[2]), .C(n32768), 
         .D(n32849), .Z(n32697)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_2_lut_rep_682_3_lut_4_lut.init = 16'h0010;
    FD1S3AX cmp_511 (.D(cmp_out), .CK(clk_c), .Q(cmp)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(117[12] 120[8])
    defparam cmp_511.GSR = "DISABLED";
    LUT4 imm_10__bdd_3_lut_28774_3_lut_4_lut (.A(n32839), .B(counter_hi[2]), 
         .C(instrret_count[1]), .D(\imm[0] ), .Z(n31616)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam imm_10__bdd_3_lut_28774_3_lut_4_lut.init = 16'h11f0;
    FD1P3AX tmp_data_i0_i0 (.D(tmp_data[4]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i0.GSR = "DISABLED";
    LUT4 cy_I_0_3_lut_rep_668_3_lut_4_lut (.A(n32839), .B(counter_hi[2]), 
         .C(cy_c), .D(instr_retired), .Z(n32683)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam cy_I_0_3_lut_rep_668_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX mepc_i0_i0 (.D(mepc[4]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i0.GSR = "DISABLED";
    LUT4 imm_10__bdd_3_lut_3_lut_4_lut (.A(n32839), .B(counter_hi[2]), .C(\imm[1] ), 
         .D(mcause[1]), .Z(n31617)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam imm_10__bdd_3_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 cy_I_0_3_lut_rep_673_3_lut_4_lut (.A(n32839), .B(counter_hi[2]), 
         .C(cy_adj_3149), .D(n32748), .Z(n32688)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam cy_I_0_3_lut_rep_673_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i27173_3_lut_3_lut_4_lut (.A(n32839), .B(counter_hi[2]), .C(instrret_count[0]), 
         .D(\imm[0] ), .Z(n29882)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i27173_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i4727_2_lut_rep_686_3_lut_4_lut (.A(n32839), .B(counter_hi[2]), 
         .C(cycle_count_wide[0]), .D(cy_adj_3150), .Z(n32701)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i4727_2_lut_rep_686_3_lut_4_lut.init = 16'hf010;
    LUT4 i4725_2_lut_3_lut_4_lut (.A(n32839), .B(counter_hi[2]), .C(cycle_count_wide[0]), 
         .D(cy_adj_3150), .Z(increment_result_3__N_1911[0])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i4725_2_lut_3_lut_4_lut.init = 16'h0fe1;
    LUT4 i28526_3_lut_4_lut (.A(n32805), .B(n32838), .C(n15), .D(n32807), 
         .Z(n30243)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i28526_3_lut_4_lut.init = 16'hffdf;
    LUT4 i1_2_lut_rep_709_4_lut (.A(\alu_op_in[2] ), .B(n32847), .C(n32846), 
         .D(n32827), .Z(n32724)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_709_4_lut.init = 16'h1000;
    PFUMX i27159 (.BLUT(n29866), .ALUT(n29867), .C0(\imm[0] ), .Z(n29868));
    LUT4 i1_2_lut_rep_721_4_lut (.A(\alu_op_in[2] ), .B(n32847), .C(n32846), 
         .D(n32849), .Z(n32736)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_721_4_lut.init = 16'h0010;
    FD1P3AX last_interrupt_req_i0_i0 (.D(\ui_in_sync[0] ), .SP(clk_c_enable_433), 
            .CK(clk_c), .Q(last_interrupt_req[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam last_interrupt_req_i0_i0.GSR = "DISABLED";
    LUT4 i28051_4_lut_4_lut (.A(n32807), .B(n15), .C(n196[0]), .D(n191[0]), 
         .Z(debug_rd_3__N_1559[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;
    defparam i28051_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i28094_3_lut_4_lut_4_lut (.A(n32807), .B(debug_rd_3__N_1559[3]), 
         .C(n32805), .D(tmp_data[3]), .Z(debug_rd_3__N_1396[3])) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam i28094_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 i15438_2_lut_3_lut_4_lut (.A(counter_hi[4]), .B(n32854), .C(interrupt_core), 
         .D(stall_core), .Z(n18087)) /* synthesis lut_function=(!(A (B (C+(D))))) */ ;
    defparam i15438_2_lut_3_lut_4_lut.init = 16'h777f;
    LUT4 cycle_count_wide_6__I_0_3_lut_4_lut (.A(counter_hi[4]), .B(n32854), 
         .C(time_hi[2]), .D(cycle_count_wide[6]), .Z(time_count[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam cycle_count_wide_6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i28316_2_lut_3_lut_4_lut (.A(counter_hi[4]), .B(n32854), .C(rst_reg_n), 
         .D(n17920), .Z(clk_c_enable_348)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i28316_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 cycle_count_wide_5__I_0_3_lut_4_lut (.A(counter_hi[4]), .B(n32854), 
         .C(time_hi[1]), .D(cycle_count_wide[5]), .Z(time_count[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam cycle_count_wide_5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut (.A(counter_hi[4]), .B(n32854), .C(n28685), 
         .D(n27294), .Z(n28687)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i8335_4_lut (.A(n34285), .B(n29009), .C(is_lui), .D(is_jal), 
         .Z(n11035)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(218[17:110])
    defparam i8335_4_lut.init = 16'haaa8;
    FD1S3AX cy_510 (.D(cy_out), .CK(clk_c), .Q(cy_adj_3149)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(117[12] 120[8])
    defparam cy_510.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_304 (.A(is_branch), .B(is_jalr), .C(is_auipc), .D(is_system), 
         .Z(n29009)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(218[17:110])
    defparam i1_4_lut_adj_304.init = 16'hfffe;
    LUT4 debug_branch_N_441_I_0_2_lut_rep_536_3_lut_4_lut (.A(n34281), .B(n32854), 
         .C(was_early_branch), .D(n27294), .Z(n32551)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam debug_branch_N_441_I_0_2_lut_rep_536_3_lut_4_lut.init = 16'hf7ff;
    FD1P3BX mstatus_mte_523 (.D(mstatus_mte_N_1703), .SP(clk_c_enable_115), 
            .CK(clk_c), .PD(n32840), .Q(mstatus_mte)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(384[18] 390[12])
    defparam mstatus_mte_523.GSR = "DISABLED";
    FD1P3AX shift_amt__i1 (.D(n92[0]), .SP(clk_c_enable_436), .CK(clk_c), 
            .Q(shift_amt[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i1.GSR = "DISABLED";
    LUT4 cycle_count_wide_4__I_0_3_lut_4_lut (.A(counter_hi[4]), .B(n32854), 
         .C(time_hi[0]), .D(cycle_count_wide[4]), .Z(time_count[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam cycle_count_wide_4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i24427_2_lut_3_lut_4_lut (.A(n34281), .B(n32854), .C(n34287), 
         .D(n27294), .Z(n27003)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i24427_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i1_4_lut_adj_305 (.A(n28179), .B(cmp_out), .C(n32821), .D(mem_op[0]), 
         .Z(n27294)) /* synthesis lut_function=(A+!(B ((D)+!C)+!B !(C (D)))) */ ;
    defparam i1_4_lut_adj_305.init = 16'hbaea;
    LUT4 i1_4_lut_adj_306 (.A(n32736), .B(n32724), .C(n32741), .D(interrupt_core), 
         .Z(n28179)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_306.init = 16'hfffe;
    LUT4 i1_4_lut_adj_307 (.A(cycle[0]), .B(n32804), .C(n32839), .D(n29411), 
         .Z(n15)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_4_lut_adj_307.init = 16'hfffd;
    LUT4 i1_3_lut_adj_308 (.A(\alu_op[3] ), .B(counter_hi[2]), .C(cycle[1]), 
         .Z(n29411)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_3_lut_adj_308.init = 16'hfefe;
    LUT4 n194_bdd_4_lut_29032 (.A(n191[1]), .B(shift_out[1]), .C(n32805), 
         .D(n32838), .Z(n31407)) /* synthesis lut_function=(A (B+((D)+!C))+!A !(((D)+!C)+!B)) */ ;
    defparam n194_bdd_4_lut_29032.init = 16'haaca;
    L6MUX21 i27144 (.D0(n29851), .D1(n29852), .SD(\imm[10] ), .Z(n29853));
    PFUMX mux_233_i1 (.BLUT(n5080[0]), .ALUT(n27861), .C0(interrupt_core), 
          .Z(n611[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 mux_73_i1_4_lut (.A(cmp), .B(tmp_data[0]), .C(n32807), .D(n32805), 
         .Z(n196[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(170[18] 174[35])
    defparam mux_73_i1_4_lut.init = 16'hca0a;
    LUT4 mux_72_i1_4_lut (.A(accum[0]), .B(alu_out[0]), .C(n32747), .D(d_3__N_1868[0]), 
         .Z(n191[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(174[17:35])
    defparam mux_72_i1_4_lut.init = 16'hc5ca;
    LUT4 i28567_3_lut (.A(data_out_3__N_1385), .B(is_timer_addr), .C(n30160), 
         .Z(n30171)) /* synthesis lut_function=(A+!(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam i28567_3_lut.init = 16'habab;
    LUT4 n31542_bdd_4_lut (.A(n31542), .B(n31541), .C(n32750), .D(n4862), 
         .Z(n32518)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n31542_bdd_4_lut.init = 16'hca00;
    LUT4 is_jal_I_0_2_lut_rep_769 (.A(is_jal), .B(is_jalr), .Z(n32784)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam is_jal_I_0_2_lut_rep_769.init = 16'heeee;
    LUT4 i1_2_lut_rep_662_3_lut (.A(\imm[6] ), .B(n10660), .C(\imm[2] ), 
         .Z(n32677)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_2_lut_rep_662_3_lut.init = 16'hefef;
    LUT4 i5893_2_lut_rep_726_3_lut (.A(is_jal), .B(is_jalr), .C(debug_instr_valid), 
         .Z(n32741)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam i5893_2_lut_rep_726_3_lut.init = 16'he0e0;
    PFUMX i27142 (.BLUT(csr_read_3__N_1439[3]), .ALUT(csr_read_3__N_1455[3]), 
          .C0(\imm[1] ), .Z(n29851));
    LUT4 debug_rd_3__I_0_i2_3_lut_4_lut (.A(n32772), .B(debug_rd_3__N_1575), 
         .C(debug_rd_3__N_1392[1]), .D(debug_rd_3__N_1571[1]), .Z(debug_rd[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(176[18] 194[12])
    defparam debug_rd_3__I_0_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mie_3__bdd_4_lut (.A(mie[3]), .B(n17982), .C(counter_hi[2]), 
         .D(counter_hi[4]), .Z(n34004)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mie_3__bdd_4_lut.init = 16'hcac0;
    LUT4 mepc_3__bdd_4_lut (.A(mepc[3]), .B(counter_hi[3]), .C(\imm[6] ), 
         .D(counter_hi[4]), .Z(n34002)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;
    defparam mepc_3__bdd_4_lut.init = 16'h20a0;
    LUT4 mie_3__bdd_4_lut_29864 (.A(mie[15]), .B(counter_hi[2]), .C(counter_hi[4]), 
         .D(mie[11]), .Z(n34003)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(B+!(C (D)))) */ ;
    defparam mie_3__bdd_4_lut_29864.init = 16'hb080;
    PFUMX i66 (.BLUT(n27933), .ALUT(n27987), .C0(\imm[11] ), .Z(n46));
    FD1P3IX time_hi__i2 (.D(n498[2]), .SP(clk_c_enable_276), .CD(n32840), 
            .CK(clk_c), .Q(time_hi[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i2.GSR = "DISABLED";
    FD1P3IX time_hi__i1 (.D(n498[1]), .SP(clk_c_enable_276), .CD(n32840), 
            .CK(clk_c), .Q(time_hi[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i1.GSR = "DISABLED";
    LUT4 i28538_2_lut_rep_775 (.A(\imm[1] ), .B(\imm[0] ), .Z(n32790)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i28538_2_lut_rep_775.init = 16'hbbbb;
    LUT4 n34005_bdd_3_lut (.A(n34005), .B(n34278), .C(\imm[6] ), .Z(n34006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n34005_bdd_3_lut.init = 16'hcaca;
    LUT4 i28540_2_lut_3_lut (.A(\imm[1] ), .B(\imm[0] ), .C(\imm[10] ), 
         .Z(n30231)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i28540_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i27016_2_lut_rep_776 (.A(fsm_state[1]), .B(fsm_state[3]), .Z(n32791)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i27016_2_lut_rep_776.init = 16'heeee;
    LUT4 i1_2_lut_rep_748_3_lut (.A(fsm_state[1]), .B(fsm_state[3]), .C(fsm_state[2]), 
         .Z(n32763)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_748_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_715_3_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[3]), 
         .C(fsm_state[0]), .D(fsm_state[2]), .Z(n32730)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_715_3_lut_4_lut.init = 16'hfffe;
    LUT4 and_454_i1_2_lut_rep_777 (.A(mip_reg[16]), .B(mie[0]), .Z(n32792)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[48:59])
    defparam and_454_i1_2_lut_rep_777.init = 16'h8888;
    LUT4 i1_4_lut_4_lut (.A(\imm[2] ), .B(n40), .C(\imm[10] ), .D(n29647), 
         .Z(n27987)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i1_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_778 (.A(mie[16]), .B(timer_interrupt), .Z(n32793)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_778.init = 16'h8888;
    LUT4 i15331_2_lut_3_lut (.A(mie[16]), .B(timer_interrupt), .C(interrupt_core), 
         .Z(n611[2])) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15331_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut (.A(mie[16]), .B(timer_interrupt), .C(interrupt_core), 
         .Z(n101)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_779 (.A(mip_reg_c[17]), .B(mie[1]), .Z(n32794)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam i1_2_lut_rep_779.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_309 (.A(mip_reg_c[17]), .B(mie[1]), .C(timer_interrupt), 
         .D(mie[16]), .Z(n29011)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam i1_2_lut_3_lut_4_lut_adj_309.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_310 (.A(\imm[6] ), .B(n10660), .C(\imm[2] ), 
         .D(n32765), .Z(n29245)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_3_lut_4_lut_adj_310.init = 16'hfffe;
    PFUMX mux_3505_i3 (.BLUT(time_count[2]), .ALUT(n5642), .C0(n30231), 
          .Z(n5652[2]));
    FD1P3IX mie__i16 (.D(n25980), .SP(clk_c_enable_310), .CD(n32650), 
            .CK(clk_c), .Q(mie[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i16.GSR = "DISABLED";
    FD1P3IX mie__i15 (.D(n25984), .SP(clk_c_enable_316), .CD(n32650), 
            .CK(clk_c), .Q(mie[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i15.GSR = "DISABLED";
    FD1P3IX mie__i14 (.D(n926), .SP(clk_c_enable_316), .CD(n32650), .CK(clk_c), 
            .Q(\mie[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i14.GSR = "DISABLED";
    LUT4 i28071_3_lut (.A(n33057), .B(\timer_data[0] ), .C(is_timer_addr), 
         .Z(debug_branch_N_840[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam i28071_3_lut.init = 16'hcaca;
    FD1P3IX mie__i13 (.D(n927), .SP(clk_c_enable_316), .CD(n32650), .CK(clk_c), 
            .Q(mie[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i13.GSR = "DISABLED";
    FD1P3IX mie__i12 (.D(n928), .SP(clk_c_enable_316), .CD(n32650), .CK(clk_c), 
            .Q(mie[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i12.GSR = "DISABLED";
    LUT4 gnd_bdd_2_lut_28673 (.A(n31407), .B(n15), .Z(n31408)) /* synthesis lut_function=(A (B)) */ ;
    defparam gnd_bdd_2_lut_28673.init = 16'h8888;
    FD1P3IX mie__i11 (.D(n25986), .SP(clk_c_enable_321), .CD(n32650), 
            .CK(clk_c), .Q(mie[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i11.GSR = "DISABLED";
    FD1P3IX mie__i10 (.D(n893), .SP(clk_c_enable_321), .CD(n32650), .CK(clk_c), 
            .Q(\mie[10] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i10.GSR = "DISABLED";
    FD1P3IX mie__i9 (.D(n894), .SP(clk_c_enable_321), .CD(n32650), .CK(clk_c), 
            .Q(mie[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i9.GSR = "DISABLED";
    FD1P3IX mie__i8 (.D(n895), .SP(clk_c_enable_321), .CD(n32650), .CK(clk_c), 
            .Q(mie[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i8.GSR = "DISABLED";
    FD1P3AX load_done_515 (.D(n8228), .SP(clk_c_enable_363), .CK(clk_c), 
            .Q(load_done)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(232[12] 235[8])
    defparam load_done_515.GSR = "DISABLED";
    FD1P3IX mie__i7 (.D(n25978), .SP(clk_c_enable_332), .CD(n32650), .CK(clk_c), 
            .Q(mie[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i7.GSR = "DISABLED";
    LUT4 i28078_3_lut (.A(n32317), .B(\timer_data[2] ), .C(is_timer_addr), 
         .Z(debug_branch_N_840[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam i28078_3_lut.init = 16'hcaca;
    LUT4 tmp_data_in_3__I_124_i3_4_lut (.A(data_rs1[2]), .B(mstatus_mte), 
         .C(n32691), .D(n32697), .Z(tmp_data_in_3__N_1514[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_124_i3_4_lut.init = 16'hca0a;
    FD1P3IX mie__i6 (.D(n860), .SP(clk_c_enable_332), .CD(n32650), .CK(clk_c), 
            .Q(\mie[6] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i6.GSR = "DISABLED";
    FD1P3IX mie__i5 (.D(n861), .SP(clk_c_enable_332), .CD(n32650), .CK(clk_c), 
            .Q(mie[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i5.GSR = "DISABLED";
    LUT4 n17983_bdd_4_lut_29419_then_4_lut (.A(timer_interrupt), .B(counter_hi[4]), 
         .C(counter_hi[3]), .D(counter_hi[2]), .Z(n34277)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam n17983_bdd_4_lut_29419_then_4_lut.init = 16'h0200;
    FD1P3IX mie__i4 (.D(n862), .SP(clk_c_enable_332), .CD(n32650), .CK(clk_c), 
            .Q(mie[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i4.GSR = "DISABLED";
    FD1P3IX mie__i3 (.D(n25982), .SP(clk_c_enable_335), .CD(n32650), .CK(clk_c), 
            .Q(mie[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i3.GSR = "DISABLED";
    FD1P3IX mie__i2 (.D(n793), .SP(clk_c_enable_335), .CD(n32650), .CK(clk_c), 
            .Q(\mie[2] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i2.GSR = "DISABLED";
    FD1P3IX mie__i1 (.D(n794), .SP(clk_c_enable_335), .CD(n32650), .CK(clk_c), 
            .Q(mie[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i1.GSR = "DISABLED";
    FD1P3IX mip_reg__i17 (.D(n979[1]), .SP(clk_c_enable_342), .CD(n32650), 
            .CK(clk_c), .Q(mip_reg_c[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mip_reg__i17.GSR = "DISABLED";
    FD1P3IX mcause__i5 (.D(interrupt_core), .SP(clk_c_enable_347), .CD(n32840), 
            .CK(clk_c), .Q(mcause[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i5.GSR = "DISABLED";
    FD1P3IX mcause__i4 (.D(n101), .SP(clk_c_enable_347), .CD(n32840), 
            .CK(clk_c), .Q(mcause[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i4.GSR = "DISABLED";
    LUT4 i6651_4_lut_4_lut (.A(n32546), .B(n28417), .C(n32580), .D(n32642), 
         .Z(n3274)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i6651_4_lut_4_lut.init = 16'hfb40;
    FD1P3IX mcause__i3 (.D(n27994), .SP(clk_c_enable_347), .CD(n32840), 
            .CK(clk_c), .Q(mcause[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i3.GSR = "DISABLED";
    FD1P3IX mcause__i2 (.D(n611[2]), .SP(clk_c_enable_347), .CD(n32840), 
            .CK(clk_c), .Q(mcause[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i2.GSR = "DISABLED";
    FD1P3IX mcause__i1 (.D(n26364), .SP(clk_c_enable_347), .CD(n32840), 
            .CK(clk_c), .Q(mcause[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i1.GSR = "DISABLED";
    FD1P3IX cycle__i1 (.D(n25410), .SP(clk_c_enable_348), .CD(n32840), 
            .CK(clk_c), .Q(cycle[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam cycle__i1.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_adj_311 (.A(n32546), .B(n28429), .C(n32543), .D(n4), 
         .Z(n27546)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_311.init = 16'h4000;
    LUT4 i1_4_lut_4_lut_adj_312 (.A(n32546), .B(n28465), .C(n32543), .D(n4), 
         .Z(n27541)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_312.init = 16'h4000;
    LUT4 i1_3_lut_adj_313 (.A(tmp_data[30]), .B(tmp_data[31]), .C(cycle[0]), 
         .Z(instr_complete_N_1656)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_adj_313.init = 16'hf7f7;
    LUT4 cycle_0__I_0_548_3_lut (.A(cycle[0]), .B(cmp_out), .C(\alu_op[0] ), 
         .Z(instr_complete_N_1654)) /* synthesis lut_function=(A+!(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(224[34:67])
    defparam cycle_0__I_0_548_3_lut.init = 16'hbebe;
    LUT4 i15321_2_lut (.A(n32404), .B(n15), .Z(debug_rd_3__N_1559[3])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[18] 174[35])
    defparam i15321_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_789 (.A(\alu_op_in[2] ), .B(\alu_op[1] ), .Z(n32804)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam i1_2_lut_rep_789.init = 16'hbbbb;
    LUT4 mux_87_i4_3_lut (.A(\debug_branch_N_450[3] ), .B(load_top_bit), 
         .C(data_out_3__N_1385), .Z(debug_rd_3__N_1571[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam mux_87_i4_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_732_3_lut (.A(\alu_op_in[2] ), .B(\alu_op[1] ), .C(\alu_op[3] ), 
         .Z(n32747)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam i1_2_lut_rep_732_3_lut.init = 16'hbfbf;
    LUT4 i28384_2_lut_rep_790 (.A(cycle[0]), .B(cycle[1]), .Z(n32805)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam i28384_2_lut_rep_790.init = 16'h2222;
    LUT4 n194_bdd_2_lut_29031_3_lut (.A(cycle[0]), .B(cycle[1]), .C(tmp_data[1]), 
         .Z(n31406)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam n194_bdd_2_lut_29031_3_lut.init = 16'h2020;
    LUT4 n193_bdd_2_lut_3_lut (.A(cycle[0]), .B(cycle[1]), .C(tmp_data[2]), 
         .Z(n31419)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam n193_bdd_2_lut_3_lut.init = 16'h2020;
    LUT4 i5881_3_lut_rep_791 (.A(n34285), .B(is_auipc), .C(is_jal), .Z(n32806)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(108[27:47])
    defparam i5881_3_lut_rep_791.init = 16'ha8a8;
    LUT4 i27342_2_lut_4_lut (.A(n34285), .B(is_auipc), .C(is_jal), .D(n32808), 
         .Z(n30051)) /* synthesis lut_function=(A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(108[27:47])
    defparam i27342_2_lut_4_lut.init = 16'ha800;
    PFUMX instr_complete_I_133 (.BLUT(instr_complete_N_1651), .ALUT(instr_complete_N_1652), 
          .C0(debug_rd_3__N_1401), .Z(instr_complete_N_1650)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_rep_792 (.A(\alu_op[1] ), .B(\alu_op_in[2] ), .C(\alu_op[3] ), 
         .Z(n32807)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_792.init = 16'h8080;
    LUT4 n17983_bdd_4_lut_29419_else_4_lut (.A(timer_interrupt), .B(counter_hi[4]), 
         .C(counter_hi[3]), .D(counter_hi[2]), .Z(n34276)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam n17983_bdd_4_lut_29419_else_4_lut.init = 16'h020c;
    FD1P3IX is_double_fault_r_520 (.D(n32736), .SP(clk_c_enable_363), .CD(n6086), 
            .CK(clk_c), .Q(is_double_fault_r)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(361[12] 364[8])
    defparam is_double_fault_r_520.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_adj_314 (.A(n32546), .B(n28441), .C(n32543), .D(n4), 
         .Z(n27545)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_314.init = 16'h4000;
    LUT4 i15313_2_lut_rep_723_3_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .Z(n32738)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i15313_2_lut_rep_723_3_lut.init = 16'h2a2a;
    LUT4 i13_3_lut_4_lut (.A(\alu_op[0] ), .B(n32732), .C(data_rs1[2]), 
         .D(n32733), .Z(n8)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i15443_3_lut_rep_733_3_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .Z(n32748)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;
    defparam i15443_3_lut_rep_733_3_lut.init = 16'h7a7a;
    LUT4 i5216_2_lut_rep_609_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in[0]), .Z(n32624)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i5216_2_lut_rep_609_4_lut_4_lut.init = 16'h857a;
    LUT4 mux_3507_i4_3_lut (.A(n29853), .B(n34007), .C(n5651), .Z(n5659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3507_i4_3_lut.init = 16'hcaca;
    LUT4 i28594_2_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), .C(\alu_op[3] ), 
         .D(debug_rd_3__N_413), .Z(n30073)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i28594_2_lut_4_lut.init = 16'hff80;
    LUT4 i5245_2_lut_rep_610_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in[2]), .Z(n32625)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i5245_2_lut_rep_610_4_lut_4_lut.init = 16'h857a;
    LUT4 i5246_2_lut_rep_611_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in[3]), .Z(n32626)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i5246_2_lut_rep_611_4_lut_4_lut.init = 16'h857a;
    LUT4 i5244_2_lut_rep_631_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in[1]), .Z(n32646)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i5244_2_lut_rep_631_4_lut_4_lut.init = 16'h857a;
    LUT4 i1_2_lut_rep_734_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), .C(\alu_op[3] ), 
         .D(\alu_op[0] ), .Z(n32749)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;
    defparam i1_2_lut_rep_734_4_lut.init = 16'h7f00;
    LUT4 mux_327_i2_4_lut (.A(data_rs1_c[1]), .B(n32702), .C(n32704), 
         .D(mip_reg_c[17]), .Z(n809[1])) /* synthesis lut_function=(A (B)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(437[22:76])
    defparam mux_327_i2_4_lut.init = 16'hdc88;
    FD1P3AX tmp_data_i0_i1 (.D(tmp_data[5]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i1.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i2 (.D(tmp_data[6]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i2.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i3 (.D(tmp_data[7]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i3.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i4 (.D(tmp_data[8]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i4.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i5 (.D(tmp_data[9]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i5.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i6 (.D(tmp_data[10]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i6.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i7 (.D(tmp_data[11]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i7.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i8 (.D(tmp_data[12]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i8.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i9 (.D(tmp_data[13]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i9.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i10 (.D(tmp_data[14]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i10.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i11 (.D(tmp_data[15]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i11.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i12 (.D(tmp_data[16]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i12.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i13 (.D(tmp_data[17]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i13.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i14 (.D(tmp_data[18]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i14.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i15 (.D(tmp_data[19]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i15.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i16 (.D(tmp_data[20]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i16.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i17 (.D(tmp_data[21]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i17.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i18 (.D(tmp_data[22]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i18.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i19 (.D(tmp_data[23]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i19.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i20 (.D(tmp_data[24]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i20.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i21 (.D(tmp_data[25]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i21.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i22 (.D(tmp_data[26]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i22.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i23 (.D(tmp_data[27]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i23.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i24 (.D(tmp_data[28]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i24.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i25 (.D(tmp_data[29]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i25.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i26 (.D(tmp_data[30]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i26.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i27 (.D(tmp_data[31]), .SP(clk_c_enable_540), .CK(clk_c), 
            .Q(tmp_data[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i27.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i30 (.D(tmp_data_in[2]), .SP(clk_c_enable_540), 
            .CK(clk_c), .Q(tmp_data[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i30.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i31 (.D(tmp_data_in[3]), .SP(clk_c_enable_540), 
            .CK(clk_c), .Q(tmp_data[31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i31.GSR = "DISABLED";
    FD1P3AX mepc_i0_i1 (.D(mepc[5]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_735_3_lut (.A(counter_hi[2]), .B(counter_hi[4]), .C(counter_hi[3]), 
         .Z(n32750)) /* synthesis lut_function=(!(A (B+(C))+!A ((C)+!B))) */ ;
    defparam i1_2_lut_rep_735_3_lut.init = 16'h0606;
    FD1P3AX mepc_i0_i2 (.D(mepc[6]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i2.GSR = "DISABLED";
    FD1P3AX mepc_i0_i3 (.D(mepc[7]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i3.GSR = "DISABLED";
    FD1P3AX mepc_i0_i4 (.D(mepc[8]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i4.GSR = "DISABLED";
    FD1P3AX mepc_i0_i5 (.D(mepc[9]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i5.GSR = "DISABLED";
    FD1P3AX mepc_i0_i6 (.D(mepc[10]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i6.GSR = "DISABLED";
    FD1P3AX mepc_i0_i7 (.D(mepc[11]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i7.GSR = "DISABLED";
    FD1P3AX mepc_i0_i8 (.D(mepc[12]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i8.GSR = "DISABLED";
    FD1P3AX mepc_i0_i9 (.D(mepc[13]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i9.GSR = "DISABLED";
    FD1P3AX mepc_i0_i10 (.D(mepc[14]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i10.GSR = "DISABLED";
    FD1P3AX mepc_i0_i11 (.D(mepc[15]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i11.GSR = "DISABLED";
    FD1P3AX mepc_i0_i12 (.D(mepc[16]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i12.GSR = "DISABLED";
    FD1P3AX mepc_i0_i13 (.D(mepc[17]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i13.GSR = "DISABLED";
    FD1P3AX mepc_i0_i14 (.D(mepc[18]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i14.GSR = "DISABLED";
    FD1P3AX mepc_i0_i15 (.D(mepc[19]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i15.GSR = "DISABLED";
    FD1P3AX mepc_i0_i16 (.D(mepc[20]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i16.GSR = "DISABLED";
    FD1P3AX mepc_i0_i17 (.D(mepc[21]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i17.GSR = "DISABLED";
    FD1P3AX mepc_i0_i18 (.D(mepc[22]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i18.GSR = "DISABLED";
    FD1P3AX mepc_i0_i19 (.D(mepc[23]), .SP(clk_c_enable_538), .CK(clk_c), 
            .Q(mepc[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i19.GSR = "DISABLED";
    LUT4 i15333_3_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[4]), .C(mie[16]), 
         .D(mie[7]), .Z(n17982)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;
    defparam i15333_3_lut_4_lut.init = 16'hf960;
    FD1P3AX last_interrupt_req_i0_i1 (.D(\ui_in_sync[1] ), .SP(clk_c_enable_433), 
            .CK(clk_c), .Q(last_interrupt_req[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam last_interrupt_req_i0_i1.GSR = "DISABLED";
    FD1P3AX shift_amt__i2 (.D(n92[1]), .SP(clk_c_enable_436), .CK(clk_c), 
            .Q(shift_amt[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i2.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_adj_315 (.A(n32546), .B(n28275), .C(n32543), .D(n1), 
         .Z(n27427)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_315.init = 16'h4000;
    LUT4 i28282_2_lut_rep_800 (.A(counter_hi[3]), .B(counter_hi[4]), .Z(clk_c_enable_538)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i28282_2_lut_rep_800.init = 16'h7777;
    LUT4 i1_2_lut_3_lut_adj_316 (.A(counter_hi[3]), .B(counter_hi[4]), .C(\imm[6] ), 
         .Z(n26850)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_316.init = 16'h7070;
    LUT4 i28436_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), .C(rst_reg_n), 
         .Z(n11722)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam i28436_2_lut_3_lut.init = 16'h0707;
    LUT4 i15092_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), .C(mepc[0]), 
         .Z(csr_read_3__N_1451[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i15092_2_lut_3_lut.init = 16'h7070;
    LUT4 i27962_3_lut_4_lut (.A(\imm[10] ), .B(\imm[1] ), .C(n31618), 
         .D(n29875), .Z(n5652[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i27962_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i24425_2_lut_rep_801 (.A(\imm[10] ), .B(\imm[4] ), .Z(n32816)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24425_2_lut_rep_801.init = 16'heeee;
    FD1P3AX shift_amt__i3 (.D(n92[2]), .SP(clk_c_enable_436), .CK(clk_c), 
            .Q(shift_amt_adj_3153[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i3.GSR = "DISABLED";
    FD1P3AX shift_amt__i4 (.D(n92[3]), .SP(clk_c_enable_436), .CK(clk_c), 
            .Q(shift_amt_adj_3153[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i4.GSR = "DISABLED";
    FD1P3AX shift_amt__i5 (.D(n92[0]), .SP(clk_c_enable_437), .CK(clk_c), 
            .Q(shift_amt_adj_3153[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i5.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_317 (.A(\imm[10] ), .B(\imm[4] ), .C(\imm[7] ), 
         .D(\imm[11] ), .Z(n27962)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_317.init = 16'hfffe;
    LUT4 mux_3482_i3_4_lut_4_lut (.A(\imm[0] ), .B(\imm[1] ), .C(instrret_count[2]), 
         .D(cycle_count_wide[2]), .Z(n5607)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam mux_3482_i3_4_lut_4_lut.init = 16'h7340;
    LUT4 mux_3482_i4_4_lut_4_lut (.A(\imm[0] ), .B(\imm[1] ), .C(instrret_count[3]), 
         .D(\cycle_count_wide[3] ), .Z(n5605[3])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam mux_3482_i4_4_lut_4_lut.init = 16'h7340;
    LUT4 i5214_2_lut (.A(time_hi[0]), .B(clk_c_enable_276), .Z(n12[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam i5214_2_lut.init = 16'h6666;
    LUT4 i3_4_lut_rep_524_4_lut (.A(n32546), .B(n28343), .C(n32543), .D(n32559), 
         .Z(n32539)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i3_4_lut_rep_524_4_lut.init = 16'h4000;
    LUT4 i15070_2_lut (.A(data_rs2[0]), .B(data_out_3__N_1385), .Z(\data_out_slice[0] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i15070_2_lut.init = 16'h2222;
    LUT4 i15330_2_lut_rep_629 (.A(data_rs2[3]), .B(data_out_3__N_1385), 
         .Z(n32644)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i15330_2_lut_rep_629.init = 16'h2222;
    LUT4 i8336_4_lut (.A(mem_op[1]), .B(mem_op[0]), .C(n34281), .D(n34283), 
         .Z(data_out_3__N_1385)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[13] 272[50])
    defparam i8336_4_lut.init = 16'h5150;
    LUT4 mtimecmp_7__I_0_3_lut_4_lut (.A(data_rs2[3]), .B(data_out_3__N_1385), 
         .C(timer_data_3__N_631), .D(\mtimecmp[7] ), .Z(mtimecmp_3__N_1935)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam mtimecmp_7__I_0_3_lut_4_lut.init = 16'h2f20;
    LUT4 i1_3_lut_4_lut_adj_318 (.A(n32676), .B(\data_rs1[3] ), .C(n14), 
         .D(mie[15]), .Z(n25984)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_318.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_319 (.A(n32676), .B(\data_rs1[3] ), .C(n14), 
         .D(mie[16]), .Z(n25980)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_319.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_320 (.A(n32676), .B(\data_rs1[3] ), .C(n14), 
         .D(mie[11]), .Z(n25986)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_320.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_321 (.A(n32676), .B(\data_rs1[3] ), .C(n14), 
         .D(mie[7]), .Z(n25978)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_321.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_322 (.A(n32676), .B(\data_rs1[3] ), .C(n14), 
         .D(mie[3]), .Z(n25982)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_322.init = 16'h8f88;
    LUT4 mstatus_mie_I_153_3_lut_4_lut (.A(n32676), .B(\data_rs1[3] ), .C(n32724), 
         .D(mstatus_mpie), .Z(mstatus_mie_N_1709)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam mstatus_mie_I_153_3_lut_4_lut.init = 16'hf808;
    LUT4 mie_0__bdd_4_lut (.A(mie[0]), .B(\data_rs1[0] ), .C(n32704), 
         .D(n32702), .Z(n31292)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B (D))) */ ;
    defparam mie_0__bdd_4_lut.init = 16'hee2a;
    LUT4 i1_2_lut_rep_812 (.A(\imm[9] ), .B(\imm[8] ), .Z(n32827)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_812.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_323 (.A(\imm[9] ), .B(\imm[8] ), .C(n10687), 
         .D(n27962), .Z(n5651)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_323.init = 16'h0080;
    LUT4 i15327_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[31]), 
         .D(n32768), .Z(\addr_out[27] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i15327_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i15324_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[28]), 
         .D(n32768), .Z(\addr_out[24] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i15324_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i15325_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[29]), 
         .D(n32768), .Z(\addr_out[25] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i15325_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i15326_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[30]), 
         .D(n32768), .Z(\addr_out[26] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i15326_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 equal_3108_i3_2_lut_rep_814 (.A(cycle[0]), .B(cycle[1]), .Z(n32829)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(234[45:57])
    defparam equal_3108_i3_2_lut_rep_814.init = 16'heeee;
    PFUMX i28679 (.BLUT(n31428), .ALUT(n31425), .C0(n32772), .Z(debug_rd[2]));
    LUT4 i28489_2_lut_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(n32839), 
         .D(counter_hi[2]), .Z(clk_c_enable_437)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(234[45:57])
    defparam i28489_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i28451_2_lut_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(counter_hi[2]), 
         .D(n32839), .Z(clk_c_enable_436)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(234[45:57])
    defparam i28451_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_324 (.A(n29445), .B(\imm[9] ), .C(\imm[8] ), .D(n29443), 
         .Z(n10660)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_324.init = 16'hffbf;
    LUT4 i1_4_lut_adj_325 (.A(\imm[0] ), .B(\imm[10] ), .C(\imm[1] ), 
         .D(\imm[11] ), .Z(n29445)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_325.init = 16'hfffe;
    PFUMX i28676 (.BLUT(debug_branch_N_840[30]), .ALUT(n31426), .C0(n30171), 
          .Z(n31427));
    LUT4 i15547_2_lut_rep_816 (.A(\imm[5] ), .B(\imm[3] ), .Z(n32831)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15547_2_lut_rep_816.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_326 (.A(\imm[5] ), .B(\imm[3] ), .C(\imm[7] ), 
         .D(\imm[4] ), .Z(n29443)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_326.init = 16'hfffe;
    LUT4 i27025_2_lut_3_lut (.A(\imm[5] ), .B(\imm[3] ), .C(\imm[2] ), 
         .Z(n29669)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i27025_2_lut_3_lut.init = 16'hfefe;
    LUT4 i27004_2_lut_3_lut (.A(\imm[5] ), .B(\imm[3] ), .C(\imm[6] ), 
         .Z(n29647)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i27004_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_327 (.A(stall_core), .B(instr_complete_N_1647), .C(clk_c_enable_285), 
         .D(n28903), .Z(n27656)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_327.init = 16'h8000;
    LUT4 i1_4_lut_adj_328 (.A(stall_core), .B(instr_complete_N_1647), .C(clk_c_enable_285), 
         .D(n28909), .Z(n27655)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_328.init = 16'h8000;
    LUT4 n29838_bdd_3_lut_29035 (.A(n29838), .B(n234[1]), .C(n30172), 
         .Z(n31410)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n29838_bdd_3_lut_29035.init = 16'hacac;
    LUT4 i1_4_lut_adj_329 (.A(stall_core), .B(instr_complete_N_1647), .C(n28897), 
         .D(clk_c_enable_285), .Z(n27657)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_329.init = 16'h8000;
    LUT4 i1_4_lut_4_lut_adj_330 (.A(n32546), .B(n28533), .C(n32548), .D(clk_c_enable_524), 
         .Z(n2559)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_330.init = 16'hf400;
    LUT4 equal_111_i4_2_lut_rep_819 (.A(counter_hi[3]), .B(counter_hi[4]), 
         .Z(n32834)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(481[33:47])
    defparam equal_111_i4_2_lut_rep_819.init = 16'hbbbb;
    LUT4 equal_111_i5_2_lut_rep_745_3_lut (.A(n34283), .B(n34281), .C(counter_hi[2]), 
         .Z(n32760)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(481[33:47])
    defparam equal_111_i5_2_lut_rep_745_3_lut.init = 16'hfbfb;
    LUT4 i28423_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n32758), .D(counter_hi[2]), .Z(clk_c_enable_187)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(481[33:47])
    defparam i28423_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i28380_2_lut_rep_731_3_lut (.A(n34283), .B(n34281), .C(counter_hi[2]), 
         .Z(n32746)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(481[33:47])
    defparam i28380_2_lut_rep_731_3_lut.init = 16'h4040;
    LUT4 n31410_bdd_3_lut_28670 (.A(n31410), .B(n31409), .C(n32772), .Z(debug_rd_3__N_1392[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31410_bdd_3_lut_28670.init = 16'hcaca;
    LUT4 i1_4_lut_rep_523_4_lut (.A(n32546), .B(n28363), .C(n28483), .D(n32543), 
         .Z(n32538)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_rep_523_4_lut.init = 16'h4000;
    PFUMX i27143 (.BLUT(time_count[3]), .ALUT(n5605[3]), .C0(n32790), 
          .Z(n29852));
    LUT4 i1_4_lut_adj_331 (.A(n32829), .B(clk_c_enable_285), .C(n9909), 
         .D(n32828), .Z(address_ready)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_331.init = 16'h4000;
    LUT4 is_load_I_0_2_lut (.A(is_load), .B(is_store), .Z(n9909)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(237[58:79])
    defparam is_load_I_0_2_lut.init = 16'heeee;
    LUT4 i27038_3_lut_4_lut (.A(\alu_op[0] ), .B(n32732), .C(\data_rs1[0] ), 
         .D(n32733), .Z(n29683)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i27038_3_lut_4_lut.init = 16'hff80;
    FD1P3AX mstatus_mie_524 (.D(mstatus_mie_N_1707), .SP(clk_c_enable_520), 
            .CK(clk_c), .Q(mstatus_mie)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam mstatus_mie_524.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_824 (.A(n34283), .B(counter_hi[4]), .Z(n32839)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_2_lut_rep_824.init = 16'heeee;
    LUT4 i15093_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(mcause[4]), .D(counter_hi[2]), .Z(csr_read_3__N_1637[0])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i15093_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i20_3_lut_4_lut (.A(\alu_op[0] ), .B(n32732), .C(\data_rs1[3] ), 
         .D(n32733), .Z(n14)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i20_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_rep_750_3_lut (.A(n34283), .B(n34281), .C(counter_hi[2]), 
         .Z(n32765)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_2_lut_rep_750_3_lut.init = 16'hfefe;
    LUT4 n29882_bdd_3_lut (.A(n29882), .B(n29881), .C(\imm[1] ), .Z(n32349)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n29882_bdd_3_lut.init = 16'hacac;
    LUT4 equal_110_i5_2_lut_rep_744_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(n32759)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam equal_110_i5_2_lut_rep_744_3_lut.init = 16'hefef;
    LUT4 i28483_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_top_bit_next_N_1731), .D(counter_hi[2]), .Z(n18385)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i28483_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 equal_107_i6_1_lut_rep_703_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(clk_c_enable_363)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam equal_107_i6_1_lut_rep_703_2_lut_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_top_bit_next_N_1731), .D(counter_hi[2]), .Z(clk_c_enable_522)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i28345_2_lut_rep_695_3_lut_3_lut_4_lut_3_lut (.A(counter_hi[3]), 
         .B(counter_hi[4]), .C(counter_hi[2]), .Z(n32710)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i28345_2_lut_rep_695_3_lut_3_lut_4_lut_3_lut.init = 16'h0404;
    LUT4 n193_bdd_4_lut_29637 (.A(n191[2]), .B(shift_out[2]), .C(n32805), 
         .D(n32838), .Z(n31420)) /* synthesis lut_function=(A (B+((D)+!C))+!A !(((D)+!C)+!B)) */ ;
    defparam n193_bdd_4_lut_29637.init = 16'haaca;
    LUT4 i3935_2_lut_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(mstatus_mte), .D(counter_hi[2]), .Z(n6086)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i3935_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    FD1P3IX load_top_bit_513 (.D(\debug_branch_N_450[3] ), .SP(clk_c_enable_522), 
            .CD(n18385), .CK(clk_c), .Q(load_top_bit)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(156[12] 157[43])
    defparam load_top_bit_513.GSR = "DISABLED";
    LUT4 i15263_2_lut_rep_716_3_lut_4_lut (.A(n34283), .B(n34281), .C(cy_adj_3150), 
         .D(counter_hi[2]), .Z(n32731)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i15263_2_lut_rep_716_3_lut_4_lut.init = 16'hf0f1;
    PFUMX i30007 (.BLUT(n34276), .ALUT(n34277), .C0(n32730), .Z(n34278));
    PFUMX i28617 (.BLUT(n31292), .ALUT(n34292), .C0(n32733), .Z(n31293));
    LUT4 i27051_3_lut_3_lut (.A(counter_hi[4]), .B(n30425), .C(n13), .Z(n29760)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i27051_3_lut_3_lut.init = 16'he4e4;
    LUT4 i15328_2_lut_rep_653 (.A(data_rs2[1]), .B(data_out_3__N_1385), 
         .Z(n32668)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i15328_2_lut_rep_653.init = 16'h2222;
    LUT4 mtimecmp_5__I_0_3_lut_4_lut (.A(data_rs2[1]), .B(data_out_3__N_1385), 
         .C(timer_data_3__N_631), .D(\mtimecmp[5] ), .Z(mtimecmp_1__N_1941)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam mtimecmp_5__I_0_3_lut_4_lut.init = 16'h2f20;
    LUT4 i1_2_lut_rep_832 (.A(\alu_op[0] ), .B(\alu_op[1] ), .Z(n32847)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_2_lut_rep_832.init = 16'heeee;
    LUT4 i1_2_lut_rep_717_3_lut_4_lut_3_lut (.A(\alu_op[1] ), .B(debug_instr_valid), 
         .C(is_system), .Z(n32732)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_2_lut_rep_717_3_lut_4_lut_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_332 (.A(n10675), .B(n32736), .C(\debug_rd_3__N_405[28] ), 
         .D(interrupt_core), .Z(n27994)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_332.init = 16'h0004;
    LUT4 i25_4_lut (.A(n32736), .B(n32793), .C(interrupt_core), .D(n26807), 
         .Z(n26364)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(351[22] 355[16])
    defparam i25_4_lut.init = 16'hfaca;
    LUT4 is_system_I_0_2_lut_rep_833 (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .C(debug_instr_valid), .D(is_system), .Z(n32848)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam is_system_I_0_2_lut_rep_833.init = 16'he000;
    LUT4 i1_2_lut_rep_661_3_lut_4_lut_4_lut_3_lut_4_lut (.A(\alu_op[0] ), 
         .B(\alu_op[1] ), .C(debug_instr_valid), .D(is_system), .Z(n32676)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_2_lut_rep_661_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h6000;
    LUT4 i15561_2_lut_rep_834 (.A(\imm[8] ), .B(\imm[9] ), .Z(n32849)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15561_2_lut_rep_834.init = 16'heeee;
    LUT4 n29844_bdd_3_lut_29640 (.A(n29844), .B(n234[2]), .C(n30172), 
         .Z(n31423)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n29844_bdd_3_lut_29640.init = 16'hacac;
    LUT4 i1_4_lut_adj_333 (.A(n32678), .B(instr_complete_N_1648), .C(n17772), 
         .D(n11035), .Z(n17920)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(220[18] 228[36])
    defparam i1_4_lut_adj_333.init = 16'hffef;
    LUT4 i15124_2_lut (.A(cycle[0]), .B(cycle[1]), .Z(n17772)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15124_2_lut.init = 16'h8888;
    LUT4 i15077_2_lut_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), .C(n10675), 
         .D(n32768), .Z(n5080[0])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i15077_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 is_trap_I_0_586_2_lut_rep_676_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), 
         .C(interrupt_core), .D(n32768), .Z(n32691)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam is_trap_I_0_586_2_lut_rep_676_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i1_2_lut_rep_690_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), .C(interrupt_core), 
         .D(n32768), .Z(n32705)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i1_2_lut_rep_690_3_lut_4_lut.init = 16'hf1f0;
    FD1P3IX mepc_i0_i23 (.D(n658[3]), .SP(clk_c_enable_538), .CD(n11722), 
            .CK(clk_c), .Q(mepc[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i23.GSR = "DISABLED";
    FD1P3IX mepc_i0_i22 (.D(n658[2]), .SP(clk_c_enable_538), .CD(n11722), 
            .CK(clk_c), .Q(mepc[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i22.GSR = "DISABLED";
    FD1P3IX mepc_i0_i21 (.D(n658[1]), .SP(clk_c_enable_538), .CD(n11722), 
            .CK(clk_c), .Q(mepc[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i21.GSR = "DISABLED";
    LUT4 debug_branch_N_840_30__bdd_4_lut (.A(n31420), .B(n31419), .C(n15), 
         .D(n32807), .Z(n31425)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (B (D))) */ ;
    defparam debug_branch_N_840_30__bdd_4_lut.init = 16'hcca0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_334 (.A(n32765), .B(n32691), .C(n32675), 
         .D(n32724), .Z(clk_c_enable_115)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(398[22:52])
    defparam i1_2_lut_3_lut_4_lut_adj_334.init = 16'hfff4;
    LUT4 i7219_3_lut_rep_757_4_lut (.A(is_alu_imm), .B(is_alu_reg), .C(is_auipc), 
         .D(debug_instr_valid), .Z(n32772)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(225[22:46])
    defparam i7219_3_lut_rep_757_4_lut.init = 16'hfe00;
    LUT4 i5901_2_lut_3_lut (.A(is_alu_imm), .B(is_alu_reg), .C(debug_instr_valid), 
         .Z(debug_rd_3__N_1401)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(225[22:46])
    defparam i5901_2_lut_3_lut.init = 16'he0e0;
    FD1P3IX mepc_i0_i20 (.D(n658[0]), .SP(clk_c_enable_538), .CD(n11722), 
            .CK(clk_c), .Q(mepc[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i20.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_335 (.A(stall_core), .B(instr_complete_N_1647), .C(clk_c_enable_285), 
         .D(n28889), .Z(n27653)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_335.init = 16'h8000;
    LUT4 i28322_3_lut_4_lut (.A(n32736), .B(interrupt_core), .C(n32765), 
         .D(rst_reg_n), .Z(clk_c_enable_347)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i28322_3_lut_4_lut.init = 16'h0eff;
    FD1P3IX tmp_data_i0_i29 (.D(tmp_data_in_3__N_1514[1]), .SP(clk_c_enable_540), 
            .CD(n11720), .CK(clk_c), .Q(tmp_data[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i29.GSR = "DISABLED";
    FD1P3IX tmp_data_i0_i28 (.D(tmp_data_in_3__N_1514[0]), .SP(clk_c_enable_540), 
            .CD(n11720), .CK(clk_c), .Q(tmp_data[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i28.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_839 (.A(counter_hi[2]), .B(n34283), .Z(n32854)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i1_2_lut_rep_839.init = 16'h8888;
    FD1S3IX instr_retired_518 (.D(instr_complete_N_1647), .CK(clk_c), .CD(n18087), 
            .Q(instr_retired)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(303[12] 305[8])
    defparam instr_retired_518.GSR = "DISABLED";
    PFUMX i28666 (.BLUT(n31408), .ALUT(n31406), .C0(n32807), .Z(n31409));
    FD1S3AX cycle__i0 (.D(n31351), .CK(clk_c), .Q(cycle[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam cycle__i0.GSR = "DISABLED";
    LUT4 debug_branch_N_840_30__bdd_3_lut (.A(n29864), .B(data_out_3__N_1385), 
         .C(load_top_bit), .Z(n31426)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam debug_branch_N_840_30__bdd_3_lut.init = 16'he2e2;
    LUT4 i15715_2_lut_rep_755_3_lut (.A(counter_hi[2]), .B(n34283), .C(n34281), 
         .Z(clk_c_enable_285)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i15715_2_lut_rep_755_3_lut.init = 16'h8080;
    LUT4 i28404_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), 
         .C(n32758), .D(counter_hi[4]), .Z(clk_c_enable_195)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i28404_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i13_4_lut_3_lut (.A(counter_hi[2]), .B(counter_hi[3]), .C(counter_hi[4]), 
         .Z(csr_read_3__N_1443[2])) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i13_4_lut_3_lut.init = 16'h8181;
    LUT4 i21720_2_lut_3_lut (.A(counter_hi[2]), .B(counter_hi[3]), .C(counter_hi[4]), 
         .Z(n18)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i21720_2_lut_3_lut.init = 16'h7878;
    LUT4 i1_4_lut_adj_336 (.A(n29317), .B(n32724), .C(n131), .D(n29671), 
         .Z(clk_c_enable_55)) /* synthesis lut_function=(A+!(B+((D)+!C))) */ ;
    defparam i1_4_lut_adj_336.init = 16'haaba;
    LUT4 i14867_4_lut (.A(n32647), .B(n32650), .C(mstatus_mie), .D(n32670), 
         .Z(n6299)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam i14867_4_lut.init = 16'h3022;
    LUT4 i28273_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), 
         .C(rst_reg_n), .D(counter_hi[4]), .Z(clk_c_enable_28)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i28273_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i24607_rep_537_3_lut_4_lut (.A(counter_hi[2]), .B(n34283), .C(n27294), 
         .D(n34281), .Z(n32552)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i24607_rep_537_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_337 (.A(counter_hi[2]), .B(counter_hi[3]), 
         .C(mcause[5]), .D(counter_hi[4]), .Z(n29227)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i1_2_lut_3_lut_4_lut_adj_337.init = 16'h8000;
    LUT4 i1_2_lut_rep_693_3_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), 
         .C(n32783), .D(counter_hi[4]), .Z(n32708)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i1_2_lut_rep_693_3_lut_4_lut.init = 16'h0800;
    LUT4 i24607_rep_142_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), 
         .C(n27294), .D(counter_hi[4]), .Z(n30928)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i24607_rep_142_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i24607_rep_141_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), 
         .C(n27294), .D(counter_hi[4]), .Z(n30927)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i24607_rep_141_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i24607_rep_140_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), 
         .C(n27294), .D(counter_hi[4]), .Z(n30926)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i24607_rep_140_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 n31423_bdd_3_lut (.A(n31423), .B(n31427), .C(debug_rd_3__N_1575), 
         .Z(n31428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31423_bdd_3_lut.init = 16'hcaca;
    LUT4 i24607_rep_139_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), 
         .C(n27294), .D(counter_hi[4]), .Z(n30925)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i24607_rep_139_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i24607_rep_138_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), 
         .C(n27294), .D(counter_hi[4]), .Z(n30924)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i24607_rep_138_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_3_lut_rep_759_4_lut (.A(counter_hi[2]), .B(n34283), .C(n34285), 
         .D(n34281), .Z(n32774)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(439[18] 459[12])
    defparam i1_3_lut_rep_759_4_lut.init = 16'hf7ff;
    LUT4 i1_4_lut_adj_338 (.A(\imm[1] ), .B(n32831), .C(\imm[0] ), .D(\imm[2] ), 
         .Z(n10687)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_adj_338.init = 16'h0110;
    LUT4 data_rs1_3__I_0_i1_2_lut (.A(\data_rs1[0] ), .B(cycle[0]), .Z(mul_out_3__N_1510[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i1_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i2_2_lut (.A(data_rs1_c[1]), .B(cycle[0]), .Z(mul_out_3__N_1510[1])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i2_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i3_2_lut (.A(data_rs1[2]), .B(cycle[0]), .Z(mul_out_3__N_1510[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i3_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i4_2_lut (.A(\data_rs1[3] ), .B(cycle[0]), .Z(mul_out_3__N_1510[3])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i4_2_lut.init = 16'h8888;
    LUT4 i2_2_lut_3_lut_4_lut (.A(\imm[2] ), .B(n32703), .C(n32746), .D(n32759), 
         .Z(clk_c_enable_332)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_339 (.A(\imm[2] ), .B(n32703), .C(clk_c_enable_285), 
         .D(n32759), .Z(clk_c_enable_316)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_2_lut_3_lut_4_lut_adj_339.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_340 (.A(\imm[2] ), .B(n32703), .C(n32760), 
         .D(n32759), .Z(clk_c_enable_335)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_2_lut_3_lut_4_lut_adj_340.init = 16'h0200;
    LUT4 i1_3_lut_4_lut_adj_341 (.A(n32705), .B(n32769), .C(n11035), .D(instr_complete_N_1648), 
         .Z(instr_complete_N_1647)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i1_3_lut_4_lut_adj_341.init = 16'hfffe;
    LUT4 i1_4_lut_adj_342 (.A(n27962), .B(n32733), .C(n29669), .D(n29425), 
         .Z(n652)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_342.init = 16'h0400;
    LUT4 i1_4_lut_adj_343 (.A(\imm[1] ), .B(\imm[0] ), .C(n32827), .D(\imm[6] ), 
         .Z(n29425)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_343.init = 16'h4000;
    LUT4 i15339_4_lut (.A(\data_rs1[3] ), .B(n32807), .C(\debug_branch_N_442[31] ), 
         .D(n32806), .Z(alu_a_in[3])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i15339_4_lut.init = 16'h3022;
    LUT4 i15338_4_lut (.A(data_rs1[2]), .B(n32807), .C(\debug_branch_N_442[30] ), 
         .D(n32806), .Z(alu_a_in[2])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i15338_4_lut.init = 16'h3022;
    LUT4 imm_3__I_0_i3_3_lut (.A(\debug_rd_3__N_405[30] ), .B(data_rs2[2]), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 i15337_4_lut (.A(data_rs1_c[1]), .B(n32807), .C(\debug_branch_N_442[29] ), 
         .D(n32806), .Z(alu_a_in[1])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i15337_4_lut.init = 16'h3022;
    LUT4 n31443_bdd_3_lut_4_lut (.A(n32710), .B(mip_reg[16]), .C(\imm[6] ), 
         .D(n32883), .Z(n32347)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n31443_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_4_lut_adj_344 (.A(stall_core), .B(clk_c_enable_285), .C(n32783), 
         .D(\addr_offset[2] ), .Z(n28963)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_344.init = 16'h8000;
    LUT4 imm_3__I_0_i2_3_lut (.A(\debug_rd_3__N_405[29] ), .B(data_rs2[1]), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 imm_3__I_0_i1_3_lut (.A(\debug_rd_3__N_405[28] ), .B(data_rs2[0]), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 i5882_3_lut (.A(n34285), .B(is_alu_reg), .C(is_branch), .Z(alu_b_in_3__N_1504)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:52])
    defparam i5882_3_lut.init = 16'ha8a8;
    LUT4 i15094_4_lut (.A(n157), .B(n32807), .C(\debug_branch_N_442[28] ), 
         .D(n30051), .Z(alu_a_in[0])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i15094_4_lut.init = 16'h2230;
    LUT4 i1_4_lut_4_lut_adj_345 (.A(n32546), .B(n28495), .C(n32548), .D(clk_c_enable_524), 
         .Z(n2124)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_345.init = 16'hf400;
    LUT4 imm_3__I_0_i4_3_lut (.A(\debug_rd_3__N_405[31] ), .B(data_rs2[3]), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 i4392_2_lut_4_lut (.A(tmp_data[6]), .B(mepc[2]), .C(n32724), 
         .D(\addr_offset[2] ), .Z(n701)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(267[23:65])
    defparam i4392_2_lut_4_lut.init = 16'h35ca;
    LUT4 i1_2_lut_rep_630_3_lut_4_lut (.A(n32736), .B(interrupt_core), .C(n32724), 
         .D(n32765), .Z(n32645)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i1_2_lut_rep_630_3_lut_4_lut.init = 16'hf0fe;
    LUT4 mux_252_i4_3_lut_4_lut (.A(n32736), .B(interrupt_core), .C(\debug_branch_N_442[31] ), 
         .D(n653[3]), .Z(n658[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15080_2_lut_3_lut_4_lut (.A(n32736), .B(interrupt_core), .C(n32675), 
         .D(n32765), .Z(mstatus_mte_N_1703)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i15080_2_lut_3_lut_4_lut.init = 16'hfff1;
    LUT4 mux_252_i3_3_lut_4_lut (.A(n32736), .B(interrupt_core), .C(\debug_branch_N_442[30] ), 
         .D(n653[2]), .Z(n658[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i2_3_lut_4_lut (.A(n32736), .B(interrupt_core), .C(\debug_branch_N_442[29] ), 
         .D(n653[1]), .Z(n658[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n30235_bdd_4_lut_28689 (.A(n32759), .B(csr_read_3__N_1451[0]), 
         .C(csr_read_3__N_1443[2]), .D(\imm[6] ), .Z(n31441)) /* synthesis lut_function=(A (B (D))+!A (B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n30235_bdd_4_lut_28689.init = 16'hcc05;
    LUT4 i15329_2_lut (.A(data_rs2[2]), .B(data_out_3__N_1385), .Z(\data_out_slice[2] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i15329_2_lut.init = 16'h2222;
    LUT4 is_double_fault_I_0_3_lut_rep_660_4_lut (.A(n32765), .B(n32736), 
         .C(is_double_fault_r), .D(mstatus_mte), .Z(n32675)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam is_double_fault_I_0_3_lut_rep_660_4_lut.init = 16'hf0f4;
    LUT4 i1_3_lut_adj_346 (.A(\debug_rd_3__N_405[30] ), .B(\debug_rd_3__N_405[29] ), 
         .C(\debug_rd_3__N_405[31] ), .Z(n10675)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(353[26:40])
    defparam i1_3_lut_adj_346.init = 16'hfefe;
    LUT4 i2_3_lut_rep_531 (.A(n32783), .B(debug_early_branch_N_955), .C(no_write_in_progress), 
         .Z(n32546)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i2_3_lut_rep_531.init = 16'h4040;
    LUT4 i1_3_lut_rep_684 (.A(n10660), .B(n24384), .C(\imm[2] ), .Z(n32699)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i1_3_lut_rep_684.init = 16'hbfbf;
    LUT4 i790_2_lut_4_lut (.A(n10660), .B(n24384), .C(\imm[2] ), .D(n32760), 
         .Z(n1152)) /* synthesis lut_function=(!(A (D)+!A (B (C+(D))+!B (D)))) */ ;
    defparam i790_2_lut_4_lut.init = 16'h00bf;
    LUT4 i27166_3_lut (.A(cycle_count_wide[1]), .B(time_count[1]), .C(\imm[0] ), 
         .Z(n29875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27166_3_lut.init = 16'hcaca;
    LUT4 mux_3503_i2_4_lut (.A(n31545), .B(mepc[1]), .C(\imm[0] ), .D(n26850), 
         .Z(n5646[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3503_i2_4_lut.init = 16'hca0a;
    PFUMX debug_rd_3__I_122_i4 (.BLUT(debug_rd_3__N_1571[3]), .ALUT(debug_rd_3__N_1396[3]), 
          .C0(n32772), .Z(debug_rd_3__N_1392[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    L6MUX21 instr_complete_I_131 (.D0(instr_complete_N_1650), .D1(instr_complete_N_1649), 
            .SD(n30073), .Z(instr_complete_N_1648)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX instr_complete_I_132 (.BLUT(instr_complete_N_1654), .ALUT(instr_complete_N_1656), 
          .C0(debug_rd_3__N_413), .Z(instr_complete_N_1649)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 mux_149_i1_3_lut_4_lut (.A(n32829), .B(n32747), .C(alu_out[0]), 
         .D(data_rs2[0]), .Z(tmp_data_in_3__N_1582[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_149_i2_3_lut_4_lut (.A(n32829), .B(n32747), .C(alu_out[1]), 
         .D(data_rs2[1]), .Z(tmp_data_in_3__N_1582[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_149_i4_3_lut_4_lut (.A(n32829), .B(n32747), .C(alu_out[3]), 
         .D(data_rs2[3]), .Z(tmp_data_in_3__N_1582[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_149_i3_3_lut_4_lut (.A(n32829), .B(n32747), .C(alu_out[2]), 
         .D(data_rs2[2]), .Z(tmp_data_in_3__N_1582[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i3_3_lut_4_lut.init = 16'hfb40;
    PFUMX tmp_data_in_3__I_0_i4 (.BLUT(tmp_data_in_3__N_1582[3]), .ALUT(tmp_data_in_3__N_1514[3]), 
          .C0(n30193), .Z(tmp_data_in[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_4_lut_adj_347 (.A(n32816), .B(n10687), .C(n32827), .D(n27960), 
         .Z(n27933)) /* synthesis lut_function=(!(A+!(B (C)+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_adj_347.init = 16'h4050;
    L6MUX21 debug_rd_3__I_122_i1 (.D0(debug_rd_3__N_1567[0]), .D1(debug_rd_3__N_1571[0]), 
            .SD(debug_rd_3__N_1575), .Z(debug_rd_3__N_1392[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_rep_534_4_lut (.A(clk_c_enable_285), .B(n32783), .C(instr_complete_N_1647), 
         .D(stall_core), .Z(n32549)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_rep_534_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_adj_348 (.A(clk_c_enable_285), .B(n32783), .C(stall_core), 
         .D(\next_pc_offset[3] ), .Z(n28237)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_4_lut_adj_348.init = 16'h2000;
    LUT4 mux_3113_i2_4_lut_4_lut (.A(n32759), .B(n32765), .C(mstatus_mpie), 
         .D(mstatus_mie), .Z(csr_read_3__N_1439[3])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(471[33:47])
    defparam mux_3113_i2_4_lut_4_lut.init = 16'h7340;
    PFUMX tmp_data_in_3__I_0_i3 (.BLUT(tmp_data_in_3__N_1582[2]), .ALUT(tmp_data_in_3__N_1514[2]), 
          .C0(n30193), .Z(tmp_data_in[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 csr_read_3__I_128_i4_4_lut (.A(mcause[3]), .B(n29227), .C(n32765), 
         .D(n32759), .Z(csr_read_3__N_1455[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(490[33] 493[57])
    defparam csr_read_3__I_128_i4_4_lut.init = 16'hca0a;
    PFUMX mux_87_i1 (.BLUT(debug_branch_N_840[28]), .ALUT(\debug_branch_N_450[0] ), 
          .C0(n30171), .Z(debug_rd_3__N_1571[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i27158_4_lut (.A(csr_read_3__N_1443[2]), .B(mepc[2]), .C(\imm[6] ), 
         .D(clk_c_enable_538), .Z(n29867)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i27158_4_lut.init = 16'hca0a;
    PFUMX i29867 (.BLUT(n34006), .ALUT(n34002), .C0(\imm[0] ), .Z(n34007));
    LUT4 i15286_4_lut (.A(mcause[0]), .B(\imm[1] ), .C(csr_read_3__N_1637[0]), 
         .D(n32765), .Z(n5632[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i15286_4_lut.init = 16'hc088;
    PFUMX i29865 (.BLUT(n34004), .ALUT(n34003), .C0(counter_hi[3]), .Z(n34005));
    LUT4 i1_4_lut_adj_349 (.A(n32792), .B(n27723), .C(n32793), .D(n32794), 
         .Z(n27861)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(331[17] 350[24])
    defparam i1_4_lut_adj_349.init = 16'hfdfc;
    LUT4 i1_4_lut_adj_350 (.A(n18098), .B(debug_rd_3__N_1575), .C(mem_op[1]), 
         .D(mem_op[2]), .Z(load_top_bit_next_N_1731)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_350.init = 16'h0004;
    LUT4 i27172_3_lut (.A(cycle_count_wide[0]), .B(\cycle_count_wide[3] ), 
         .C(\imm[0] ), .Z(n29881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27172_3_lut.init = 16'hcaca;
    PFUMX mux_93_i1 (.BLUT(\debug_branch_N_446[28] ), .ALUT(n238), .C0(n30070), 
          .Z(debug_rd_3__N_1567[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX debug_rd_3__I_121_i1 (.BLUT(shift_out[0]), .ALUT(debug_rd_3__N_1559[0]), 
          .C0(n30243), .Z(debug_rd_3__N_1396[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i4753_2_lut_4_lut_4_lut (.A(n32765), .B(instrret_count[0]), .C(instr_retired), 
         .D(cy_c), .Z(increment_result_3__N_1925[0])) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i4753_2_lut_4_lut_4_lut.init = 16'h369c;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n32765), .B(alu_b_in[0]), .C(n32748), 
         .D(cy_adj_3149), .Z(n29121)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hc66c;
    LUT4 i4755_2_lut_rep_650_4_lut_4_lut (.A(n32765), .B(instrret_count[0]), 
         .C(instr_retired), .D(cy_c), .Z(n32665)) /* synthesis lut_function=(A (B (D))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i4755_2_lut_rep_650_4_lut_4_lut.init = 16'hc840;
    LUT4 i1_4_lut_adj_351 (.A(interrupt_pending_N_1671), .B(instr_complete_N_1647), 
         .C(clk_c_enable_285), .D(mstatus_mie), .Z(debug_early_branch_N_955)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_351.init = 16'h8000;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n32765), .B(cmp), .C(alu_b_in[1]), .D(alu_a_in[1]), 
         .Z(n28225)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd00d;
    LUT4 i1_4_lut_adj_352 (.A(n76), .B(n10727), .C(n29011), .D(n32792), 
         .Z(interrupt_pending_N_1671)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[47:59])
    defparam i1_4_lut_adj_352.init = 16'hfffe;
    LUT4 i4701_2_lut_rep_577_3_lut_4_lut_4_lut (.A(n32765), .B(alu_b_in[0]), 
         .C(n32748), .D(cy_adj_3149), .Z(n32592)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i4701_2_lut_rep_577_3_lut_4_lut_4_lut.init = 16'h3810;
    LUT4 i4836_2_lut_rep_648_4_lut_4_lut (.A(n32765), .B(\mtime_out[0] ), 
         .C(n32717), .D(cy), .Z(n32663)) /* synthesis lut_function=(A (B (D))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i4836_2_lut_rep_648_4_lut_4_lut.init = 16'hc840;
    LUT4 debug_rd_3__N_1575_bdd_4_lut_29201 (.A(\alu_op[3] ), .B(\alu_op[1] ), 
         .C(\alu_op_in[2] ), .D(cycle[0]), .Z(n32352)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam debug_rd_3__N_1575_bdd_4_lut_29201.init = 16'hfff7;
    LUT4 debug_rd_3__N_1575_bdd_4_lut_29351 (.A(n32848), .B(n32784), .C(debug_instr_valid), 
         .D(is_lui), .Z(n32353)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam debug_rd_3__N_1575_bdd_4_lut_29351.init = 16'hfaea;
    LUT4 i15579_4_lut_4_lut (.A(n32765), .B(\imm[1] ), .C(mcause[2]), 
         .D(mstatus_mte), .Z(n9620)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i15579_4_lut_4_lut.init = 16'h5140;
    LUT4 tmp_data_in_3__I_124_i4_4_lut_4_lut_4_lut (.A(n32765), .B(\data_rs1[3] ), 
         .C(interrupt_core), .D(n32736), .Z(tmp_data_in_3__N_1514[3])) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam tmp_data_in_3__I_124_i4_4_lut_4_lut_4_lut.init = 16'h505c;
    LUT4 cy_I_0_3_lut_rep_665_4_lut_4_lut (.A(n32765), .B(cy), .C(time_pulse_r), 
         .D(n10737), .Z(n32680)) /* synthesis lut_function=(A (B)+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam cy_I_0_3_lut_rep_665_4_lut_4_lut.init = 16'hd8dd;
    LUT4 debug_branch_N_446_31__bdd_3_lut (.A(\next_pc_for_core[7] ), .B(\next_pc_for_core[3] ), 
         .C(counter_hi[2]), .Z(n33042)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam debug_branch_N_446_31__bdd_3_lut.init = 16'hacac;
    LUT4 next_pc_for_core_23__bdd_4_lut (.A(\next_pc_for_core[23] ), .B(\next_pc_for_core[19] ), 
         .C(counter_hi[3]), .D(counter_hi[2]), .Z(n33039)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam next_pc_for_core_23__bdd_4_lut.init = 16'h0a0c;
    LUT4 i1_4_lut_adj_353 (.A(n32831), .B(n7739), .C(\imm[0] ), .D(\imm[2] ), 
         .Z(n27960)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_353.init = 16'hfffe;
    LUT4 i5176_2_lut (.A(\imm[6] ), .B(\imm[1] ), .Z(n7739)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5176_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_354 (.A(fsm_state[2]), .B(n32791), .C(fsm_state[0]), 
         .D(mie[3]), .Z(n10727)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_354.init = 16'h0100;
    LUT4 i67_4_lut (.A(n17891), .B(n32827), .C(\imm[4] ), .D(n32849), 
         .Z(n40)) /* synthesis lut_function=(A (B (C))+!A !(C+(D))) */ ;
    defparam i67_4_lut.init = 16'h8085;
    LUT4 i15242_2_lut (.A(\imm[1] ), .B(\imm[0] ), .Z(n17891)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15242_2_lut.init = 16'h8888;
    LUT4 i4513_3_lut (.A(time_hi[2]), .B(time_hi[1]), .C(time_hi[0]), 
         .Z(n498[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(295[55:71])
    defparam i4513_3_lut.init = 16'h6a6a;
    LUT4 i4506_2_lut (.A(time_hi[1]), .B(time_hi[0]), .Z(n498[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(295[55:71])
    defparam i4506_2_lut.init = 16'h6666;
    LUT4 tmp_data_31__I_0_542_i2_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[1]), 
         .D(tmp_data[5]), .Z(\addr_out[1] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i1_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[0]), 
         .D(tmp_data[4]), .Z(\addr_out[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i3_3_lut_rep_675_4_lut (.A(n32827), .B(n32768), 
         .C(mepc[2]), .D(tmp_data[6]), .Z(n32690)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i3_3_lut_rep_675_4_lut.init = 16'hf780;
    LUT4 n32353_bdd_2_lut (.A(n32353), .B(debug_rd_3__N_1575), .Z(n32354)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n32353_bdd_2_lut.init = 16'heeee;
    LUT4 tmp_data_31__I_0_542_i24_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[23]), 
         .D(tmp_data[27]), .Z(\addr_out[23] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i23_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[22]), 
         .D(tmp_data[26]), .Z(\addr_out[22] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i22_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[21]), 
         .D(tmp_data[25]), .Z(\addr_out[21] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i21_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[20]), 
         .D(tmp_data[24]), .Z(\addr_out[20] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i20_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[19]), 
         .D(tmp_data[23]), .Z(\addr_out[19] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i19_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[18]), 
         .D(tmp_data[22]), .Z(\addr_out[18] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i18_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[17]), 
         .D(tmp_data[21]), .Z(\addr_out[17] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i17_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[16]), 
         .D(tmp_data[20]), .Z(\addr_out[16] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i16_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[15]), 
         .D(tmp_data[19]), .Z(\addr_out[15] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i15_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[14]), 
         .D(tmp_data[18]), .Z(\addr_out[14] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i14_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[13]), 
         .D(tmp_data[17]), .Z(\addr_out[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i13_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[12]), 
         .D(tmp_data[16]), .Z(\addr_out[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i12_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[11]), 
         .D(tmp_data[15]), .Z(\addr_out[11] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i11_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[10]), 
         .D(tmp_data[14]), .Z(\addr_out[10] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i10_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[9]), 
         .D(tmp_data[13]), .Z(\addr_out[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i9_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[8]), 
         .D(tmp_data[12]), .Z(\addr_out[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i8_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[7]), 
         .D(tmp_data[11]), .Z(\addr_out[7] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i7_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[6]), 
         .D(tmp_data[10]), .Z(\addr_out[6] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i6_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[5]), 
         .D(tmp_data[9]), .Z(\addr_out[5] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i5_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[4]), 
         .D(tmp_data[8]), .Z(\addr_out[4] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i4_3_lut_4_lut (.A(n32827), .B(n32768), .C(mepc[3]), 
         .D(tmp_data[7]), .Z(\addr_out[3] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_355 (.A(n32733), .B(n32702), .C(n32704), .D(data_rs1_c[1]), 
         .Z(n57)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[25:55])
    defparam i1_4_lut_adj_355.init = 16'h4555;
    LUT4 n4841_bdd_3_lut (.A(n4826[1]), .B(counter_hi[2]), .C(mie[9]), 
         .Z(n31542)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n4841_bdd_3_lut.init = 16'hb8b8;
    LUT4 mux_328_i2_3_lut_4_lut (.A(n32848), .B(n32838), .C(data_rs1_c[1]), 
         .D(n809[1]), .Z(n812[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[25:55])
    defparam mux_328_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_251_i1_3_lut (.A(mepc[0]), .B(\data_rs1[0] ), .C(n652), .Z(n653[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i1_3_lut.init = 16'hcaca;
    LUT4 tmp_data_in_3__N_1581_I_0_588_2_lut_rep_655_3_lut_4_lut (.A(n32849), 
         .B(n32768), .C(n32765), .D(interrupt_core), .Z(n32670)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C)+!B (C+!(D))))) */ ;
    defparam tmp_data_in_3__N_1581_I_0_588_2_lut_rep_655_3_lut_4_lut.init = 16'h0f04;
    LUT4 n4841_bdd_2_lut_28730 (.A(counter_hi[2]), .B(mie[1]), .Z(n31541)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam n4841_bdd_2_lut_28730.init = 16'h4444;
    LUT4 i9012_2_lut_3_lut_4_lut (.A(n32849), .B(n32768), .C(clk_c_enable_540), 
         .D(interrupt_core), .Z(n11720)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i9012_2_lut_3_lut_4_lut.init = 16'hf040;
    LUT4 i28554_2_lut_3_lut_4_lut (.A(n32849), .B(n32768), .C(n5721), 
         .D(interrupt_core), .Z(n30193)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i28554_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 debug_rd_3__I_0_i4_4_lut (.A(debug_rd_3__N_1567[3]), .B(debug_rd_3__N_1392[3]), 
         .C(n32772), .D(debug_rd_3__N_1575), .Z(debug_rd[3])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(176[18] 194[12])
    defparam debug_rd_3__I_0_i4_4_lut.init = 16'hccca;
    PFUMX i28775 (.BLUT(n31617), .ALUT(n31616), .C0(\imm[10] ), .Z(n31618));
    LUT4 i1_3_lut_4_lut_adj_356 (.A(n32792), .B(n32794), .C(n76), .D(n10727), 
         .Z(n27723)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_356.init = 16'h0100;
    LUT4 i1_3_lut_4_lut_adj_357 (.A(n32792), .B(n32794), .C(n76), .D(n10727), 
         .Z(n26807)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_357.init = 16'h1110;
    LUT4 n13_bdd_3_lut_29175 (.A(\mem_data_from_read[17] ), .B(counter_hi[2]), 
         .C(\mem_data_from_read[21] ), .Z(n32308)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n13_bdd_3_lut_29175.init = 16'he2e2;
    LUT4 mux_251_i4_3_lut (.A(mepc[3]), .B(\data_rs1[3] ), .C(n652), .Z(n653[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i4_3_lut.init = 16'hcaca;
    LUT4 n32310_bdd_3_lut (.A(n32310), .B(\timer_data[1] ), .C(is_timer_addr), 
         .Z(n32311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n32310_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_251_i3_3_lut (.A(mepc[2]), .B(data_rs1[2]), .C(n652), .Z(n653[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i3_3_lut.init = 16'hcaca;
    LUT4 mux_251_i2_3_lut (.A(mepc[1]), .B(data_rs1_c[1]), .C(n652), .Z(n653[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_rep_533 (.A(stall_core), .B(instr_complete_N_1647), .C(clk_c_enable_285), 
         .D(n32783), .Z(n32548)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_rep_533.init = 16'h8000;
    LUT4 dr_3__N_1864_31__bdd_3_lut_29227_4_lut (.A(\alu_op[3] ), .B(n32804), 
         .C(\mul_out[3] ), .D(alu_out[3]), .Z(n32401)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam dr_3__N_1864_31__bdd_3_lut_29227_4_lut.init = 16'hfd20;
    LUT4 i15067_3_lut_4_lut (.A(\alu_op[3] ), .B(n32804), .C(n32838), 
         .D(n32805), .Z(clk_c_enable_540)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam i15067_3_lut_4_lut.init = 16'hd0ff;
    LUT4 mux_72_i3_3_lut_4_lut (.A(\alu_op[3] ), .B(n32804), .C(alu_out[2]), 
         .D(\mul_out[2] ), .Z(n191[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam mux_72_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i1_4_lut_adj_358 (.A(rd[3]), .B(n32783), .C(rd[2]), .D(n32776), 
         .Z(n28897)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_358.init = 16'h4888;
    LUT4 mux_72_i2_3_lut_4_lut (.A(\alu_op[3] ), .B(n32804), .C(alu_out[1]), 
         .D(\mul_out[1] ), .Z(n191[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam mux_72_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 tmp_data_in_3__I_124_i2_3_lut (.A(tmp_data_in_3__N_1582[1]), .B(data_rs1_c[1]), 
         .C(n5721), .Z(tmp_data_in_3__N_1514[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_124_i2_3_lut.init = 16'hcaca;
    LUT4 n31760_bdd_3_lut_4_lut (.A(n32807), .B(\alu_op[0] ), .C(n31758), 
         .D(n31760), .Z(cmp_out)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam n31760_bdd_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_3024_i2_3_lut_4_lut (.A(n32807), .B(\alu_op[0] ), .C(alu_b_in[1]), 
         .D(alu_a_in[1]), .Z(n4901[1])) /* synthesis lut_function=(A (C+(D))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam mux_3024_i2_3_lut_4_lut.init = 16'hfbb0;
    LUT4 i12470_4_lut (.A(\alu_op[0] ), .B(\alu_op[3] ), .C(\alu_op[1] ), 
         .D(\alu_op_in[2] ), .Z(n5721)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    defparam i12470_4_lut.init = 16'hca0a;
    LUT4 mux_3024_i3_3_lut_4_lut (.A(n32807), .B(\alu_op[0] ), .C(alu_b_in[2]), 
         .D(alu_a_in[2]), .Z(n4901[2])) /* synthesis lut_function=(A (C+(D))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam mux_3024_i3_3_lut_4_lut.init = 16'hfbb0;
    LUT4 mux_3024_i4_3_lut_4_lut (.A(n32807), .B(\alu_op[0] ), .C(alu_b_in[3]), 
         .D(alu_a_in[3]), .Z(n4901[3])) /* synthesis lut_function=(A (C+(D))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam mux_3024_i4_3_lut_4_lut.init = 16'hfbb0;
    LUT4 mux_3024_i1_3_lut_4_lut (.A(n32807), .B(\alu_op[0] ), .C(alu_b_in[0]), 
         .D(alu_a_in[0]), .Z(n4901[0])) /* synthesis lut_function=(A (C+(D))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam mux_3024_i1_3_lut_4_lut.init = 16'hfbb0;
    LUT4 tmp_data_in_3__I_124_i1_3_lut (.A(tmp_data_in_3__N_1582[0]), .B(\data_rs1[0] ), 
         .C(n5721), .Z(tmp_data_in_3__N_1514[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_124_i1_3_lut.init = 16'hcaca;
    L6MUX21 i29408 (.D0(n33043), .D1(n33041), .SD(n30172), .Z(debug_rd_3__N_1567[3]));
    PFUMX i29406 (.BLUT(n33042), .ALUT(\debug_branch_N_446[31] ), .C0(n30175), 
          .Z(n33043));
    PFUMX i29404 (.BLUT(n33040), .ALUT(n33039), .C0(counter_hi[4]), .Z(n33041));
    PFUMX mux_91_i3 (.BLUT(n29842), .ALUT(\debug_branch_N_446[30] ), .C0(n30175), 
          .Z(n234[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_adj_359 (.A(n32783), .B(rd[1]), .C(rd[0]), .Z(n28903)) /* synthesis lut_function=(!((B (C)+!B !(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_adj_359.init = 16'h2828;
    PFUMX i29328 (.BLUT(n32893), .ALUT(n32894), .C0(counter_hi[3]), .Z(\csr_read_3__N_1447[2] ));
    PFUMX mux_91_i2 (.BLUT(n29836), .ALUT(\debug_branch_N_446[29] ), .C0(n30175), 
          .Z(n234[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX i29228 (.BLUT(n32403), .ALUT(n32401), .C0(n32767), .Z(n32404));
    PFUMX i29320 (.BLUT(n32881), .ALUT(n32882), .C0(counter_hi[2]), .Z(n32883));
    PFUMX mux_443_i1 (.BLUT(n822[0]), .ALUT(n948[0]), .C0(n32760), .Z(n979[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX mux_443_i2 (.BLUT(n27929), .ALUT(n948[1]), .C0(n32760), .Z(n979[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    tinyqv_mul multiplier (.accum({accum}), .\next_accum[5] (\next_accum[5] ), 
            .clk_c(clk_c), .mul_out_3__N_1510({mul_out_3__N_1510}), .\tmp_data[0] (tmp_data[0]), 
            .\tmp_data[1] (tmp_data[1]), .\tmp_data[2] (tmp_data[2]), .\tmp_data[3] (tmp_data[3]), 
            .\tmp_data[4] (tmp_data[4]), .\tmp_data[5] (tmp_data[5]), .\tmp_data[6] (tmp_data[6]), 
            .\tmp_data[7] (tmp_data[7]), .\tmp_data[8] (tmp_data[8]), .\tmp_data[9] (tmp_data[9]), 
            .\tmp_data[10] (tmp_data[10]), .\tmp_data[11] (tmp_data[11]), 
            .\tmp_data[12] (tmp_data[12]), .\tmp_data[13] (tmp_data[13]), 
            .\tmp_data[14] (tmp_data[14]), .\tmp_data[15] (tmp_data[15]), 
            .d_3__N_1868({d_3__N_1868}), .GND_net(GND_net), .VCC_net(VCC_net), 
            .\next_accum[16] (\next_accum[16] ), .\next_accum[17] (\next_accum[17] ), 
            .\next_accum[18] (\next_accum[18] ), .\next_accum[19] (\next_accum[19] ), 
            .\next_accum[6] (\next_accum[6] ), .\next_accum[7] (\next_accum[7] ), 
            .\next_accum[8] (\next_accum[8] ), .\next_accum[9] (\next_accum[9] ), 
            .\next_accum[10] (\next_accum[10] ), .\next_accum[11] (\next_accum[11] ), 
            .\next_accum[12] (\next_accum[12] ), .\next_accum[13] (\next_accum[13] ), 
            .\next_accum[14] (\next_accum[14] ), .\next_accum[15] (\next_accum[15] ), 
            .\next_accum[4] (\next_accum[4] ), .\cycle[0] (cycle[0]), .data_rs1({\data_rs1[3] , 
            data_rs1[2], data_rs1_c[1], \data_rs1[0] })) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[31:97])
    tinyqv_shifter i_shift (.\dr_3__N_1864[31] (dr_3__N_1864[31]), .\shift_amt[0] (shift_amt[0]), 
            .\shift_amt[1] (shift_amt[1]), .\dr_3__N_1864[34] (dr_3__N_1864[34]), 
            .\alu_op_in[2] (\alu_op_in[2] ), .\counter_hi[4] (counter_hi[4]), 
            .\shift_amt[4] (shift_amt_adj_3153[4]), .n34281(n34281), .\counter_hi[2] (counter_hi[2]), 
            .\shift_amt[2] (shift_amt_adj_3153[2]), .tmp_data({tmp_data}), 
            .\alu_op[3] (\alu_op[3] ), .\shift_out[0] (shift_out[0]), .\shift_out[1] (shift_out[1]), 
            .\shift_out[2] (shift_out[2]), .n32402(n32402), .n32403(n32403), 
            .n34283(n34283), .\shift_amt[3] (shift_amt_adj_3153[3])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(133[20:81])
    tinyqv_registers i_registers (.rd({rd}), .debug_reg_wen(debug_reg_wen), 
            .n32699(n32699), .n21667(n21667), .data_rs1({\data_rs1[3] , 
            data_rs1[2], data_rs1_c[1], \data_rs1[0] }), .n32733(n32733), 
            .n824(n822[0]), .debug_rd({debug_rd}), .rs1({rs1}), .rs2({rs2}), 
            .\reg_access[3][2] (\reg_access[3][2] ), .data_rs2({data_rs2}), 
            .clk_c(clk_c), .return_addr({return_addr}), .n32676(n32676), 
            .n57(n57), .\mie[13] (mie[13]), .n927(n927), .\mie[9] (mie[9]), 
            .n894(n894), .\mie[5] (mie[5]), .n861(n861), .\mie[1] (mie[1]), 
            .n794(n794), .n29683(n29683), .\mie[12] (mie[12]), .n928(n928), 
            .\mie[8] (mie[8]), .n895(n895), .\mie[4] (mie[4]), .n862(n862), 
            .n34281(n34281), .n34283(n34283), .\counter_hi[2] (counter_hi[2]), 
            .\reg_access[4][3] (\reg_access[4][3] ), .\counter_hi[3] (counter_hi[3]), 
            .n4829(n4826[1]), .n34292(n34292)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(91[9:103])
    tinyqv_counter_U0 i_instrret (.cy(cy_c), .clk_c(clk_c), .n32840(n32840), 
            .\increment_result_3__N_1925[0] (increment_result_3__N_1925[0]), 
            .instrret_count({instrret_count}), .n32665(n32665), .n32683(n32683)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(307[20] 315[6])
    \tinyqv_counter(OUTPUT_WIDTH=7)  i_cycles (.cy(cy_adj_3150), .clk_c(clk_c), 
            .n32840(n32840), .\increment_result_3__N_1911[0] (increment_result_3__N_1911[0]), 
            .cycle_count_wide({cycle_count_wide[6:4], \cycle_count_wide[3] , 
            cycle_count_wide[2:0]}), .n32701(n32701), .n32731(n32731), 
            .n32652(n32652), .n32765(n32765)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(281[40] 290[6])
    tinyqv_alu i_alu (.alu_a_in({alu_a_in}), .n32625(n32625), .n29121(n29121), 
            .alu_b_in({alu_b_in}), .\alu_op_in[2] (\alu_op_in[2] ), .n32748(n32748), 
            .n32688(n32688), .n32592(n32592), .n32646(n32646), .n32626(n32626), 
            .cy_out(cy_out), .n28225(n28225), .n31758(n31758), .n32738(n32738), 
            .n31760(n31760), .n32624(n32624), .n32749(n32749), .alu_out({alu_out}), 
            .n4901({n4901})) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(115[16:93])
    
endmodule
//
// Verilog Description of module tinyqv_mul
//

module tinyqv_mul (accum, \next_accum[5] , clk_c, mul_out_3__N_1510, 
            \tmp_data[0] , \tmp_data[1] , \tmp_data[2] , \tmp_data[3] , 
            \tmp_data[4] , \tmp_data[5] , \tmp_data[6] , \tmp_data[7] , 
            \tmp_data[8] , \tmp_data[9] , \tmp_data[10] , \tmp_data[11] , 
            \tmp_data[12] , \tmp_data[13] , \tmp_data[14] , \tmp_data[15] , 
            d_3__N_1868, GND_net, VCC_net, \next_accum[16] , \next_accum[17] , 
            \next_accum[18] , \next_accum[19] , \next_accum[6] , \next_accum[7] , 
            \next_accum[8] , \next_accum[9] , \next_accum[10] , \next_accum[11] , 
            \next_accum[12] , \next_accum[13] , \next_accum[14] , \next_accum[15] , 
            \next_accum[4] , \cycle[0] , data_rs1) /* synthesis syn_module_defined=1 */ ;
    output [15:0]accum;
    input \next_accum[5] ;
    input clk_c;
    input [3:0]mul_out_3__N_1510;
    input \tmp_data[0] ;
    input \tmp_data[1] ;
    input \tmp_data[2] ;
    input \tmp_data[3] ;
    input \tmp_data[4] ;
    input \tmp_data[5] ;
    input \tmp_data[6] ;
    input \tmp_data[7] ;
    input \tmp_data[8] ;
    input \tmp_data[9] ;
    input \tmp_data[10] ;
    input \tmp_data[11] ;
    input \tmp_data[12] ;
    input \tmp_data[13] ;
    input \tmp_data[14] ;
    input \tmp_data[15] ;
    output [19:0]d_3__N_1868;
    input GND_net;
    input VCC_net;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[4] ;
    input \cycle[0] ;
    input [3:0]data_rs1;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n7;
    wire [15:0]accum_15__N_1888;
    
    wire n29349;
    
    LUT4 accum_15__I_0_i2_3_lut (.A(accum[5]), .B(\next_accum[5] ), .C(n7), 
         .Z(accum_15__N_1888[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i2_3_lut.init = 16'hacac;
    FD1S3AX accum_i0 (.D(accum_15__N_1888[0]), .CK(clk_c), .Q(accum[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i0.GSR = "DISABLED";
    MULT18X18D a_3__I_0_11_mult_2 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(mul_out_3__N_1510[3]), 
            .A2(mul_out_3__N_1510[2]), .A1(mul_out_3__N_1510[1]), .A0(mul_out_3__N_1510[0]), 
            .B17(GND_net), .B16(GND_net), .B15(\tmp_data[15] ), .B14(\tmp_data[14] ), 
            .B13(\tmp_data[13] ), .B12(\tmp_data[12] ), .B11(\tmp_data[11] ), 
            .B10(\tmp_data[10] ), .B9(\tmp_data[9] ), .B8(\tmp_data[8] ), 
            .B7(\tmp_data[7] ), .B6(\tmp_data[6] ), .B5(\tmp_data[5] ), 
            .B4(\tmp_data[4] ), .B3(\tmp_data[3] ), .B2(\tmp_data[2] ), 
            .B1(\tmp_data[1] ), .B0(\tmp_data[0] ), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .P19(d_3__N_1868[19]), .P18(d_3__N_1868[18]), .P17(d_3__N_1868[17]), 
            .P16(d_3__N_1868[16]), .P15(d_3__N_1868[15]), .P14(d_3__N_1868[14]), 
            .P13(d_3__N_1868[13]), .P12(d_3__N_1868[12]), .P11(d_3__N_1868[11]), 
            .P10(d_3__N_1868[10]), .P9(d_3__N_1868[9]), .P8(d_3__N_1868[8]), 
            .P7(d_3__N_1868[7]), .P6(d_3__N_1868[6]), .P5(d_3__N_1868[5]), 
            .P4(d_3__N_1868[4]), .P3(d_3__N_1868[3]), .P2(d_3__N_1868[2]), 
            .P1(d_3__N_1868[1]), .P0(d_3__N_1868[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[52:83])
    defparam a_3__I_0_11_mult_2.REG_INPUTA_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTA_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTA_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_RST = "RST0";
    defparam a_3__I_0_11_mult_2.CLK0_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK1_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK2_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK3_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.HIGHSPEED_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.GSR = "DISABLED";
    defparam a_3__I_0_11_mult_2.CAS_MATCH_REG = "FALSE";
    defparam a_3__I_0_11_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam a_3__I_0_11_mult_2.MULT_BYPASS = "DISABLED";
    defparam a_3__I_0_11_mult_2.RESETMODE = "SYNC";
    FD1S3IX accum_i12 (.D(\next_accum[16] ), .CK(clk_c), .CD(n7), .Q(accum[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i12.GSR = "DISABLED";
    FD1S3AX accum_i1 (.D(accum_15__N_1888[1]), .CK(clk_c), .Q(accum[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i1.GSR = "DISABLED";
    FD1S3AX accum_i2 (.D(accum_15__N_1888[2]), .CK(clk_c), .Q(accum[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i2.GSR = "DISABLED";
    FD1S3AX accum_i3 (.D(accum_15__N_1888[3]), .CK(clk_c), .Q(accum[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i3.GSR = "DISABLED";
    FD1S3AX accum_i4 (.D(accum_15__N_1888[4]), .CK(clk_c), .Q(accum[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i4.GSR = "DISABLED";
    FD1S3AX accum_i5 (.D(accum_15__N_1888[5]), .CK(clk_c), .Q(accum[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i5.GSR = "DISABLED";
    FD1S3AX accum_i6 (.D(accum_15__N_1888[6]), .CK(clk_c), .Q(accum[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i6.GSR = "DISABLED";
    FD1S3AX accum_i7 (.D(accum_15__N_1888[7]), .CK(clk_c), .Q(accum[7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i7.GSR = "DISABLED";
    FD1S3AX accum_i8 (.D(accum_15__N_1888[8]), .CK(clk_c), .Q(accum[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i8.GSR = "DISABLED";
    FD1S3AX accum_i9 (.D(accum_15__N_1888[9]), .CK(clk_c), .Q(accum[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i9.GSR = "DISABLED";
    FD1S3AX accum_i10 (.D(accum_15__N_1888[10]), .CK(clk_c), .Q(accum[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i10.GSR = "DISABLED";
    FD1S3AX accum_i11 (.D(accum_15__N_1888[11]), .CK(clk_c), .Q(accum[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i11.GSR = "DISABLED";
    FD1S3IX accum_i13 (.D(\next_accum[17] ), .CK(clk_c), .CD(n7), .Q(accum[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i13.GSR = "DISABLED";
    FD1S3IX accum_i14 (.D(\next_accum[18] ), .CK(clk_c), .CD(n7), .Q(accum[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i14.GSR = "DISABLED";
    FD1S3IX accum_i15 (.D(\next_accum[19] ), .CK(clk_c), .CD(n7), .Q(accum[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i15.GSR = "DISABLED";
    LUT4 accum_15__I_0_i3_3_lut (.A(accum[6]), .B(\next_accum[6] ), .C(n7), 
         .Z(accum_15__N_1888[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i3_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i4_3_lut (.A(accum[7]), .B(\next_accum[7] ), .C(n7), 
         .Z(accum_15__N_1888[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i4_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i5_3_lut (.A(accum[8]), .B(\next_accum[8] ), .C(n7), 
         .Z(accum_15__N_1888[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i5_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i6_3_lut (.A(accum[9]), .B(\next_accum[9] ), .C(n7), 
         .Z(accum_15__N_1888[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i6_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i7_3_lut (.A(accum[10]), .B(\next_accum[10] ), .C(n7), 
         .Z(accum_15__N_1888[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i7_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i8_3_lut (.A(accum[11]), .B(\next_accum[11] ), .C(n7), 
         .Z(accum_15__N_1888[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i8_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i9_3_lut (.A(accum[12]), .B(\next_accum[12] ), .C(n7), 
         .Z(accum_15__N_1888[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i9_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i10_3_lut (.A(accum[13]), .B(\next_accum[13] ), .C(n7), 
         .Z(accum_15__N_1888[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i10_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i11_3_lut (.A(accum[14]), .B(\next_accum[14] ), .C(n7), 
         .Z(accum_15__N_1888[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i11_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i12_3_lut (.A(accum[15]), .B(\next_accum[15] ), .C(n7), 
         .Z(accum_15__N_1888[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i12_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i1_3_lut (.A(accum[4]), .B(\next_accum[4] ), .C(n7), 
         .Z(accum_15__N_1888[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i1_3_lut.init = 16'hacac;
    LUT4 i28476_4_lut (.A(\cycle[0] ), .B(n29349), .C(data_rs1[3]), .D(data_rs1[0]), 
         .Z(n7)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:32])
    defparam i28476_4_lut.init = 16'h5557;
    LUT4 i1_2_lut (.A(data_rs1[2]), .B(data_rs1[1]), .Z(n29349)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:32])
    defparam i1_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module tinyqv_shifter
//

module tinyqv_shifter (\dr_3__N_1864[31] , \shift_amt[0] , \shift_amt[1] , 
            \dr_3__N_1864[34] , \alu_op_in[2] , \counter_hi[4] , \shift_amt[4] , 
            n34281, \counter_hi[2] , \shift_amt[2] , tmp_data, \alu_op[3] , 
            \shift_out[0] , \shift_out[1] , \shift_out[2] , n32402, 
            n32403, n34283, \shift_amt[3] ) /* synthesis syn_module_defined=1 */ ;
    output \dr_3__N_1864[31] ;
    input \shift_amt[0] ;
    input \shift_amt[1] ;
    output \dr_3__N_1864[34] ;
    input \alu_op_in[2] ;
    input \counter_hi[4] ;
    input \shift_amt[4] ;
    input n34281;
    input \counter_hi[2] ;
    input \shift_amt[2] ;
    input [31:0]tmp_data;
    input \alu_op[3] ;
    output \shift_out[0] ;
    output \shift_out[1] ;
    output \shift_out[2] ;
    input n32402;
    output n32403;
    input n34283;
    input \shift_amt[3] ;
    
    
    wire n30403, n30404, n30921, n30408, n109, n113, n30413, n30342, 
        n30343;
    wire [5:0]shift_amt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[16:25])
    wire [31:0]a_for_shift_right;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[17:34])
    
    wire n41, n30357, n30358;
    wire [65:0]dr_3__N_1864;
    
    wire n46, n48, n30400, n30409, n30410, n42, n44, n30399, 
        n30416, n30417, n38, n40, n30398, n33, n117, n121, n30414, 
        n35, n34, n36, n30397, n37, n125, n129, n30415, n9550, 
        n9548, n8985, n39, n105, n101, n30338, n30339, n30340, 
        n30341, n30353, n30354, n30355, n30356, n30405, n30406, 
        n30407, n30412, n30330, n30331, n30332, n30333, n61, n63, 
        n30352, n30334, n30335, n57, n59, n30351, n4, n32813, 
        n30923, n30922, n32814, n62, n53, n55, n30350, n49, 
        n51, n30349, n30336, n30337, n45, n47, n30348, n43, 
        n30347, n30346, n30345, n50, n52, n60, n54, n56, n32, 
        n58, n30539, n30402, n30401;
    
    PFUMX i27699 (.BLUT(n30403), .ALUT(n30404), .C0(n30921), .Z(n30408));
    PFUMX i27704 (.BLUT(n109), .ALUT(n113), .C0(n30921), .Z(n30413));
    L6MUX21 i27635 (.D0(n30342), .D1(n30343), .SD(shift_amt[4]), .Z(\dr_3__N_1864[31] ));
    LUT4 top_bit_I_0_i41_3_lut (.A(a_for_shift_right[9]), .B(a_for_shift_right[10]), 
         .C(\shift_amt[0] ), .Z(n41)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i41_3_lut.init = 16'hcaca;
    L6MUX21 i27650 (.D0(n30357), .D1(n30358), .SD(shift_amt[4]), .Z(dr_3__N_1864[32]));
    LUT4 i27691_3_lut (.A(n46), .B(n48), .C(\shift_amt[1] ), .Z(n30400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27691_3_lut.init = 16'hcaca;
    L6MUX21 i27702 (.D0(n30409), .D1(n30410), .SD(shift_amt[4]), .Z(dr_3__N_1864[33]));
    LUT4 i27690_3_lut (.A(n42), .B(n44), .C(\shift_amt[1] ), .Z(n30399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27690_3_lut.init = 16'hcaca;
    L6MUX21 i27709 (.D0(n30416), .D1(n30417), .SD(shift_amt[4]), .Z(\dr_3__N_1864[34] ));
    LUT4 i27689_3_lut (.A(n38), .B(n40), .C(\shift_amt[1] ), .Z(n30398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27689_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i33_3_lut (.A(a_for_shift_right[1]), .B(a_for_shift_right[2]), 
         .C(\shift_amt[0] ), .Z(n33)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i33_3_lut.init = 16'hcaca;
    PFUMX i27705 (.BLUT(n117), .ALUT(n121), .C0(n30921), .Z(n30414));
    LUT4 top_bit_I_0_i35_3_lut (.A(a_for_shift_right[3]), .B(a_for_shift_right[4]), 
         .C(\shift_amt[0] ), .Z(n35)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i35_3_lut.init = 16'hcaca;
    LUT4 i27688_3_lut (.A(n34), .B(n36), .C(\shift_amt[1] ), .Z(n30397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27688_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i37_3_lut (.A(a_for_shift_right[5]), .B(a_for_shift_right[6]), 
         .C(\shift_amt[0] ), .Z(n37)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i37_3_lut.init = 16'hcaca;
    PFUMX i27706 (.BLUT(n125), .ALUT(n129), .C0(n30921), .Z(n30415));
    LUT4 i6868_3_lut (.A(dr_3__N_1864[32]), .B(dr_3__N_1864[33]), .C(\alu_op_in[2] ), 
         .Z(n9550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i6868_3_lut.init = 16'hcaca;
    LUT4 i6866_3_lut (.A(dr_3__N_1864[33]), .B(dr_3__N_1864[32]), .C(\alu_op_in[2] ), 
         .Z(n9548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i6866_3_lut.init = 16'hcaca;
    LUT4 i6307_3_lut (.A(\dr_3__N_1864[34] ), .B(\dr_3__N_1864[31] ), .C(\alu_op_in[2] ), 
         .Z(n8985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i6307_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i105_3_lut (.A(n39), .B(n41), .C(\shift_amt[1] ), 
         .Z(n105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i105_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i101_3_lut (.A(n35), .B(n37), .C(\shift_amt[1] ), 
         .Z(n101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i101_3_lut.init = 16'hcaca;
    L6MUX21 i27633 (.D0(n30338), .D1(n30339), .SD(shift_amt[3]), .Z(n30342));
    L6MUX21 i27634 (.D0(n30340), .D1(n30341), .SD(shift_amt[3]), .Z(n30343));
    L6MUX21 i27648 (.D0(n30353), .D1(n30354), .SD(shift_amt[3]), .Z(n30357));
    L6MUX21 i27649 (.D0(n30355), .D1(n30356), .SD(shift_amt[3]), .Z(n30358));
    L6MUX21 i27700 (.D0(n30405), .D1(n30406), .SD(shift_amt[3]), .Z(n30409));
    L6MUX21 i27701 (.D0(n30407), .D1(n30408), .SD(shift_amt[3]), .Z(n30410));
    L6MUX21 i27707 (.D0(n30412), .D1(n30413), .SD(shift_amt[3]), .Z(n30416));
    L6MUX21 i27708 (.D0(n30414), .D1(n30415), .SD(shift_amt[3]), .Z(n30417));
    PFUMX i27629 (.BLUT(n30330), .ALUT(n30331), .C0(shift_amt[2]), .Z(n30338));
    PFUMX i27630 (.BLUT(n30332), .ALUT(n30333), .C0(shift_amt[2]), .Z(n30339));
    LUT4 i27643_3_lut (.A(n61), .B(n63), .C(\shift_amt[1] ), .Z(n30352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27643_3_lut.init = 16'hcaca;
    PFUMX i27631 (.BLUT(n30334), .ALUT(n30335), .C0(shift_amt[2]), .Z(n30340));
    LUT4 i27642_3_lut (.A(n57), .B(n59), .C(\shift_amt[1] ), .Z(n30351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27642_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(\counter_hi[4] ), .B(\alu_op_in[2] ), .C(n4), 
         .D(\shift_amt[4] ), .Z(shift_amt[4])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i2_3_lut_4_lut.init = 16'h9669;
    LUT4 i4696_3_lut_4_lut (.A(n34281), .B(\alu_op_in[2] ), .C(n4), .D(\shift_amt[4] ), 
         .Z(shift_amt[5])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4696_3_lut_4_lut.init = 16'hf990;
    LUT4 i28235_2_lut_rep_798 (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .Z(n32813)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i28235_2_lut_rep_798.init = 16'h6666;
    LUT4 i4676_rep_135_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .C(\shift_amt[2] ), .Z(n30921)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4676_rep_135_2_lut_3_lut.init = 16'h6969;
    LUT4 i4676_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), .C(\shift_amt[2] ), 
         .Z(shift_amt[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4676_2_lut_3_lut.init = 16'h6969;
    LUT4 i4676_rep_137_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .C(\shift_amt[2] ), .Z(n30923)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4676_rep_137_2_lut_3_lut.init = 16'h6969;
    LUT4 i4676_rep_136_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .C(\shift_amt[2] ), .Z(n30922)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4676_rep_136_2_lut_3_lut.init = 16'h6969;
    LUT4 i15262_2_lut_rep_799 (.A(tmp_data[31]), .B(\alu_op[3] ), .Z(n32814)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i15262_2_lut_rep_799.init = 16'h8888;
    LUT4 i6308_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n8985), .Z(\shift_out[0] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i6308_3_lut_4_lut.init = 16'h8f80;
    LUT4 i6867_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n9548), .Z(\shift_out[1] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i6867_3_lut_4_lut.init = 16'h8f80;
    LUT4 i27695_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(\shift_amt[1] ), 
         .D(n62), .Z(n30404)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i27695_3_lut_4_lut.init = 16'h8f80;
    LUT4 i6869_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n9550), .Z(\shift_out[2] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i6869_3_lut_4_lut.init = 16'h8f80;
    LUT4 n32402_bdd_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n32402), .Z(n32403)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam n32402_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 top_bit_I_0_i63_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), 
         .C(\shift_amt[0] ), .D(a_for_shift_right[31]), .Z(n63)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam top_bit_I_0_i63_3_lut_4_lut.init = 16'h8f80;
    LUT4 i27641_3_lut (.A(n53), .B(n55), .C(\shift_amt[1] ), .Z(n30350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27641_3_lut.init = 16'hcaca;
    LUT4 i27640_3_lut (.A(n49), .B(n51), .C(\shift_amt[1] ), .Z(n30349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27640_3_lut.init = 16'hcaca;
    PFUMX i27632 (.BLUT(n30336), .ALUT(n30337), .C0(shift_amt[2]), .Z(n30341));
    LUT4 top_bit_I_0_i39_3_lut (.A(a_for_shift_right[7]), .B(a_for_shift_right[8]), 
         .C(\shift_amt[0] ), .Z(n39)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i39_3_lut.init = 16'hcaca;
    LUT4 i27639_3_lut (.A(n45), .B(n47), .C(\shift_amt[1] ), .Z(n30348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27639_3_lut.init = 16'hcaca;
    LUT4 i27638_3_lut (.A(n41), .B(n43), .C(\shift_amt[1] ), .Z(n30347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27638_3_lut.init = 16'hcaca;
    LUT4 i27637_3_lut (.A(n37), .B(n39), .C(\shift_amt[1] ), .Z(n30346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27637_3_lut.init = 16'hcaca;
    LUT4 i27636_3_lut (.A(n33), .B(n35), .C(\shift_amt[1] ), .Z(n30345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27636_3_lut.init = 16'hcaca;
    PFUMX i27644 (.BLUT(n30345), .ALUT(n30346), .C0(n30923), .Z(n30353));
    LUT4 top_bit_I_0_i50_3_lut (.A(a_for_shift_right[18]), .B(a_for_shift_right[19]), 
         .C(\shift_amt[0] ), .Z(n50)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i50_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i52_3_lut (.A(a_for_shift_right[20]), .B(a_for_shift_right[21]), 
         .C(\shift_amt[0] ), .Z(n52)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i52_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i21_3_lut (.A(tmp_data[11]), .B(tmp_data[20]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i22_3_lut (.A(tmp_data[10]), .B(tmp_data[21]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i19_3_lut (.A(tmp_data[13]), .B(tmp_data[18]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i20_3_lut (.A(tmp_data[12]), .B(tmp_data[19]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 i27628_3_lut (.A(n60), .B(n62), .C(\shift_amt[1] ), .Z(n30337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27628_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i54_3_lut (.A(a_for_shift_right[22]), .B(a_for_shift_right[23]), 
         .C(\shift_amt[0] ), .Z(n54)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i54_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i56_3_lut (.A(a_for_shift_right[24]), .B(a_for_shift_right[25]), 
         .C(\shift_amt[0] ), .Z(n56)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i56_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i25_3_lut (.A(tmp_data[7]), .B(tmp_data[24]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i26_3_lut (.A(tmp_data[6]), .B(tmp_data[25]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i23_3_lut (.A(tmp_data[9]), .B(tmp_data[22]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i24_3_lut (.A(tmp_data[8]), .B(tmp_data[23]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i32_3_lut (.A(a_for_shift_right[0]), .B(a_for_shift_right[1]), 
         .C(\shift_amt[0] ), .Z(n32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i32_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i1_3_lut (.A(tmp_data[31]), .B(tmp_data[0]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i34_3_lut (.A(a_for_shift_right[2]), .B(a_for_shift_right[3]), 
         .C(\shift_amt[0] ), .Z(n34)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i34_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i3_3_lut (.A(tmp_data[29]), .B(tmp_data[2]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i4_3_lut (.A(tmp_data[28]), .B(tmp_data[3]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i2_3_lut (.A(tmp_data[30]), .B(tmp_data[1]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i36_3_lut (.A(a_for_shift_right[4]), .B(a_for_shift_right[5]), 
         .C(\shift_amt[0] ), .Z(n36)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i36_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i38_3_lut (.A(a_for_shift_right[6]), .B(a_for_shift_right[7]), 
         .C(\shift_amt[0] ), .Z(n38)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i38_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i7_3_lut (.A(tmp_data[25]), .B(tmp_data[6]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i8_3_lut (.A(tmp_data[24]), .B(tmp_data[7]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i5_3_lut (.A(tmp_data[27]), .B(tmp_data[4]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i6_3_lut (.A(tmp_data[26]), .B(tmp_data[5]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i40_3_lut (.A(a_for_shift_right[8]), .B(a_for_shift_right[9]), 
         .C(\shift_amt[0] ), .Z(n40)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i40_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i42_3_lut (.A(a_for_shift_right[10]), .B(a_for_shift_right[11]), 
         .C(\shift_amt[0] ), .Z(n42)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i42_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i9_3_lut (.A(tmp_data[23]), .B(tmp_data[8]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i10_3_lut (.A(tmp_data[22]), .B(tmp_data[9]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i11_3_lut (.A(tmp_data[21]), .B(tmp_data[10]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i44_3_lut (.A(a_for_shift_right[12]), .B(a_for_shift_right[13]), 
         .C(\shift_amt[0] ), .Z(n44)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i44_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i46_3_lut (.A(a_for_shift_right[14]), .B(a_for_shift_right[15]), 
         .C(\shift_amt[0] ), .Z(n46)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i46_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i16_3_lut (.A(tmp_data[16]), .B(tmp_data[15]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i16_3_lut.init = 16'hcaca;
    PFUMX i27645 (.BLUT(n30347), .ALUT(n30348), .C0(n30923), .Z(n30354));
    LUT4 top_bit_I_0_i58_3_lut (.A(a_for_shift_right[26]), .B(a_for_shift_right[27]), 
         .C(\shift_amt[0] ), .Z(n58)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i58_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i60_3_lut (.A(a_for_shift_right[28]), .B(a_for_shift_right[29]), 
         .C(\shift_amt[0] ), .Z(n60)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i60_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i29_3_lut (.A(tmp_data[3]), .B(tmp_data[28]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i30_3_lut (.A(tmp_data[2]), .B(tmp_data[29]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i27_3_lut (.A(tmp_data[5]), .B(tmp_data[26]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i28_3_lut (.A(tmp_data[4]), .B(tmp_data[27]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i62_3_lut (.A(a_for_shift_right[30]), .B(a_for_shift_right[31]), 
         .C(\shift_amt[0] ), .Z(n62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i62_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i31_3_lut (.A(tmp_data[1]), .B(tmp_data[30]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i32_3_lut (.A(tmp_data[0]), .B(tmp_data[31]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i43_3_lut (.A(a_for_shift_right[11]), .B(a_for_shift_right[12]), 
         .C(\shift_amt[0] ), .Z(n43)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i43_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i45_3_lut (.A(a_for_shift_right[13]), .B(a_for_shift_right[14]), 
         .C(\shift_amt[0] ), .Z(n45)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i45_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i14_3_lut (.A(tmp_data[18]), .B(tmp_data[13]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i15_3_lut (.A(tmp_data[17]), .B(tmp_data[14]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i12_3_lut (.A(tmp_data[20]), .B(tmp_data[11]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i13_3_lut (.A(tmp_data[19]), .B(tmp_data[12]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i47_4_lut (.A(tmp_data[16]), .B(tmp_data[15]), .C(\alu_op_in[2] ), 
         .D(\shift_amt[0] ), .Z(n47)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A !((C (D)+!C !(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i47_4_lut.init = 16'hacca;
    LUT4 top_bit_I_0_i49_3_lut (.A(a_for_shift_right[17]), .B(a_for_shift_right[18]), 
         .C(\shift_amt[0] ), .Z(n49)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i49_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i18_3_lut (.A(tmp_data[14]), .B(tmp_data[17]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 i28237_2_lut (.A(n34283), .B(\alu_op_in[2] ), .Z(n30539)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i28237_2_lut.init = 16'h6666;
    LUT4 top_bit_I_0_i48_3_lut (.A(a_for_shift_right[16]), .B(a_for_shift_right[17]), 
         .C(\shift_amt[0] ), .Z(n48)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i48_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i17_3_lut (.A(tmp_data[15]), .B(tmp_data[16]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i17_3_lut.init = 16'hcaca;
    PFUMX i27646 (.BLUT(n30349), .ALUT(n30350), .C0(n30922), .Z(n30355));
    LUT4 i27627_3_lut (.A(n56), .B(n58), .C(\shift_amt[1] ), .Z(n30336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27627_3_lut.init = 16'hcaca;
    LUT4 i27626_3_lut (.A(n52), .B(n54), .C(\shift_amt[1] ), .Z(n30335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27626_3_lut.init = 16'hcaca;
    PFUMX i27647 (.BLUT(n30351), .ALUT(n30352), .C0(n30922), .Z(n30356));
    LUT4 top_bit_I_0_i51_3_lut (.A(a_for_shift_right[19]), .B(a_for_shift_right[20]), 
         .C(\shift_amt[0] ), .Z(n51)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i51_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i53_3_lut (.A(a_for_shift_right[21]), .B(a_for_shift_right[22]), 
         .C(\shift_amt[0] ), .Z(n53)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i53_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i55_3_lut (.A(a_for_shift_right[23]), .B(a_for_shift_right[24]), 
         .C(\shift_amt[0] ), .Z(n55)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i55_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i57_3_lut (.A(a_for_shift_right[25]), .B(a_for_shift_right[26]), 
         .C(\shift_amt[0] ), .Z(n57)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i57_3_lut.init = 16'hcaca;
    LUT4 i27625_3_lut (.A(n48), .B(n50), .C(\shift_amt[1] ), .Z(n30334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27625_3_lut.init = 16'hcaca;
    LUT4 i27624_3_lut (.A(n44), .B(n46), .C(\shift_amt[1] ), .Z(n30333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27624_3_lut.init = 16'hcaca;
    LUT4 i27623_3_lut (.A(n40), .B(n42), .C(\shift_amt[1] ), .Z(n30332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27623_3_lut.init = 16'hcaca;
    LUT4 i27622_3_lut (.A(n36), .B(n38), .C(\shift_amt[1] ), .Z(n30331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27622_3_lut.init = 16'hcaca;
    LUT4 i27621_3_lut (.A(n32), .B(n34), .C(\shift_amt[1] ), .Z(n30330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27621_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i59_3_lut (.A(a_for_shift_right[27]), .B(a_for_shift_right[28]), 
         .C(\shift_amt[0] ), .Z(n59)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i59_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i61_3_lut (.A(a_for_shift_right[29]), .B(a_for_shift_right[30]), 
         .C(\shift_amt[0] ), .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i61_3_lut.init = 16'hcaca;
    PFUMX i27703 (.BLUT(n101), .ALUT(n105), .C0(n30923), .Z(n30412));
    LUT4 i6334_4_lut (.A(a_for_shift_right[31]), .B(n32814), .C(\shift_amt[0] ), 
         .D(\shift_amt[1] ), .Z(n129)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam i6334_4_lut.init = 16'hccca;
    LUT4 top_bit_I_0_i125_3_lut (.A(n59), .B(n61), .C(\shift_amt[1] ), 
         .Z(n125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i125_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i121_3_lut (.A(n55), .B(n57), .C(\shift_amt[1] ), 
         .Z(n121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i121_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i117_3_lut (.A(n51), .B(n53), .C(\shift_amt[1] ), 
         .Z(n117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i117_3_lut.init = 16'hcaca;
    PFUMX i27696 (.BLUT(n30397), .ALUT(n30398), .C0(n30923), .Z(n30405));
    LUT4 top_bit_I_0_i113_3_lut (.A(n47), .B(n49), .C(\shift_amt[1] ), 
         .Z(n113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i113_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i109_3_lut (.A(n43), .B(n45), .C(\shift_amt[1] ), 
         .Z(n109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i109_3_lut.init = 16'hcaca;
    LUT4 i27694_3_lut (.A(n58), .B(n60), .C(\shift_amt[1] ), .Z(n30403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27694_3_lut.init = 16'hcaca;
    LUT4 i27693_3_lut (.A(n54), .B(n56), .C(\shift_amt[1] ), .Z(n30402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27693_3_lut.init = 16'hcaca;
    LUT4 i4689_3_lut_4_lut (.A(\shift_amt[2] ), .B(n32813), .C(n30539), 
         .D(\shift_amt[3] ), .Z(n4)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[28:55])
    defparam i4689_3_lut_4_lut.init = 16'h2f02;
    LUT4 i2_3_lut_4_lut_adj_299 (.A(\shift_amt[2] ), .B(n32813), .C(n30539), 
         .D(\shift_amt[3] ), .Z(shift_amt[3])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[28:55])
    defparam i2_3_lut_4_lut_adj_299.init = 16'hd22d;
    PFUMX i27697 (.BLUT(n30399), .ALUT(n30400), .C0(n30922), .Z(n30406));
    LUT4 i27692_3_lut (.A(n50), .B(n52), .C(\shift_amt[1] ), .Z(n30401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27692_3_lut.init = 16'hcaca;
    PFUMX i27698 (.BLUT(n30401), .ALUT(n30402), .C0(n30922), .Z(n30407));
    
endmodule
//
// Verilog Description of module tinyqv_registers
//

module tinyqv_registers (rd, debug_reg_wen, n32699, n21667, data_rs1, 
            n32733, n824, debug_rd, rs1, rs2, \reg_access[3][2] , 
            data_rs2, clk_c, return_addr, n32676, n57, \mie[13] , 
            n927, \mie[9] , n894, \mie[5] , n861, \mie[1] , n794, 
            n29683, \mie[12] , n928, \mie[8] , n895, \mie[4] , n862, 
            n34281, n34283, \counter_hi[2] , \reg_access[4][3] , \counter_hi[3] , 
            n4829, n34292) /* synthesis syn_module_defined=1 */ ;
    input [3:0]rd;
    input debug_reg_wen;
    input n32699;
    input n21667;
    output [3:0]data_rs1;
    input n32733;
    output n824;
    input [3:0]debug_rd;
    input [3:0]rs1;
    input [3:0]rs2;
    output \reg_access[3][2] ;
    output [3:0]data_rs2;
    input clk_c;
    output [23:1]return_addr;
    input n32676;
    input n57;
    input \mie[13] ;
    output n927;
    input \mie[9] ;
    output n894;
    input \mie[5] ;
    output n861;
    input \mie[1] ;
    output n794;
    input n29683;
    input \mie[12] ;
    output n928;
    input \mie[8] ;
    output n895;
    input \mie[4] ;
    output n862;
    input n34281;
    input n34283;
    input \counter_hi[2] ;
    output \reg_access[4][3] ;
    input \counter_hi[3] ;
    output n4829;
    output n34292;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n32556, n32555, n32554, n32553, n32779;
    wire [31:0]\registers[15] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_15__3__N_1825, registers_15__2__N_1828, registers_15__1__N_1829, 
        registers_15__0__N_1830;
    wire [31:0]\registers[14] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_14__3__N_1819, registers_14__2__N_1822, registers_14__1__N_1823, 
        registers_14__0__N_1824;
    wire [31:0]\registers[13] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_13__3__N_1813, registers_13__2__N_1816, registers_13__1__N_1817, 
        registers_13__0__N_1818;
    wire [31:0]\registers[12] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_12__3__N_1807, registers_12__2__N_1810, registers_12__1__N_1811, 
        registers_12__0__N_1812, n32780;
    wire [31:0]\registers[11] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_11__3__N_1801, registers_11__2__N_1804, registers_11__1__N_1805, 
        registers_11__0__N_1806;
    wire [31:0]\registers[10] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_10__3__N_1795, registers_10__2__N_1798, registers_10__1__N_1799, 
        registers_10__0__N_1800;
    wire [31:0]\registers[9] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_9__3__N_1789, registers_9__2__N_1792, registers_9__1__N_1793, 
        registers_9__0__N_1794;
    wire [31:0]\registers[8] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_8__3__N_1783, registers_8__2__N_1786, registers_8__1__N_1787, 
        registers_8__0__N_1788, n32781;
    wire [31:0]\registers[7] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_7__3__N_1777, registers_7__2__N_1780, registers_7__1__N_1781, 
        registers_7__0__N_1782;
    wire [31:0]\registers[6] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_6__3__N_1771, registers_6__2__N_1774, registers_6__1__N_1775, 
        registers_6__0__N_1776;
    wire [31:0]\registers[5] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_5__0__N_1770, registers_5__2__N_1768, registers_5__3__N_1765, 
        registers_5__1__N_1769, n32786;
    wire [31:0]\registers[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_2__3__N_1759, registers_2__2__N_1762, registers_2__1__N_1763, 
        registers_2__0__N_1764;
    wire [31:0]\registers[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_1__2__N_1756, registers_1__1__N_1757, registers_1__0__N_1758, 
        n12, n11, registers_1__3__N_1753, n9, n8, n5, n12_adj_3130, 
        n11_adj_3131, n9_adj_3132, n8_adj_3133, n5_adj_3134, n30426, 
        n12_adj_3135, n30383, n11_adj_3136, n9_adj_3137, n8_adj_3138, 
        n12_adj_3139, n11_adj_3140, n9_adj_3141, n8_adj_3142, n30389, 
        n30298, n30299, n30388, n30387, n30382, n30386, n30385, 
        n30384, n30374, n30373, n30372, n30379, n30380, n30394, 
        n30395, n30371, n30370, n30369, n30294, n30295, n30309, 
        n30310, n30313, n30375, n30376, n30390, n30391, n30427, 
        n30430, n30433, n30434, n30437, n30286, n30287, n30301, 
        n30302, n30368, n30367, n30308, n30307, n30306, n30305, 
        n30447, n30440, n30304, n30303, n30314, n30293, n30292, 
        n30291, n30290, n30289, n30288, n30296, n30297, n30311, 
        n30312, n30377, n30378, n30392, n30393, n30428, n30429, 
        n30431, n30435, n30436, n30438, n30441, n30444, n30442, 
        n30443, n30445, n30448, n30451, n30449, n30450, n30452, 
        n5_adj_3143, n4, n5_adj_3144, n4_adj_3145;
    
    LUT4 i1_2_lut_rep_541_3_lut (.A(rd[0]), .B(debug_reg_wen), .C(rd[1]), 
         .Z(n32556)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_541_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_540_3_lut (.A(rd[0]), .B(rd[1]), .C(debug_reg_wen), 
         .Z(n32555)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_rep_540_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_539_3_lut (.A(rd[0]), .B(rd[1]), .C(debug_reg_wen), 
         .Z(n32554)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_539_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_538_3_lut (.A(rd[0]), .B(debug_reg_wen), .C(rd[1]), 
         .Z(n32553)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_rep_538_3_lut.init = 16'h0404;
    LUT4 i1_4_lut (.A(n32699), .B(n21667), .C(data_rs1[0]), .D(n32733), 
         .Z(n824)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam i1_4_lut.init = 16'h5044;
    LUT4 registers_15__7__I_0_3_lut_4_lut (.A(n32779), .B(n32554), .C(debug_rd[3]), 
         .D(\registers[15] [7]), .Z(registers_15__3__N_1825)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_15__6__I_0_3_lut_4_lut (.A(n32779), .B(n32554), .C(debug_rd[2]), 
         .D(\registers[15] [6]), .Z(registers_15__2__N_1828)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_15__5__I_0_3_lut_4_lut (.A(n32779), .B(n32554), .C(debug_rd[1]), 
         .D(\registers[15] [5]), .Z(registers_15__1__N_1829)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_15__4__I_0_3_lut_4_lut (.A(n32779), .B(n32554), .C(debug_rd[0]), 
         .D(\registers[15] [4]), .Z(registers_15__0__N_1830)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__7__I_0_3_lut_4_lut (.A(n32779), .B(n32555), .C(debug_rd[3]), 
         .D(\registers[14] [7]), .Z(registers_14__3__N_1819)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__6__I_0_3_lut_4_lut (.A(n32779), .B(n32555), .C(debug_rd[2]), 
         .D(\registers[14] [6]), .Z(registers_14__2__N_1822)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__5__I_0_3_lut_4_lut (.A(n32779), .B(n32555), .C(debug_rd[1]), 
         .D(\registers[14] [5]), .Z(registers_14__1__N_1823)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__4__I_0_3_lut_4_lut (.A(n32779), .B(n32555), .C(debug_rd[0]), 
         .D(\registers[14] [4]), .Z(registers_14__0__N_1824)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__7__I_0_3_lut_4_lut (.A(n32779), .B(n32556), .C(debug_rd[3]), 
         .D(\registers[13] [7]), .Z(registers_13__3__N_1813)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__6__I_0_3_lut_4_lut (.A(n32779), .B(n32556), .C(debug_rd[2]), 
         .D(\registers[13] [6]), .Z(registers_13__2__N_1816)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__5__I_0_3_lut_4_lut (.A(n32779), .B(n32556), .C(debug_rd[1]), 
         .D(\registers[13] [5]), .Z(registers_13__1__N_1817)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__4__I_0_3_lut_4_lut (.A(n32779), .B(n32556), .C(debug_rd[0]), 
         .D(\registers[13] [4]), .Z(registers_13__0__N_1818)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__7__I_0_3_lut_4_lut (.A(n32779), .B(n32553), .C(debug_rd[3]), 
         .D(\registers[12] [7]), .Z(registers_12__3__N_1807)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__6__I_0_3_lut_4_lut (.A(n32779), .B(n32553), .C(debug_rd[2]), 
         .D(\registers[12] [6]), .Z(registers_12__2__N_1810)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__5__I_0_3_lut_4_lut (.A(n32779), .B(n32553), .C(debug_rd[1]), 
         .D(\registers[12] [5]), .Z(registers_12__1__N_1811)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__4__I_0_3_lut_4_lut (.A(n32779), .B(n32553), .C(debug_rd[0]), 
         .D(\registers[12] [4]), .Z(registers_12__0__N_1812)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_11__7__I_0_3_lut_4_lut (.A(n32780), .B(n32554), .C(debug_rd[3]), 
         .D(\registers[11] [7]), .Z(registers_11__3__N_1801)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__6__I_0_3_lut_4_lut (.A(n32780), .B(n32554), .C(debug_rd[2]), 
         .D(\registers[11] [6]), .Z(registers_11__2__N_1804)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__5__I_0_3_lut_4_lut (.A(n32780), .B(n32554), .C(debug_rd[1]), 
         .D(\registers[11] [5]), .Z(registers_11__1__N_1805)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__4__I_0_3_lut_4_lut (.A(n32780), .B(n32554), .C(debug_rd[0]), 
         .D(\registers[11] [4]), .Z(registers_11__0__N_1806)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__7__I_0_3_lut_4_lut (.A(n32780), .B(n32555), .C(debug_rd[3]), 
         .D(\registers[10] [7]), .Z(registers_10__3__N_1795)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__6__I_0_3_lut_4_lut (.A(n32780), .B(n32555), .C(debug_rd[2]), 
         .D(\registers[10] [6]), .Z(registers_10__2__N_1798)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__5__I_0_3_lut_4_lut (.A(n32780), .B(n32555), .C(debug_rd[1]), 
         .D(\registers[10] [5]), .Z(registers_10__1__N_1799)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__4__I_0_3_lut_4_lut (.A(n32780), .B(n32555), .C(debug_rd[0]), 
         .D(\registers[10] [4]), .Z(registers_10__0__N_1800)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__7__I_0_3_lut_4_lut (.A(n32780), .B(n32556), .C(debug_rd[3]), 
         .D(\registers[9] [7]), .Z(registers_9__3__N_1789)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__6__I_0_3_lut_4_lut (.A(n32780), .B(n32556), .C(debug_rd[2]), 
         .D(\registers[9] [6]), .Z(registers_9__2__N_1792)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__5__I_0_3_lut_4_lut (.A(n32780), .B(n32556), .C(debug_rd[1]), 
         .D(\registers[9] [5]), .Z(registers_9__1__N_1793)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__4__I_0_3_lut_4_lut (.A(n32780), .B(n32556), .C(debug_rd[0]), 
         .D(\registers[9] [4]), .Z(registers_9__0__N_1794)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__7__I_0_3_lut_4_lut (.A(n32780), .B(n32553), .C(debug_rd[3]), 
         .D(\registers[8] [7]), .Z(registers_8__3__N_1783)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__6__I_0_3_lut_4_lut (.A(n32780), .B(n32553), .C(debug_rd[2]), 
         .D(\registers[8] [6]), .Z(registers_8__2__N_1786)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__5__I_0_3_lut_4_lut (.A(n32780), .B(n32553), .C(debug_rd[1]), 
         .D(\registers[8] [5]), .Z(registers_8__1__N_1787)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__4__I_0_3_lut_4_lut (.A(n32780), .B(n32553), .C(debug_rd[0]), 
         .D(\registers[8] [4]), .Z(registers_8__0__N_1788)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__7__I_0_3_lut_4_lut (.A(n32781), .B(n32554), .C(debug_rd[3]), 
         .D(\registers[7] [7]), .Z(registers_7__3__N_1777)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__6__I_0_3_lut_4_lut (.A(n32781), .B(n32554), .C(debug_rd[2]), 
         .D(\registers[7] [6]), .Z(registers_7__2__N_1780)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__5__I_0_3_lut_4_lut (.A(n32781), .B(n32554), .C(debug_rd[1]), 
         .D(\registers[7] [5]), .Z(registers_7__1__N_1781)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__4__I_0_3_lut_4_lut (.A(n32781), .B(n32554), .C(debug_rd[0]), 
         .D(\registers[7] [4]), .Z(registers_7__0__N_1782)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__7__I_0_3_lut_4_lut (.A(n32781), .B(n32555), .C(debug_rd[3]), 
         .D(\registers[6] [7]), .Z(registers_6__3__N_1771)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__6__I_0_3_lut_4_lut (.A(n32781), .B(n32555), .C(debug_rd[2]), 
         .D(\registers[6] [6]), .Z(registers_6__2__N_1774)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__5__I_0_3_lut_4_lut (.A(n32781), .B(n32555), .C(debug_rd[1]), 
         .D(\registers[6] [5]), .Z(registers_6__1__N_1775)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__4__I_0_3_lut_4_lut (.A(n32781), .B(n32555), .C(debug_rd[0]), 
         .D(\registers[6] [4]), .Z(registers_6__0__N_1776)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__4__I_0_3_lut_4_lut (.A(n32781), .B(n32556), .C(debug_rd[0]), 
         .D(\registers[5] [4]), .Z(registers_5__0__N_1770)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__6__I_0_3_lut_4_lut (.A(n32781), .B(n32556), .C(debug_rd[2]), 
         .D(\registers[5] [6]), .Z(registers_5__2__N_1768)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__7__I_0_3_lut_4_lut (.A(n32781), .B(n32556), .C(debug_rd[3]), 
         .D(\registers[5] [7]), .Z(registers_5__3__N_1765)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__5__I_0_3_lut_4_lut (.A(n32781), .B(n32556), .C(debug_rd[1]), 
         .D(\registers[5] [5]), .Z(registers_5__1__N_1769)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_2__7__I_0_3_lut_4_lut (.A(n32555), .B(n32786), .C(debug_rd[3]), 
         .D(\registers[2] [7]), .Z(registers_2__3__N_1759)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__7__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__6__I_0_3_lut_4_lut (.A(n32555), .B(n32786), .C(debug_rd[2]), 
         .D(\registers[2] [6]), .Z(registers_2__2__N_1762)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__5__I_0_3_lut_4_lut (.A(n32555), .B(n32786), .C(debug_rd[1]), 
         .D(\registers[2] [5]), .Z(registers_2__1__N_1763)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__4__I_0_3_lut_4_lut (.A(n32555), .B(n32786), .C(debug_rd[0]), 
         .D(\registers[2] [4]), .Z(registers_2__0__N_1764)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__4__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__6__I_0_3_lut_4_lut (.A(n32556), .B(n32786), .C(debug_rd[2]), 
         .D(\registers[1] [6]), .Z(registers_1__2__N_1756)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__5__I_0_3_lut_4_lut (.A(n32556), .B(n32786), .C(debug_rd[1]), 
         .D(\registers[1] [5]), .Z(registers_1__1__N_1757)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__4__I_0_3_lut_4_lut (.A(n32556), .B(n32786), .C(debug_rd[0]), 
         .D(\registers[1] [4]), .Z(registers_1__0__N_1758)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__4__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 rs1_3__I_0_Mux_1_i12_3_lut (.A(\registers[14] [5]), .B(\registers[15] [5]), 
         .C(rs1[0]), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i12_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i11_3_lut (.A(\registers[12] [5]), .B(\registers[13] [5]), 
         .C(rs1[0]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i11_3_lut.init = 16'hcaca;
    LUT4 registers_1__7__I_0_3_lut_4_lut (.A(n32556), .B(n32786), .C(debug_rd[3]), 
         .D(\registers[1] [7]), .Z(registers_1__3__N_1753)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__7__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 rs1_3__I_0_Mux_1_i9_3_lut (.A(\registers[10] [5]), .B(\registers[11] [5]), 
         .C(rs1[0]), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i8_3_lut (.A(\registers[8] [5]), .B(\registers[9] [5]), 
         .C(rs1[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i8_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i5_3_lut (.A(\registers[6] [5]), .B(\registers[7] [5]), 
         .C(rs1[0]), .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i12_3_lut (.A(\registers[14] [5]), .B(\registers[15] [5]), 
         .C(rs2[0]), .Z(n12_adj_3130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i12_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i11_3_lut (.A(\registers[12] [5]), .B(\registers[13] [5]), 
         .C(rs2[0]), .Z(n11_adj_3131)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i11_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i9_3_lut (.A(\registers[10] [5]), .B(\registers[11] [5]), 
         .C(rs2[0]), .Z(n9_adj_3132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i8_3_lut (.A(\registers[8] [5]), .B(\registers[9] [5]), 
         .C(rs2[0]), .Z(n8_adj_3133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i8_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i5_3_lut (.A(\registers[6] [5]), .B(\registers[7] [5]), 
         .C(rs2[0]), .Z(n5_adj_3134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 i27717_4_lut_4_lut (.A(\registers[2] [7]), .B(rs1[0]), .C(rs1[1]), 
         .D(\registers[1] [7]), .Z(n30426)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i27717_4_lut_4_lut.init = 16'h2c20;
    LUT4 rs2_3__I_0_Mux_3_i12_3_lut (.A(\registers[14] [7]), .B(\registers[15] [7]), 
         .C(rs2[0]), .Z(n12_adj_3135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i12_3_lut.init = 16'hcaca;
    LUT4 i27674_3_lut (.A(\registers[2] [6]), .B(\reg_access[3][2] ), .C(rs2[0]), 
         .Z(n30383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27674_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i11_3_lut (.A(\registers[12] [7]), .B(\registers[13] [7]), 
         .C(rs2[0]), .Z(n11_adj_3136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i9_3_lut (.A(\registers[10] [7]), .B(\registers[11] [7]), 
         .C(rs2[0]), .Z(n9_adj_3137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i8_3_lut (.A(\registers[8] [7]), .B(\registers[9] [7]), 
         .C(rs2[0]), .Z(n8_adj_3138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i12_3_lut (.A(\registers[14] [7]), .B(\registers[15] [7]), 
         .C(rs1[0]), .Z(n12_adj_3139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i12_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i11_3_lut (.A(\registers[12] [7]), .B(\registers[13] [7]), 
         .C(rs1[0]), .Z(n11_adj_3140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i9_3_lut (.A(\registers[10] [7]), .B(\registers[11] [7]), 
         .C(rs1[0]), .Z(n9_adj_3141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i8_3_lut (.A(\registers[8] [7]), .B(\registers[9] [7]), 
         .C(rs1[0]), .Z(n8_adj_3142)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 i15113_2_lut_rep_764 (.A(rd[2]), .B(rd[3]), .Z(n32779)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15113_2_lut_rep_764.init = 16'h8888;
    LUT4 equal_148_i6_2_lut_rep_765 (.A(rd[2]), .B(rd[3]), .Z(n32780)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam equal_148_i6_2_lut_rep_765.init = 16'hbbbb;
    LUT4 equal_143_i6_2_lut_rep_766 (.A(rd[2]), .B(rd[3]), .Z(n32781)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam equal_143_i6_2_lut_rep_766.init = 16'hdddd;
    LUT4 i27680_3_lut (.A(\registers[14] [6]), .B(\registers[15] [6]), .C(rs2[0]), 
         .Z(n30389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27680_3_lut.init = 16'hcaca;
    L6MUX21 i27591 (.D0(n30298), .D1(n30299), .SD(rs2[3]), .Z(data_rs2[0]));
    LUT4 i27679_3_lut (.A(\registers[12] [6]), .B(\registers[13] [6]), .C(rs2[0]), 
         .Z(n30388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27679_3_lut.init = 16'hcaca;
    LUT4 i27678_3_lut (.A(\registers[10] [6]), .B(\registers[11] [6]), .C(rs2[0]), 
         .Z(n30387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27678_3_lut.init = 16'hcaca;
    LUT4 i27673_3_lut (.A(\registers[1] [6]), .B(rs2[0]), .Z(n30382)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27673_3_lut.init = 16'h8888;
    LUT4 i27677_3_lut (.A(\registers[8] [6]), .B(\registers[9] [6]), .C(rs2[0]), 
         .Z(n30386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27677_3_lut.init = 16'hcaca;
    LUT4 i27676_3_lut (.A(\registers[6] [6]), .B(\registers[7] [6]), .C(rs2[0]), 
         .Z(n30385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27676_3_lut.init = 16'hcaca;
    LUT4 i15542_2_lut_rep_771 (.A(rd[3]), .B(rd[2]), .Z(n32786)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15542_2_lut_rep_771.init = 16'heeee;
    LUT4 i27675_3_lut (.A(\registers[5] [6]), .B(rs2[0]), .Z(n30384)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27675_3_lut.init = 16'h8888;
    LUT4 i27665_3_lut (.A(\registers[14] [6]), .B(\registers[15] [6]), .C(rs1[0]), 
         .Z(n30374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27665_3_lut.init = 16'hcaca;
    LUT4 i27664_3_lut (.A(\registers[12] [6]), .B(\registers[13] [6]), .C(rs1[0]), 
         .Z(n30373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27664_3_lut.init = 16'hcaca;
    LUT4 i27663_3_lut (.A(\registers[10] [6]), .B(\registers[11] [6]), .C(rs1[0]), 
         .Z(n30372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27663_3_lut.init = 16'hcaca;
    L6MUX21 i27672 (.D0(n30379), .D1(n30380), .SD(rs1[3]), .Z(data_rs1[2]));
    L6MUX21 i27687 (.D0(n30394), .D1(n30395), .SD(rs2[3]), .Z(data_rs2[2]));
    LUT4 i27662_3_lut (.A(\registers[8] [6]), .B(\registers[9] [6]), .C(rs1[0]), 
         .Z(n30371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27662_3_lut.init = 16'hcaca;
    LUT4 i27661_3_lut (.A(\registers[6] [6]), .B(\registers[7] [6]), .C(rs1[0]), 
         .Z(n30370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27661_3_lut.init = 16'hcaca;
    LUT4 i27660_3_lut (.A(\registers[5] [6]), .B(rs1[0]), .Z(n30369)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27660_3_lut.init = 16'h8888;
    L6MUX21 i27589 (.D0(n30294), .D1(n30295), .SD(rs2[2]), .Z(n30298));
    L6MUX21 i27604 (.D0(n30309), .D1(n30310), .SD(rs1[2]), .Z(n30313));
    FD1S3AX \registers_1[[2__504  (.D(registers_1__2__N_1756), .CK(clk_c), 
            .Q(\registers[1] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[2__504 .GSR = "DISABLED";
    FD1S3AX \registers_1[[1__505  (.D(registers_1__1__N_1757), .CK(clk_c), 
            .Q(\registers[1] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[1__505 .GSR = "DISABLED";
    FD1S3AX \registers_1[[0__506  (.D(registers_1__0__N_1758), .CK(clk_c), 
            .Q(\registers[1] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[0__506 .GSR = "DISABLED";
    FD1S3AX \registers_1[[31__507  (.D(\registers[1] [3]), .CK(clk_c), .Q(return_addr[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[31__507 .GSR = "DISABLED";
    FD1S3AX \registers_1[[30__508  (.D(\registers[1] [2]), .CK(clk_c), .Q(return_addr[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[30__508 .GSR = "DISABLED";
    FD1S3AX \registers_1[[29__509  (.D(\registers[1] [1]), .CK(clk_c), .Q(return_addr[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[29__509 .GSR = "DISABLED";
    FD1S3AX \registers_1[[28__510  (.D(\registers[1] [0]), .CK(clk_c), .Q(return_addr[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[28__510 .GSR = "DISABLED";
    FD1S3AX \registers_1[[27__511  (.D(return_addr[23]), .CK(clk_c), .Q(return_addr[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[27__511 .GSR = "DISABLED";
    FD1S3AX \registers_1[[26__512  (.D(return_addr[22]), .CK(clk_c), .Q(return_addr[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[26__512 .GSR = "DISABLED";
    FD1S3AX \registers_1[[25__513  (.D(return_addr[21]), .CK(clk_c), .Q(return_addr[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[25__513 .GSR = "DISABLED";
    FD1S3AX \registers_1[[24__514  (.D(return_addr[20]), .CK(clk_c), .Q(return_addr[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[24__514 .GSR = "DISABLED";
    FD1S3AX \registers_1[[23__515  (.D(return_addr[19]), .CK(clk_c), .Q(return_addr[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[23__515 .GSR = "DISABLED";
    FD1S3AX \registers_1[[22__516  (.D(return_addr[18]), .CK(clk_c), .Q(return_addr[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[22__516 .GSR = "DISABLED";
    FD1S3AX \registers_1[[21__517  (.D(return_addr[17]), .CK(clk_c), .Q(return_addr[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[21__517 .GSR = "DISABLED";
    FD1S3AX \registers_1[[20__518  (.D(return_addr[16]), .CK(clk_c), .Q(return_addr[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[20__518 .GSR = "DISABLED";
    FD1S3AX \registers_1[[19__519  (.D(return_addr[15]), .CK(clk_c), .Q(return_addr[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[19__519 .GSR = "DISABLED";
    FD1S3AX \registers_1[[18__520  (.D(return_addr[14]), .CK(clk_c), .Q(return_addr[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[18__520 .GSR = "DISABLED";
    FD1S3AX \registers_1[[17__521  (.D(return_addr[13]), .CK(clk_c), .Q(return_addr[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[17__521 .GSR = "DISABLED";
    FD1S3AX \registers_1[[16__522  (.D(return_addr[12]), .CK(clk_c), .Q(return_addr[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[16__522 .GSR = "DISABLED";
    FD1S3AX \registers_1[[15__523  (.D(return_addr[11]), .CK(clk_c), .Q(return_addr[7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[15__523 .GSR = "DISABLED";
    FD1S3AX \registers_1[[14__524  (.D(return_addr[10]), .CK(clk_c), .Q(return_addr[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[14__524 .GSR = "DISABLED";
    FD1S3AX \registers_1[[13__525  (.D(return_addr[9]), .CK(clk_c), .Q(return_addr[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[13__525 .GSR = "DISABLED";
    FD1S3AX \registers_1[[12__526  (.D(return_addr[8]), .CK(clk_c), .Q(return_addr[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[12__526 .GSR = "DISABLED";
    FD1S3AX \registers_1[[11__527  (.D(return_addr[7]), .CK(clk_c), .Q(return_addr[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[11__527 .GSR = "DISABLED";
    FD1S3AX \registers_1[[10__528  (.D(return_addr[6]), .CK(clk_c), .Q(return_addr[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[10__528 .GSR = "DISABLED";
    FD1S3AX \registers_1[[9__529  (.D(return_addr[5]), .CK(clk_c), .Q(return_addr[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[9__529 .GSR = "DISABLED";
    FD1S3AX \registers_1[[8__530  (.D(return_addr[4]), .CK(clk_c), .Q(\registers[1] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[8__530 .GSR = "DISABLED";
    FD1S3AX \registers_1[[7__531  (.D(return_addr[3]), .CK(clk_c), .Q(\registers[1] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[7__531 .GSR = "DISABLED";
    FD1S3AX \registers_1[[6__532  (.D(return_addr[2]), .CK(clk_c), .Q(\registers[1] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[6__532 .GSR = "DISABLED";
    FD1S3AX \registers_1[[5__533  (.D(return_addr[1]), .CK(clk_c), .Q(\registers[1] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[5__533 .GSR = "DISABLED";
    FD1S3AX \registers_1[[4__534  (.D(\registers[1] [8]), .CK(clk_c), .Q(\registers[1] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[4__534 .GSR = "DISABLED";
    FD1S3AX \registers_2[[3__535  (.D(registers_2__3__N_1759), .CK(clk_c), 
            .Q(\registers[2] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[3__535 .GSR = "DISABLED";
    FD1S3AX \registers_2[[2__536  (.D(registers_2__2__N_1762), .CK(clk_c), 
            .Q(\registers[2] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[2__536 .GSR = "DISABLED";
    FD1S3AX \registers_2[[1__537  (.D(registers_2__1__N_1763), .CK(clk_c), 
            .Q(\registers[2] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[1__537 .GSR = "DISABLED";
    FD1S3AX \registers_2[[0__538  (.D(registers_2__0__N_1764), .CK(clk_c), 
            .Q(\registers[2] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[0__538 .GSR = "DISABLED";
    FD1S3AX \registers_2[[31__539  (.D(\registers[2] [3]), .CK(clk_c), .Q(\registers[2] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[31__539 .GSR = "DISABLED";
    FD1S3AX \registers_2[[30__540  (.D(\registers[2] [2]), .CK(clk_c), .Q(\registers[2] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[30__540 .GSR = "DISABLED";
    FD1S3AX \registers_2[[29__541  (.D(\registers[2] [1]), .CK(clk_c), .Q(\registers[2] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[29__541 .GSR = "DISABLED";
    FD1S3AX \registers_2[[28__542  (.D(\registers[2] [0]), .CK(clk_c), .Q(\registers[2] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[28__542 .GSR = "DISABLED";
    FD1S3AX \registers_2[[27__543  (.D(\registers[2] [31]), .CK(clk_c), 
            .Q(\registers[2] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[27__543 .GSR = "DISABLED";
    FD1S3AX \registers_2[[26__544  (.D(\registers[2] [30]), .CK(clk_c), 
            .Q(\registers[2] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[26__544 .GSR = "DISABLED";
    FD1S3AX \registers_2[[25__545  (.D(\registers[2] [29]), .CK(clk_c), 
            .Q(\registers[2] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[25__545 .GSR = "DISABLED";
    FD1S3AX \registers_2[[24__546  (.D(\registers[2] [28]), .CK(clk_c), 
            .Q(\registers[2] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[24__546 .GSR = "DISABLED";
    FD1S3AX \registers_2[[23__547  (.D(\registers[2] [27]), .CK(clk_c), 
            .Q(\registers[2] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[23__547 .GSR = "DISABLED";
    FD1S3AX \registers_2[[22__548  (.D(\registers[2] [26]), .CK(clk_c), 
            .Q(\registers[2] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[22__548 .GSR = "DISABLED";
    FD1S3AX \registers_2[[21__549  (.D(\registers[2] [25]), .CK(clk_c), 
            .Q(\registers[2] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[21__549 .GSR = "DISABLED";
    FD1S3AX \registers_2[[20__550  (.D(\registers[2] [24]), .CK(clk_c), 
            .Q(\registers[2] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[20__550 .GSR = "DISABLED";
    FD1S3AX \registers_2[[19__551  (.D(\registers[2] [23]), .CK(clk_c), 
            .Q(\registers[2] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[19__551 .GSR = "DISABLED";
    FD1S3AX \registers_2[[18__552  (.D(\registers[2] [22]), .CK(clk_c), 
            .Q(\registers[2] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[18__552 .GSR = "DISABLED";
    FD1S3AX \registers_2[[17__553  (.D(\registers[2] [21]), .CK(clk_c), 
            .Q(\registers[2] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[17__553 .GSR = "DISABLED";
    FD1S3AX \registers_2[[16__554  (.D(\registers[2] [20]), .CK(clk_c), 
            .Q(\registers[2] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[16__554 .GSR = "DISABLED";
    FD1S3AX \registers_2[[15__555  (.D(\registers[2] [19]), .CK(clk_c), 
            .Q(\registers[2] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[15__555 .GSR = "DISABLED";
    FD1S3AX \registers_2[[14__556  (.D(\registers[2] [18]), .CK(clk_c), 
            .Q(\registers[2] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[14__556 .GSR = "DISABLED";
    FD1S3AX \registers_2[[13__557  (.D(\registers[2] [17]), .CK(clk_c), 
            .Q(\registers[2] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[13__557 .GSR = "DISABLED";
    FD1S3AX \registers_2[[12__558  (.D(\registers[2] [16]), .CK(clk_c), 
            .Q(\registers[2] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[12__558 .GSR = "DISABLED";
    FD1S3AX \registers_2[[11__559  (.D(\registers[2] [15]), .CK(clk_c), 
            .Q(\registers[2] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[11__559 .GSR = "DISABLED";
    FD1S3AX \registers_2[[10__560  (.D(\registers[2] [14]), .CK(clk_c), 
            .Q(\registers[2] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[10__560 .GSR = "DISABLED";
    FD1S3AX \registers_2[[9__561  (.D(\registers[2] [13]), .CK(clk_c), .Q(\registers[2] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[9__561 .GSR = "DISABLED";
    FD1S3AX \registers_2[[8__562  (.D(\registers[2] [12]), .CK(clk_c), .Q(\registers[2] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[8__562 .GSR = "DISABLED";
    FD1S3AX \registers_2[[7__563  (.D(\registers[2] [11]), .CK(clk_c), .Q(\registers[2] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[7__563 .GSR = "DISABLED";
    FD1S3AX \registers_2[[6__564  (.D(\registers[2] [10]), .CK(clk_c), .Q(\registers[2] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[6__564 .GSR = "DISABLED";
    FD1S3AX \registers_2[[5__565  (.D(\registers[2] [9]), .CK(clk_c), .Q(\registers[2] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[5__565 .GSR = "DISABLED";
    FD1S3AX \registers_2[[4__566  (.D(\registers[2] [8]), .CK(clk_c), .Q(\registers[2] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[4__566 .GSR = "DISABLED";
    FD1S3AX \registers_5[[3__567  (.D(registers_5__3__N_1765), .CK(clk_c), 
            .Q(\registers[5] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[3__567 .GSR = "DISABLED";
    FD1S3AX \registers_5[[2__568  (.D(registers_5__2__N_1768), .CK(clk_c), 
            .Q(\registers[5] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[2__568 .GSR = "DISABLED";
    FD1S3AX \registers_5[[1__569  (.D(registers_5__1__N_1769), .CK(clk_c), 
            .Q(\registers[5] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[1__569 .GSR = "DISABLED";
    FD1S3AX \registers_5[[0__570  (.D(registers_5__0__N_1770), .CK(clk_c), 
            .Q(\registers[5] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[0__570 .GSR = "DISABLED";
    FD1S3AX \registers_5[[31__571  (.D(\registers[5] [3]), .CK(clk_c), .Q(\registers[5] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[31__571 .GSR = "DISABLED";
    FD1S3AX \registers_5[[30__572  (.D(\registers[5] [2]), .CK(clk_c), .Q(\registers[5] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[30__572 .GSR = "DISABLED";
    FD1S3AX \registers_5[[29__573  (.D(\registers[5] [1]), .CK(clk_c), .Q(\registers[5] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[29__573 .GSR = "DISABLED";
    FD1S3AX \registers_5[[28__574  (.D(\registers[5] [0]), .CK(clk_c), .Q(\registers[5] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[28__574 .GSR = "DISABLED";
    FD1S3AX \registers_5[[27__575  (.D(\registers[5] [31]), .CK(clk_c), 
            .Q(\registers[5] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[27__575 .GSR = "DISABLED";
    FD1S3AX \registers_5[[26__576  (.D(\registers[5] [30]), .CK(clk_c), 
            .Q(\registers[5] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[26__576 .GSR = "DISABLED";
    FD1S3AX \registers_5[[25__577  (.D(\registers[5] [29]), .CK(clk_c), 
            .Q(\registers[5] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[25__577 .GSR = "DISABLED";
    FD1S3AX \registers_5[[24__578  (.D(\registers[5] [28]), .CK(clk_c), 
            .Q(\registers[5] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[24__578 .GSR = "DISABLED";
    FD1S3AX \registers_5[[23__579  (.D(\registers[5] [27]), .CK(clk_c), 
            .Q(\registers[5] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[23__579 .GSR = "DISABLED";
    FD1S3AX \registers_5[[22__580  (.D(\registers[5] [26]), .CK(clk_c), 
            .Q(\registers[5] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[22__580 .GSR = "DISABLED";
    FD1S3AX \registers_5[[21__581  (.D(\registers[5] [25]), .CK(clk_c), 
            .Q(\registers[5] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[21__581 .GSR = "DISABLED";
    FD1S3AX \registers_5[[20__582  (.D(\registers[5] [24]), .CK(clk_c), 
            .Q(\registers[5] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[20__582 .GSR = "DISABLED";
    FD1S3AX \registers_5[[19__583  (.D(\registers[5] [23]), .CK(clk_c), 
            .Q(\registers[5] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[19__583 .GSR = "DISABLED";
    FD1S3AX \registers_5[[18__584  (.D(\registers[5] [22]), .CK(clk_c), 
            .Q(\registers[5] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[18__584 .GSR = "DISABLED";
    FD1S3AX \registers_5[[17__585  (.D(\registers[5] [21]), .CK(clk_c), 
            .Q(\registers[5] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[17__585 .GSR = "DISABLED";
    FD1S3AX \registers_5[[16__586  (.D(\registers[5] [20]), .CK(clk_c), 
            .Q(\registers[5] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[16__586 .GSR = "DISABLED";
    FD1S3AX \registers_5[[15__587  (.D(\registers[5] [19]), .CK(clk_c), 
            .Q(\registers[5] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[15__587 .GSR = "DISABLED";
    FD1S3AX \registers_5[[14__588  (.D(\registers[5] [18]), .CK(clk_c), 
            .Q(\registers[5] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[14__588 .GSR = "DISABLED";
    FD1S3AX \registers_5[[13__589  (.D(\registers[5] [17]), .CK(clk_c), 
            .Q(\registers[5] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[13__589 .GSR = "DISABLED";
    FD1S3AX \registers_5[[12__590  (.D(\registers[5] [16]), .CK(clk_c), 
            .Q(\registers[5] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[12__590 .GSR = "DISABLED";
    FD1S3AX \registers_5[[11__591  (.D(\registers[5] [15]), .CK(clk_c), 
            .Q(\registers[5] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[11__591 .GSR = "DISABLED";
    FD1S3AX \registers_5[[10__592  (.D(\registers[5] [14]), .CK(clk_c), 
            .Q(\registers[5] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[10__592 .GSR = "DISABLED";
    FD1S3AX \registers_5[[9__593  (.D(\registers[5] [13]), .CK(clk_c), .Q(\registers[5] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[9__593 .GSR = "DISABLED";
    FD1S3AX \registers_5[[8__594  (.D(\registers[5] [12]), .CK(clk_c), .Q(\registers[5] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[8__594 .GSR = "DISABLED";
    FD1S3AX \registers_5[[7__595  (.D(\registers[5] [11]), .CK(clk_c), .Q(\registers[5] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[7__595 .GSR = "DISABLED";
    FD1S3AX \registers_5[[6__596  (.D(\registers[5] [10]), .CK(clk_c), .Q(\registers[5] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[6__596 .GSR = "DISABLED";
    FD1S3AX \registers_5[[5__597  (.D(\registers[5] [9]), .CK(clk_c), .Q(\registers[5] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[5__597 .GSR = "DISABLED";
    FD1S3AX \registers_5[[4__598  (.D(\registers[5] [8]), .CK(clk_c), .Q(\registers[5] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[4__598 .GSR = "DISABLED";
    FD1S3AX \registers_6[[3__599  (.D(registers_6__3__N_1771), .CK(clk_c), 
            .Q(\registers[6] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[3__599 .GSR = "DISABLED";
    FD1S3AX \registers_6[[2__600  (.D(registers_6__2__N_1774), .CK(clk_c), 
            .Q(\registers[6] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[2__600 .GSR = "DISABLED";
    FD1S3AX \registers_6[[1__601  (.D(registers_6__1__N_1775), .CK(clk_c), 
            .Q(\registers[6] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[1__601 .GSR = "DISABLED";
    FD1S3AX \registers_6[[0__602  (.D(registers_6__0__N_1776), .CK(clk_c), 
            .Q(\registers[6] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[0__602 .GSR = "DISABLED";
    FD1S3AX \registers_6[[31__603  (.D(\registers[6] [3]), .CK(clk_c), .Q(\registers[6] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[31__603 .GSR = "DISABLED";
    FD1S3AX \registers_6[[30__604  (.D(\registers[6] [2]), .CK(clk_c), .Q(\registers[6] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[30__604 .GSR = "DISABLED";
    FD1S3AX \registers_6[[29__605  (.D(\registers[6] [1]), .CK(clk_c), .Q(\registers[6] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[29__605 .GSR = "DISABLED";
    FD1S3AX \registers_6[[28__606  (.D(\registers[6] [0]), .CK(clk_c), .Q(\registers[6] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[28__606 .GSR = "DISABLED";
    FD1S3AX \registers_6[[27__607  (.D(\registers[6] [31]), .CK(clk_c), 
            .Q(\registers[6] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[27__607 .GSR = "DISABLED";
    FD1S3AX \registers_6[[26__608  (.D(\registers[6] [30]), .CK(clk_c), 
            .Q(\registers[6] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[26__608 .GSR = "DISABLED";
    FD1S3AX \registers_6[[25__609  (.D(\registers[6] [29]), .CK(clk_c), 
            .Q(\registers[6] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[25__609 .GSR = "DISABLED";
    FD1S3AX \registers_6[[24__610  (.D(\registers[6] [28]), .CK(clk_c), 
            .Q(\registers[6] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[24__610 .GSR = "DISABLED";
    FD1S3AX \registers_6[[23__611  (.D(\registers[6] [27]), .CK(clk_c), 
            .Q(\registers[6] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[23__611 .GSR = "DISABLED";
    FD1S3AX \registers_6[[22__612  (.D(\registers[6] [26]), .CK(clk_c), 
            .Q(\registers[6] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[22__612 .GSR = "DISABLED";
    FD1S3AX \registers_6[[21__613  (.D(\registers[6] [25]), .CK(clk_c), 
            .Q(\registers[6] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[21__613 .GSR = "DISABLED";
    FD1S3AX \registers_6[[20__614  (.D(\registers[6] [24]), .CK(clk_c), 
            .Q(\registers[6] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[20__614 .GSR = "DISABLED";
    FD1S3AX \registers_6[[19__615  (.D(\registers[6] [23]), .CK(clk_c), 
            .Q(\registers[6] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[19__615 .GSR = "DISABLED";
    FD1S3AX \registers_6[[18__616  (.D(\registers[6] [22]), .CK(clk_c), 
            .Q(\registers[6] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[18__616 .GSR = "DISABLED";
    FD1S3AX \registers_6[[17__617  (.D(\registers[6] [21]), .CK(clk_c), 
            .Q(\registers[6] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[17__617 .GSR = "DISABLED";
    FD1S3AX \registers_6[[16__618  (.D(\registers[6] [20]), .CK(clk_c), 
            .Q(\registers[6] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[16__618 .GSR = "DISABLED";
    FD1S3AX \registers_6[[15__619  (.D(\registers[6] [19]), .CK(clk_c), 
            .Q(\registers[6] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[15__619 .GSR = "DISABLED";
    FD1S3AX \registers_6[[14__620  (.D(\registers[6] [18]), .CK(clk_c), 
            .Q(\registers[6] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[14__620 .GSR = "DISABLED";
    FD1S3AX \registers_6[[13__621  (.D(\registers[6] [17]), .CK(clk_c), 
            .Q(\registers[6] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[13__621 .GSR = "DISABLED";
    FD1S3AX \registers_6[[12__622  (.D(\registers[6] [16]), .CK(clk_c), 
            .Q(\registers[6] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[12__622 .GSR = "DISABLED";
    FD1S3AX \registers_6[[11__623  (.D(\registers[6] [15]), .CK(clk_c), 
            .Q(\registers[6] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[11__623 .GSR = "DISABLED";
    FD1S3AX \registers_6[[10__624  (.D(\registers[6] [14]), .CK(clk_c), 
            .Q(\registers[6] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[10__624 .GSR = "DISABLED";
    FD1S3AX \registers_6[[9__625  (.D(\registers[6] [13]), .CK(clk_c), .Q(\registers[6] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[9__625 .GSR = "DISABLED";
    FD1S3AX \registers_6[[8__626  (.D(\registers[6] [12]), .CK(clk_c), .Q(\registers[6] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[8__626 .GSR = "DISABLED";
    FD1S3AX \registers_6[[7__627  (.D(\registers[6] [11]), .CK(clk_c), .Q(\registers[6] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[7__627 .GSR = "DISABLED";
    FD1S3AX \registers_6[[6__628  (.D(\registers[6] [10]), .CK(clk_c), .Q(\registers[6] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[6__628 .GSR = "DISABLED";
    FD1S3AX \registers_6[[5__629  (.D(\registers[6] [9]), .CK(clk_c), .Q(\registers[6] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[5__629 .GSR = "DISABLED";
    FD1S3AX \registers_6[[4__630  (.D(\registers[6] [8]), .CK(clk_c), .Q(\registers[6] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[4__630 .GSR = "DISABLED";
    FD1S3AX \registers_7[[3__631  (.D(registers_7__3__N_1777), .CK(clk_c), 
            .Q(\registers[7] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[3__631 .GSR = "DISABLED";
    FD1S3AX \registers_7[[2__632  (.D(registers_7__2__N_1780), .CK(clk_c), 
            .Q(\registers[7] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[2__632 .GSR = "DISABLED";
    FD1S3AX \registers_7[[1__633  (.D(registers_7__1__N_1781), .CK(clk_c), 
            .Q(\registers[7] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[1__633 .GSR = "DISABLED";
    FD1S3AX \registers_7[[0__634  (.D(registers_7__0__N_1782), .CK(clk_c), 
            .Q(\registers[7] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[0__634 .GSR = "DISABLED";
    FD1S3AX \registers_7[[31__635  (.D(\registers[7] [3]), .CK(clk_c), .Q(\registers[7] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[31__635 .GSR = "DISABLED";
    FD1S3AX \registers_7[[30__636  (.D(\registers[7] [2]), .CK(clk_c), .Q(\registers[7] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[30__636 .GSR = "DISABLED";
    FD1S3AX \registers_7[[29__637  (.D(\registers[7] [1]), .CK(clk_c), .Q(\registers[7] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[29__637 .GSR = "DISABLED";
    FD1S3AX \registers_7[[28__638  (.D(\registers[7] [0]), .CK(clk_c), .Q(\registers[7] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[28__638 .GSR = "DISABLED";
    FD1S3AX \registers_7[[27__639  (.D(\registers[7] [31]), .CK(clk_c), 
            .Q(\registers[7] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[27__639 .GSR = "DISABLED";
    FD1S3AX \registers_7[[26__640  (.D(\registers[7] [30]), .CK(clk_c), 
            .Q(\registers[7] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[26__640 .GSR = "DISABLED";
    FD1S3AX \registers_7[[25__641  (.D(\registers[7] [29]), .CK(clk_c), 
            .Q(\registers[7] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[25__641 .GSR = "DISABLED";
    FD1S3AX \registers_7[[24__642  (.D(\registers[7] [28]), .CK(clk_c), 
            .Q(\registers[7] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[24__642 .GSR = "DISABLED";
    FD1S3AX \registers_7[[23__643  (.D(\registers[7] [27]), .CK(clk_c), 
            .Q(\registers[7] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[23__643 .GSR = "DISABLED";
    FD1S3AX \registers_7[[22__644  (.D(\registers[7] [26]), .CK(clk_c), 
            .Q(\registers[7] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[22__644 .GSR = "DISABLED";
    FD1S3AX \registers_7[[21__645  (.D(\registers[7] [25]), .CK(clk_c), 
            .Q(\registers[7] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[21__645 .GSR = "DISABLED";
    FD1S3AX \registers_7[[20__646  (.D(\registers[7] [24]), .CK(clk_c), 
            .Q(\registers[7] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[20__646 .GSR = "DISABLED";
    FD1S3AX \registers_7[[19__647  (.D(\registers[7] [23]), .CK(clk_c), 
            .Q(\registers[7] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[19__647 .GSR = "DISABLED";
    FD1S3AX \registers_7[[18__648  (.D(\registers[7] [22]), .CK(clk_c), 
            .Q(\registers[7] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[18__648 .GSR = "DISABLED";
    FD1S3AX \registers_7[[17__649  (.D(\registers[7] [21]), .CK(clk_c), 
            .Q(\registers[7] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[17__649 .GSR = "DISABLED";
    FD1S3AX \registers_7[[16__650  (.D(\registers[7] [20]), .CK(clk_c), 
            .Q(\registers[7] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[16__650 .GSR = "DISABLED";
    FD1S3AX \registers_7[[15__651  (.D(\registers[7] [19]), .CK(clk_c), 
            .Q(\registers[7] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[15__651 .GSR = "DISABLED";
    FD1S3AX \registers_7[[14__652  (.D(\registers[7] [18]), .CK(clk_c), 
            .Q(\registers[7] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[14__652 .GSR = "DISABLED";
    FD1S3AX \registers_7[[13__653  (.D(\registers[7] [17]), .CK(clk_c), 
            .Q(\registers[7] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[13__653 .GSR = "DISABLED";
    FD1S3AX \registers_7[[12__654  (.D(\registers[7] [16]), .CK(clk_c), 
            .Q(\registers[7] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[12__654 .GSR = "DISABLED";
    FD1S3AX \registers_7[[11__655  (.D(\registers[7] [15]), .CK(clk_c), 
            .Q(\registers[7] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[11__655 .GSR = "DISABLED";
    FD1S3AX \registers_7[[10__656  (.D(\registers[7] [14]), .CK(clk_c), 
            .Q(\registers[7] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[10__656 .GSR = "DISABLED";
    FD1S3AX \registers_7[[9__657  (.D(\registers[7] [13]), .CK(clk_c), .Q(\registers[7] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[9__657 .GSR = "DISABLED";
    FD1S3AX \registers_7[[8__658  (.D(\registers[7] [12]), .CK(clk_c), .Q(\registers[7] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[8__658 .GSR = "DISABLED";
    FD1S3AX \registers_7[[7__659  (.D(\registers[7] [11]), .CK(clk_c), .Q(\registers[7] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[7__659 .GSR = "DISABLED";
    FD1S3AX \registers_7[[6__660  (.D(\registers[7] [10]), .CK(clk_c), .Q(\registers[7] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[6__660 .GSR = "DISABLED";
    FD1S3AX \registers_7[[5__661  (.D(\registers[7] [9]), .CK(clk_c), .Q(\registers[7] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[5__661 .GSR = "DISABLED";
    FD1S3AX \registers_7[[4__662  (.D(\registers[7] [8]), .CK(clk_c), .Q(\registers[7] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[4__662 .GSR = "DISABLED";
    FD1S3AX \registers_8[[3__663  (.D(registers_8__3__N_1783), .CK(clk_c), 
            .Q(\registers[8] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[3__663 .GSR = "DISABLED";
    FD1S3AX \registers_8[[2__664  (.D(registers_8__2__N_1786), .CK(clk_c), 
            .Q(\registers[8] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[2__664 .GSR = "DISABLED";
    FD1S3AX \registers_8[[1__665  (.D(registers_8__1__N_1787), .CK(clk_c), 
            .Q(\registers[8] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[1__665 .GSR = "DISABLED";
    FD1S3AX \registers_8[[0__666  (.D(registers_8__0__N_1788), .CK(clk_c), 
            .Q(\registers[8] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[0__666 .GSR = "DISABLED";
    FD1S3AX \registers_8[[31__667  (.D(\registers[8] [3]), .CK(clk_c), .Q(\registers[8] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[31__667 .GSR = "DISABLED";
    FD1S3AX \registers_8[[30__668  (.D(\registers[8] [2]), .CK(clk_c), .Q(\registers[8] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[30__668 .GSR = "DISABLED";
    FD1S3AX \registers_8[[29__669  (.D(\registers[8] [1]), .CK(clk_c), .Q(\registers[8] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[29__669 .GSR = "DISABLED";
    FD1S3AX \registers_8[[28__670  (.D(\registers[8] [0]), .CK(clk_c), .Q(\registers[8] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[28__670 .GSR = "DISABLED";
    FD1S3AX \registers_8[[27__671  (.D(\registers[8] [31]), .CK(clk_c), 
            .Q(\registers[8] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[27__671 .GSR = "DISABLED";
    FD1S3AX \registers_8[[26__672  (.D(\registers[8] [30]), .CK(clk_c), 
            .Q(\registers[8] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[26__672 .GSR = "DISABLED";
    FD1S3AX \registers_8[[25__673  (.D(\registers[8] [29]), .CK(clk_c), 
            .Q(\registers[8] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[25__673 .GSR = "DISABLED";
    FD1S3AX \registers_8[[24__674  (.D(\registers[8] [28]), .CK(clk_c), 
            .Q(\registers[8] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[24__674 .GSR = "DISABLED";
    FD1S3AX \registers_8[[23__675  (.D(\registers[8] [27]), .CK(clk_c), 
            .Q(\registers[8] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[23__675 .GSR = "DISABLED";
    FD1S3AX \registers_8[[22__676  (.D(\registers[8] [26]), .CK(clk_c), 
            .Q(\registers[8] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[22__676 .GSR = "DISABLED";
    FD1S3AX \registers_8[[21__677  (.D(\registers[8] [25]), .CK(clk_c), 
            .Q(\registers[8] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[21__677 .GSR = "DISABLED";
    FD1S3AX \registers_8[[20__678  (.D(\registers[8] [24]), .CK(clk_c), 
            .Q(\registers[8] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[20__678 .GSR = "DISABLED";
    FD1S3AX \registers_8[[19__679  (.D(\registers[8] [23]), .CK(clk_c), 
            .Q(\registers[8] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[19__679 .GSR = "DISABLED";
    FD1S3AX \registers_8[[18__680  (.D(\registers[8] [22]), .CK(clk_c), 
            .Q(\registers[8] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[18__680 .GSR = "DISABLED";
    FD1S3AX \registers_8[[17__681  (.D(\registers[8] [21]), .CK(clk_c), 
            .Q(\registers[8] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[17__681 .GSR = "DISABLED";
    FD1S3AX \registers_8[[16__682  (.D(\registers[8] [20]), .CK(clk_c), 
            .Q(\registers[8] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[16__682 .GSR = "DISABLED";
    FD1S3AX \registers_8[[15__683  (.D(\registers[8] [19]), .CK(clk_c), 
            .Q(\registers[8] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[15__683 .GSR = "DISABLED";
    FD1S3AX \registers_8[[14__684  (.D(\registers[8] [18]), .CK(clk_c), 
            .Q(\registers[8] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[14__684 .GSR = "DISABLED";
    FD1S3AX \registers_8[[13__685  (.D(\registers[8] [17]), .CK(clk_c), 
            .Q(\registers[8] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[13__685 .GSR = "DISABLED";
    FD1S3AX \registers_8[[12__686  (.D(\registers[8] [16]), .CK(clk_c), 
            .Q(\registers[8] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[12__686 .GSR = "DISABLED";
    FD1S3AX \registers_8[[11__687  (.D(\registers[8] [15]), .CK(clk_c), 
            .Q(\registers[8] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[11__687 .GSR = "DISABLED";
    FD1S3AX \registers_8[[10__688  (.D(\registers[8] [14]), .CK(clk_c), 
            .Q(\registers[8] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[10__688 .GSR = "DISABLED";
    FD1S3AX \registers_8[[9__689  (.D(\registers[8] [13]), .CK(clk_c), .Q(\registers[8] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[9__689 .GSR = "DISABLED";
    FD1S3AX \registers_8[[8__690  (.D(\registers[8] [12]), .CK(clk_c), .Q(\registers[8] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[8__690 .GSR = "DISABLED";
    FD1S3AX \registers_8[[7__691  (.D(\registers[8] [11]), .CK(clk_c), .Q(\registers[8] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[7__691 .GSR = "DISABLED";
    FD1S3AX \registers_8[[6__692  (.D(\registers[8] [10]), .CK(clk_c), .Q(\registers[8] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[6__692 .GSR = "DISABLED";
    FD1S3AX \registers_8[[5__693  (.D(\registers[8] [9]), .CK(clk_c), .Q(\registers[8] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[5__693 .GSR = "DISABLED";
    FD1S3AX \registers_8[[4__694  (.D(\registers[8] [8]), .CK(clk_c), .Q(\registers[8] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[4__694 .GSR = "DISABLED";
    FD1S3AX \registers_9[[3__695  (.D(registers_9__3__N_1789), .CK(clk_c), 
            .Q(\registers[9] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[3__695 .GSR = "DISABLED";
    FD1S3AX \registers_9[[2__696  (.D(registers_9__2__N_1792), .CK(clk_c), 
            .Q(\registers[9] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[2__696 .GSR = "DISABLED";
    FD1S3AX \registers_9[[1__697  (.D(registers_9__1__N_1793), .CK(clk_c), 
            .Q(\registers[9] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[1__697 .GSR = "DISABLED";
    FD1S3AX \registers_9[[0__698  (.D(registers_9__0__N_1794), .CK(clk_c), 
            .Q(\registers[9] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[0__698 .GSR = "DISABLED";
    FD1S3AX \registers_9[[31__699  (.D(\registers[9] [3]), .CK(clk_c), .Q(\registers[9] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[31__699 .GSR = "DISABLED";
    FD1S3AX \registers_9[[30__700  (.D(\registers[9] [2]), .CK(clk_c), .Q(\registers[9] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[30__700 .GSR = "DISABLED";
    FD1S3AX \registers_9[[29__701  (.D(\registers[9] [1]), .CK(clk_c), .Q(\registers[9] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[29__701 .GSR = "DISABLED";
    FD1S3AX \registers_9[[28__702  (.D(\registers[9] [0]), .CK(clk_c), .Q(\registers[9] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[28__702 .GSR = "DISABLED";
    FD1S3AX \registers_9[[27__703  (.D(\registers[9] [31]), .CK(clk_c), 
            .Q(\registers[9] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[27__703 .GSR = "DISABLED";
    FD1S3AX \registers_9[[26__704  (.D(\registers[9] [30]), .CK(clk_c), 
            .Q(\registers[9] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[26__704 .GSR = "DISABLED";
    FD1S3AX \registers_9[[25__705  (.D(\registers[9] [29]), .CK(clk_c), 
            .Q(\registers[9] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[25__705 .GSR = "DISABLED";
    FD1S3AX \registers_9[[24__706  (.D(\registers[9] [28]), .CK(clk_c), 
            .Q(\registers[9] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[24__706 .GSR = "DISABLED";
    FD1S3AX \registers_9[[23__707  (.D(\registers[9] [27]), .CK(clk_c), 
            .Q(\registers[9] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[23__707 .GSR = "DISABLED";
    FD1S3AX \registers_9[[22__708  (.D(\registers[9] [26]), .CK(clk_c), 
            .Q(\registers[9] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[22__708 .GSR = "DISABLED";
    FD1S3AX \registers_9[[21__709  (.D(\registers[9] [25]), .CK(clk_c), 
            .Q(\registers[9] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[21__709 .GSR = "DISABLED";
    FD1S3AX \registers_9[[20__710  (.D(\registers[9] [24]), .CK(clk_c), 
            .Q(\registers[9] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[20__710 .GSR = "DISABLED";
    FD1S3AX \registers_9[[19__711  (.D(\registers[9] [23]), .CK(clk_c), 
            .Q(\registers[9] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[19__711 .GSR = "DISABLED";
    FD1S3AX \registers_9[[18__712  (.D(\registers[9] [22]), .CK(clk_c), 
            .Q(\registers[9] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[18__712 .GSR = "DISABLED";
    FD1S3AX \registers_9[[17__713  (.D(\registers[9] [21]), .CK(clk_c), 
            .Q(\registers[9] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[17__713 .GSR = "DISABLED";
    FD1S3AX \registers_9[[16__714  (.D(\registers[9] [20]), .CK(clk_c), 
            .Q(\registers[9] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[16__714 .GSR = "DISABLED";
    FD1S3AX \registers_9[[15__715  (.D(\registers[9] [19]), .CK(clk_c), 
            .Q(\registers[9] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[15__715 .GSR = "DISABLED";
    FD1S3AX \registers_9[[14__716  (.D(\registers[9] [18]), .CK(clk_c), 
            .Q(\registers[9] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[14__716 .GSR = "DISABLED";
    FD1S3AX \registers_9[[13__717  (.D(\registers[9] [17]), .CK(clk_c), 
            .Q(\registers[9] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[13__717 .GSR = "DISABLED";
    FD1S3AX \registers_9[[12__718  (.D(\registers[9] [16]), .CK(clk_c), 
            .Q(\registers[9] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[12__718 .GSR = "DISABLED";
    FD1S3AX \registers_9[[11__719  (.D(\registers[9] [15]), .CK(clk_c), 
            .Q(\registers[9] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[11__719 .GSR = "DISABLED";
    FD1S3AX \registers_9[[10__720  (.D(\registers[9] [14]), .CK(clk_c), 
            .Q(\registers[9] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[10__720 .GSR = "DISABLED";
    FD1S3AX \registers_9[[9__721  (.D(\registers[9] [13]), .CK(clk_c), .Q(\registers[9] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[9__721 .GSR = "DISABLED";
    FD1S3AX \registers_9[[8__722  (.D(\registers[9] [12]), .CK(clk_c), .Q(\registers[9] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[8__722 .GSR = "DISABLED";
    FD1S3AX \registers_9[[7__723  (.D(\registers[9] [11]), .CK(clk_c), .Q(\registers[9] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[7__723 .GSR = "DISABLED";
    FD1S3AX \registers_9[[6__724  (.D(\registers[9] [10]), .CK(clk_c), .Q(\registers[9] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[6__724 .GSR = "DISABLED";
    FD1S3AX \registers_9[[5__725  (.D(\registers[9] [9]), .CK(clk_c), .Q(\registers[9] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[5__725 .GSR = "DISABLED";
    FD1S3AX \registers_9[[4__726  (.D(\registers[9] [8]), .CK(clk_c), .Q(\registers[9] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[4__726 .GSR = "DISABLED";
    FD1S3AX \registers_10[[3__727  (.D(registers_10__3__N_1795), .CK(clk_c), 
            .Q(\registers[10] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[3__727 .GSR = "DISABLED";
    FD1S3AX \registers_10[[2__728  (.D(registers_10__2__N_1798), .CK(clk_c), 
            .Q(\registers[10] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[2__728 .GSR = "DISABLED";
    FD1S3AX \registers_10[[1__729  (.D(registers_10__1__N_1799), .CK(clk_c), 
            .Q(\registers[10] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[1__729 .GSR = "DISABLED";
    FD1S3AX \registers_10[[0__730  (.D(registers_10__0__N_1800), .CK(clk_c), 
            .Q(\registers[10] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[0__730 .GSR = "DISABLED";
    FD1S3AX \registers_10[[31__731  (.D(\registers[10] [3]), .CK(clk_c), 
            .Q(\registers[10] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[31__731 .GSR = "DISABLED";
    FD1S3AX \registers_10[[30__732  (.D(\registers[10] [2]), .CK(clk_c), 
            .Q(\registers[10] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[30__732 .GSR = "DISABLED";
    FD1S3AX \registers_10[[29__733  (.D(\registers[10] [1]), .CK(clk_c), 
            .Q(\registers[10] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[29__733 .GSR = "DISABLED";
    FD1S3AX \registers_10[[28__734  (.D(\registers[10] [0]), .CK(clk_c), 
            .Q(\registers[10] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[28__734 .GSR = "DISABLED";
    FD1S3AX \registers_10[[27__735  (.D(\registers[10] [31]), .CK(clk_c), 
            .Q(\registers[10] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[27__735 .GSR = "DISABLED";
    FD1S3AX \registers_10[[26__736  (.D(\registers[10] [30]), .CK(clk_c), 
            .Q(\registers[10] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[26__736 .GSR = "DISABLED";
    FD1S3AX \registers_10[[25__737  (.D(\registers[10] [29]), .CK(clk_c), 
            .Q(\registers[10] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[25__737 .GSR = "DISABLED";
    FD1S3AX \registers_10[[24__738  (.D(\registers[10] [28]), .CK(clk_c), 
            .Q(\registers[10] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[24__738 .GSR = "DISABLED";
    FD1S3AX \registers_10[[23__739  (.D(\registers[10] [27]), .CK(clk_c), 
            .Q(\registers[10] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[23__739 .GSR = "DISABLED";
    FD1S3AX \registers_10[[22__740  (.D(\registers[10] [26]), .CK(clk_c), 
            .Q(\registers[10] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[22__740 .GSR = "DISABLED";
    FD1S3AX \registers_10[[21__741  (.D(\registers[10] [25]), .CK(clk_c), 
            .Q(\registers[10] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[21__741 .GSR = "DISABLED";
    FD1S3AX \registers_10[[20__742  (.D(\registers[10] [24]), .CK(clk_c), 
            .Q(\registers[10] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[20__742 .GSR = "DISABLED";
    FD1S3AX \registers_10[[19__743  (.D(\registers[10] [23]), .CK(clk_c), 
            .Q(\registers[10] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[19__743 .GSR = "DISABLED";
    FD1S3AX \registers_10[[18__744  (.D(\registers[10] [22]), .CK(clk_c), 
            .Q(\registers[10] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[18__744 .GSR = "DISABLED";
    FD1S3AX \registers_10[[17__745  (.D(\registers[10] [21]), .CK(clk_c), 
            .Q(\registers[10] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[17__745 .GSR = "DISABLED";
    FD1S3AX \registers_10[[16__746  (.D(\registers[10] [20]), .CK(clk_c), 
            .Q(\registers[10] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[16__746 .GSR = "DISABLED";
    FD1S3AX \registers_10[[15__747  (.D(\registers[10] [19]), .CK(clk_c), 
            .Q(\registers[10] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[15__747 .GSR = "DISABLED";
    FD1S3AX \registers_10[[14__748  (.D(\registers[10] [18]), .CK(clk_c), 
            .Q(\registers[10] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[14__748 .GSR = "DISABLED";
    FD1S3AX \registers_10[[13__749  (.D(\registers[10] [17]), .CK(clk_c), 
            .Q(\registers[10] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[13__749 .GSR = "DISABLED";
    FD1S3AX \registers_10[[12__750  (.D(\registers[10] [16]), .CK(clk_c), 
            .Q(\registers[10] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[12__750 .GSR = "DISABLED";
    FD1S3AX \registers_10[[11__751  (.D(\registers[10] [15]), .CK(clk_c), 
            .Q(\registers[10] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[11__751 .GSR = "DISABLED";
    FD1S3AX \registers_10[[10__752  (.D(\registers[10] [14]), .CK(clk_c), 
            .Q(\registers[10] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[10__752 .GSR = "DISABLED";
    FD1S3AX \registers_10[[9__753  (.D(\registers[10] [13]), .CK(clk_c), 
            .Q(\registers[10] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[9__753 .GSR = "DISABLED";
    FD1S3AX \registers_10[[8__754  (.D(\registers[10] [12]), .CK(clk_c), 
            .Q(\registers[10] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[8__754 .GSR = "DISABLED";
    FD1S3AX \registers_10[[7__755  (.D(\registers[10] [11]), .CK(clk_c), 
            .Q(\registers[10] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[7__755 .GSR = "DISABLED";
    FD1S3AX \registers_10[[6__756  (.D(\registers[10] [10]), .CK(clk_c), 
            .Q(\registers[10] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[6__756 .GSR = "DISABLED";
    FD1S3AX \registers_10[[5__757  (.D(\registers[10] [9]), .CK(clk_c), 
            .Q(\registers[10] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[5__757 .GSR = "DISABLED";
    FD1S3AX \registers_10[[4__758  (.D(\registers[10] [8]), .CK(clk_c), 
            .Q(\registers[10] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[4__758 .GSR = "DISABLED";
    FD1S3AX \registers_11[[3__759  (.D(registers_11__3__N_1801), .CK(clk_c), 
            .Q(\registers[11] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[3__759 .GSR = "DISABLED";
    FD1S3AX \registers_11[[2__760  (.D(registers_11__2__N_1804), .CK(clk_c), 
            .Q(\registers[11] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[2__760 .GSR = "DISABLED";
    FD1S3AX \registers_11[[1__761  (.D(registers_11__1__N_1805), .CK(clk_c), 
            .Q(\registers[11] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[1__761 .GSR = "DISABLED";
    FD1S3AX \registers_11[[0__762  (.D(registers_11__0__N_1806), .CK(clk_c), 
            .Q(\registers[11] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[0__762 .GSR = "DISABLED";
    FD1S3AX \registers_11[[31__763  (.D(\registers[11] [3]), .CK(clk_c), 
            .Q(\registers[11] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[31__763 .GSR = "DISABLED";
    FD1S3AX \registers_11[[30__764  (.D(\registers[11] [2]), .CK(clk_c), 
            .Q(\registers[11] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[30__764 .GSR = "DISABLED";
    FD1S3AX \registers_11[[29__765  (.D(\registers[11] [1]), .CK(clk_c), 
            .Q(\registers[11] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[29__765 .GSR = "DISABLED";
    FD1S3AX \registers_11[[28__766  (.D(\registers[11] [0]), .CK(clk_c), 
            .Q(\registers[11] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[28__766 .GSR = "DISABLED";
    FD1S3AX \registers_11[[27__767  (.D(\registers[11] [31]), .CK(clk_c), 
            .Q(\registers[11] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[27__767 .GSR = "DISABLED";
    FD1S3AX \registers_11[[26__768  (.D(\registers[11] [30]), .CK(clk_c), 
            .Q(\registers[11] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[26__768 .GSR = "DISABLED";
    FD1S3AX \registers_11[[25__769  (.D(\registers[11] [29]), .CK(clk_c), 
            .Q(\registers[11] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[25__769 .GSR = "DISABLED";
    FD1S3AX \registers_11[[24__770  (.D(\registers[11] [28]), .CK(clk_c), 
            .Q(\registers[11] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[24__770 .GSR = "DISABLED";
    FD1S3AX \registers_11[[23__771  (.D(\registers[11] [27]), .CK(clk_c), 
            .Q(\registers[11] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[23__771 .GSR = "DISABLED";
    FD1S3AX \registers_11[[22__772  (.D(\registers[11] [26]), .CK(clk_c), 
            .Q(\registers[11] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[22__772 .GSR = "DISABLED";
    FD1S3AX \registers_11[[21__773  (.D(\registers[11] [25]), .CK(clk_c), 
            .Q(\registers[11] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[21__773 .GSR = "DISABLED";
    FD1S3AX \registers_11[[20__774  (.D(\registers[11] [24]), .CK(clk_c), 
            .Q(\registers[11] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[20__774 .GSR = "DISABLED";
    FD1S3AX \registers_11[[19__775  (.D(\registers[11] [23]), .CK(clk_c), 
            .Q(\registers[11] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[19__775 .GSR = "DISABLED";
    FD1S3AX \registers_11[[18__776  (.D(\registers[11] [22]), .CK(clk_c), 
            .Q(\registers[11] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[18__776 .GSR = "DISABLED";
    FD1S3AX \registers_11[[17__777  (.D(\registers[11] [21]), .CK(clk_c), 
            .Q(\registers[11] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[17__777 .GSR = "DISABLED";
    FD1S3AX \registers_11[[16__778  (.D(\registers[11] [20]), .CK(clk_c), 
            .Q(\registers[11] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[16__778 .GSR = "DISABLED";
    FD1S3AX \registers_11[[15__779  (.D(\registers[11] [19]), .CK(clk_c), 
            .Q(\registers[11] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[15__779 .GSR = "DISABLED";
    FD1S3AX \registers_11[[14__780  (.D(\registers[11] [18]), .CK(clk_c), 
            .Q(\registers[11] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[14__780 .GSR = "DISABLED";
    FD1S3AX \registers_11[[13__781  (.D(\registers[11] [17]), .CK(clk_c), 
            .Q(\registers[11] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[13__781 .GSR = "DISABLED";
    FD1S3AX \registers_11[[12__782  (.D(\registers[11] [16]), .CK(clk_c), 
            .Q(\registers[11] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[12__782 .GSR = "DISABLED";
    FD1S3AX \registers_11[[11__783  (.D(\registers[11] [15]), .CK(clk_c), 
            .Q(\registers[11] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[11__783 .GSR = "DISABLED";
    FD1S3AX \registers_11[[10__784  (.D(\registers[11] [14]), .CK(clk_c), 
            .Q(\registers[11] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[10__784 .GSR = "DISABLED";
    FD1S3AX \registers_11[[9__785  (.D(\registers[11] [13]), .CK(clk_c), 
            .Q(\registers[11] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[9__785 .GSR = "DISABLED";
    FD1S3AX \registers_11[[8__786  (.D(\registers[11] [12]), .CK(clk_c), 
            .Q(\registers[11] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[8__786 .GSR = "DISABLED";
    FD1S3AX \registers_11[[7__787  (.D(\registers[11] [11]), .CK(clk_c), 
            .Q(\registers[11] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[7__787 .GSR = "DISABLED";
    FD1S3AX \registers_11[[6__788  (.D(\registers[11] [10]), .CK(clk_c), 
            .Q(\registers[11] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[6__788 .GSR = "DISABLED";
    FD1S3AX \registers_11[[5__789  (.D(\registers[11] [9]), .CK(clk_c), 
            .Q(\registers[11] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[5__789 .GSR = "DISABLED";
    FD1S3AX \registers_11[[4__790  (.D(\registers[11] [8]), .CK(clk_c), 
            .Q(\registers[11] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[4__790 .GSR = "DISABLED";
    FD1S3AX \registers_12[[3__791  (.D(registers_12__3__N_1807), .CK(clk_c), 
            .Q(\registers[12] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[3__791 .GSR = "DISABLED";
    FD1S3AX \registers_12[[2__792  (.D(registers_12__2__N_1810), .CK(clk_c), 
            .Q(\registers[12] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[2__792 .GSR = "DISABLED";
    FD1S3AX \registers_12[[1__793  (.D(registers_12__1__N_1811), .CK(clk_c), 
            .Q(\registers[12] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[1__793 .GSR = "DISABLED";
    FD1S3AX \registers_12[[0__794  (.D(registers_12__0__N_1812), .CK(clk_c), 
            .Q(\registers[12] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[0__794 .GSR = "DISABLED";
    FD1S3AX \registers_12[[31__795  (.D(\registers[12] [3]), .CK(clk_c), 
            .Q(\registers[12] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[31__795 .GSR = "DISABLED";
    FD1S3AX \registers_12[[30__796  (.D(\registers[12] [2]), .CK(clk_c), 
            .Q(\registers[12] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[30__796 .GSR = "DISABLED";
    FD1S3AX \registers_12[[29__797  (.D(\registers[12] [1]), .CK(clk_c), 
            .Q(\registers[12] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[29__797 .GSR = "DISABLED";
    FD1S3AX \registers_12[[28__798  (.D(\registers[12] [0]), .CK(clk_c), 
            .Q(\registers[12] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[28__798 .GSR = "DISABLED";
    FD1S3AX \registers_12[[27__799  (.D(\registers[12] [31]), .CK(clk_c), 
            .Q(\registers[12] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[27__799 .GSR = "DISABLED";
    FD1S3AX \registers_12[[26__800  (.D(\registers[12] [30]), .CK(clk_c), 
            .Q(\registers[12] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[26__800 .GSR = "DISABLED";
    FD1S3AX \registers_12[[25__801  (.D(\registers[12] [29]), .CK(clk_c), 
            .Q(\registers[12] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[25__801 .GSR = "DISABLED";
    FD1S3AX \registers_12[[24__802  (.D(\registers[12] [28]), .CK(clk_c), 
            .Q(\registers[12] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[24__802 .GSR = "DISABLED";
    FD1S3AX \registers_12[[23__803  (.D(\registers[12] [27]), .CK(clk_c), 
            .Q(\registers[12] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[23__803 .GSR = "DISABLED";
    FD1S3AX \registers_12[[22__804  (.D(\registers[12] [26]), .CK(clk_c), 
            .Q(\registers[12] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[22__804 .GSR = "DISABLED";
    FD1S3AX \registers_12[[21__805  (.D(\registers[12] [25]), .CK(clk_c), 
            .Q(\registers[12] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[21__805 .GSR = "DISABLED";
    FD1S3AX \registers_12[[20__806  (.D(\registers[12] [24]), .CK(clk_c), 
            .Q(\registers[12] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[20__806 .GSR = "DISABLED";
    FD1S3AX \registers_12[[19__807  (.D(\registers[12] [23]), .CK(clk_c), 
            .Q(\registers[12] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[19__807 .GSR = "DISABLED";
    FD1S3AX \registers_12[[18__808  (.D(\registers[12] [22]), .CK(clk_c), 
            .Q(\registers[12] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[18__808 .GSR = "DISABLED";
    FD1S3AX \registers_12[[17__809  (.D(\registers[12] [21]), .CK(clk_c), 
            .Q(\registers[12] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[17__809 .GSR = "DISABLED";
    FD1S3AX \registers_12[[16__810  (.D(\registers[12] [20]), .CK(clk_c), 
            .Q(\registers[12] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[16__810 .GSR = "DISABLED";
    FD1S3AX \registers_12[[15__811  (.D(\registers[12] [19]), .CK(clk_c), 
            .Q(\registers[12] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[15__811 .GSR = "DISABLED";
    FD1S3AX \registers_12[[14__812  (.D(\registers[12] [18]), .CK(clk_c), 
            .Q(\registers[12] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[14__812 .GSR = "DISABLED";
    FD1S3AX \registers_12[[13__813  (.D(\registers[12] [17]), .CK(clk_c), 
            .Q(\registers[12] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[13__813 .GSR = "DISABLED";
    FD1S3AX \registers_12[[12__814  (.D(\registers[12] [16]), .CK(clk_c), 
            .Q(\registers[12] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[12__814 .GSR = "DISABLED";
    FD1S3AX \registers_12[[11__815  (.D(\registers[12] [15]), .CK(clk_c), 
            .Q(\registers[12] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[11__815 .GSR = "DISABLED";
    FD1S3AX \registers_12[[10__816  (.D(\registers[12] [14]), .CK(clk_c), 
            .Q(\registers[12] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[10__816 .GSR = "DISABLED";
    FD1S3AX \registers_12[[9__817  (.D(\registers[12] [13]), .CK(clk_c), 
            .Q(\registers[12] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[9__817 .GSR = "DISABLED";
    FD1S3AX \registers_12[[8__818  (.D(\registers[12] [12]), .CK(clk_c), 
            .Q(\registers[12] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[8__818 .GSR = "DISABLED";
    FD1S3AX \registers_12[[7__819  (.D(\registers[12] [11]), .CK(clk_c), 
            .Q(\registers[12] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[7__819 .GSR = "DISABLED";
    FD1S3AX \registers_12[[6__820  (.D(\registers[12] [10]), .CK(clk_c), 
            .Q(\registers[12] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[6__820 .GSR = "DISABLED";
    FD1S3AX \registers_12[[5__821  (.D(\registers[12] [9]), .CK(clk_c), 
            .Q(\registers[12] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[5__821 .GSR = "DISABLED";
    FD1S3AX \registers_12[[4__822  (.D(\registers[12] [8]), .CK(clk_c), 
            .Q(\registers[12] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[4__822 .GSR = "DISABLED";
    FD1S3AX \registers_13[[3__823  (.D(registers_13__3__N_1813), .CK(clk_c), 
            .Q(\registers[13] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[3__823 .GSR = "DISABLED";
    FD1S3AX \registers_13[[2__824  (.D(registers_13__2__N_1816), .CK(clk_c), 
            .Q(\registers[13] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[2__824 .GSR = "DISABLED";
    FD1S3AX \registers_13[[1__825  (.D(registers_13__1__N_1817), .CK(clk_c), 
            .Q(\registers[13] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[1__825 .GSR = "DISABLED";
    FD1S3AX \registers_13[[0__826  (.D(registers_13__0__N_1818), .CK(clk_c), 
            .Q(\registers[13] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[0__826 .GSR = "DISABLED";
    FD1S3AX \registers_13[[31__827  (.D(\registers[13] [3]), .CK(clk_c), 
            .Q(\registers[13] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[31__827 .GSR = "DISABLED";
    FD1S3AX \registers_13[[30__828  (.D(\registers[13] [2]), .CK(clk_c), 
            .Q(\registers[13] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[30__828 .GSR = "DISABLED";
    FD1S3AX \registers_13[[29__829  (.D(\registers[13] [1]), .CK(clk_c), 
            .Q(\registers[13] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[29__829 .GSR = "DISABLED";
    FD1S3AX \registers_13[[28__830  (.D(\registers[13] [0]), .CK(clk_c), 
            .Q(\registers[13] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[28__830 .GSR = "DISABLED";
    FD1S3AX \registers_13[[27__831  (.D(\registers[13] [31]), .CK(clk_c), 
            .Q(\registers[13] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[27__831 .GSR = "DISABLED";
    FD1S3AX \registers_13[[26__832  (.D(\registers[13] [30]), .CK(clk_c), 
            .Q(\registers[13] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[26__832 .GSR = "DISABLED";
    FD1S3AX \registers_13[[25__833  (.D(\registers[13] [29]), .CK(clk_c), 
            .Q(\registers[13] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[25__833 .GSR = "DISABLED";
    FD1S3AX \registers_13[[24__834  (.D(\registers[13] [28]), .CK(clk_c), 
            .Q(\registers[13] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[24__834 .GSR = "DISABLED";
    FD1S3AX \registers_13[[23__835  (.D(\registers[13] [27]), .CK(clk_c), 
            .Q(\registers[13] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[23__835 .GSR = "DISABLED";
    FD1S3AX \registers_13[[22__836  (.D(\registers[13] [26]), .CK(clk_c), 
            .Q(\registers[13] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[22__836 .GSR = "DISABLED";
    FD1S3AX \registers_13[[21__837  (.D(\registers[13] [25]), .CK(clk_c), 
            .Q(\registers[13] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[21__837 .GSR = "DISABLED";
    FD1S3AX \registers_13[[20__838  (.D(\registers[13] [24]), .CK(clk_c), 
            .Q(\registers[13] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[20__838 .GSR = "DISABLED";
    FD1S3AX \registers_13[[19__839  (.D(\registers[13] [23]), .CK(clk_c), 
            .Q(\registers[13] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[19__839 .GSR = "DISABLED";
    FD1S3AX \registers_13[[18__840  (.D(\registers[13] [22]), .CK(clk_c), 
            .Q(\registers[13] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[18__840 .GSR = "DISABLED";
    FD1S3AX \registers_13[[17__841  (.D(\registers[13] [21]), .CK(clk_c), 
            .Q(\registers[13] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[17__841 .GSR = "DISABLED";
    FD1S3AX \registers_13[[16__842  (.D(\registers[13] [20]), .CK(clk_c), 
            .Q(\registers[13] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[16__842 .GSR = "DISABLED";
    FD1S3AX \registers_13[[15__843  (.D(\registers[13] [19]), .CK(clk_c), 
            .Q(\registers[13] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[15__843 .GSR = "DISABLED";
    FD1S3AX \registers_13[[14__844  (.D(\registers[13] [18]), .CK(clk_c), 
            .Q(\registers[13] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[14__844 .GSR = "DISABLED";
    FD1S3AX \registers_13[[13__845  (.D(\registers[13] [17]), .CK(clk_c), 
            .Q(\registers[13] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[13__845 .GSR = "DISABLED";
    FD1S3AX \registers_13[[12__846  (.D(\registers[13] [16]), .CK(clk_c), 
            .Q(\registers[13] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[12__846 .GSR = "DISABLED";
    FD1S3AX \registers_13[[11__847  (.D(\registers[13] [15]), .CK(clk_c), 
            .Q(\registers[13] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[11__847 .GSR = "DISABLED";
    FD1S3AX \registers_13[[10__848  (.D(\registers[13] [14]), .CK(clk_c), 
            .Q(\registers[13] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[10__848 .GSR = "DISABLED";
    FD1S3AX \registers_13[[9__849  (.D(\registers[13] [13]), .CK(clk_c), 
            .Q(\registers[13] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[9__849 .GSR = "DISABLED";
    FD1S3AX \registers_13[[8__850  (.D(\registers[13] [12]), .CK(clk_c), 
            .Q(\registers[13] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[8__850 .GSR = "DISABLED";
    FD1S3AX \registers_13[[7__851  (.D(\registers[13] [11]), .CK(clk_c), 
            .Q(\registers[13] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[7__851 .GSR = "DISABLED";
    FD1S3AX \registers_13[[6__852  (.D(\registers[13] [10]), .CK(clk_c), 
            .Q(\registers[13] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[6__852 .GSR = "DISABLED";
    FD1S3AX \registers_13[[5__853  (.D(\registers[13] [9]), .CK(clk_c), 
            .Q(\registers[13] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[5__853 .GSR = "DISABLED";
    FD1S3AX \registers_13[[4__854  (.D(\registers[13] [8]), .CK(clk_c), 
            .Q(\registers[13] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[4__854 .GSR = "DISABLED";
    FD1S3AX \registers_14[[3__855  (.D(registers_14__3__N_1819), .CK(clk_c), 
            .Q(\registers[14] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[3__855 .GSR = "DISABLED";
    FD1S3AX \registers_14[[2__856  (.D(registers_14__2__N_1822), .CK(clk_c), 
            .Q(\registers[14] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[2__856 .GSR = "DISABLED";
    FD1S3AX \registers_14[[1__857  (.D(registers_14__1__N_1823), .CK(clk_c), 
            .Q(\registers[14] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[1__857 .GSR = "DISABLED";
    FD1S3AX \registers_14[[0__858  (.D(registers_14__0__N_1824), .CK(clk_c), 
            .Q(\registers[14] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[0__858 .GSR = "DISABLED";
    FD1S3AX \registers_14[[31__859  (.D(\registers[14] [3]), .CK(clk_c), 
            .Q(\registers[14] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[31__859 .GSR = "DISABLED";
    FD1S3AX \registers_14[[30__860  (.D(\registers[14] [2]), .CK(clk_c), 
            .Q(\registers[14] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[30__860 .GSR = "DISABLED";
    FD1S3AX \registers_14[[29__861  (.D(\registers[14] [1]), .CK(clk_c), 
            .Q(\registers[14] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[29__861 .GSR = "DISABLED";
    FD1S3AX \registers_14[[28__862  (.D(\registers[14] [0]), .CK(clk_c), 
            .Q(\registers[14] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[28__862 .GSR = "DISABLED";
    FD1S3AX \registers_14[[27__863  (.D(\registers[14] [31]), .CK(clk_c), 
            .Q(\registers[14] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[27__863 .GSR = "DISABLED";
    FD1S3AX \registers_14[[26__864  (.D(\registers[14] [30]), .CK(clk_c), 
            .Q(\registers[14] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[26__864 .GSR = "DISABLED";
    FD1S3AX \registers_14[[25__865  (.D(\registers[14] [29]), .CK(clk_c), 
            .Q(\registers[14] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[25__865 .GSR = "DISABLED";
    FD1S3AX \registers_14[[24__866  (.D(\registers[14] [28]), .CK(clk_c), 
            .Q(\registers[14] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[24__866 .GSR = "DISABLED";
    FD1S3AX \registers_14[[23__867  (.D(\registers[14] [27]), .CK(clk_c), 
            .Q(\registers[14] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[23__867 .GSR = "DISABLED";
    FD1S3AX \registers_14[[22__868  (.D(\registers[14] [26]), .CK(clk_c), 
            .Q(\registers[14] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[22__868 .GSR = "DISABLED";
    FD1S3AX \registers_14[[21__869  (.D(\registers[14] [25]), .CK(clk_c), 
            .Q(\registers[14] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[21__869 .GSR = "DISABLED";
    FD1S3AX \registers_14[[20__870  (.D(\registers[14] [24]), .CK(clk_c), 
            .Q(\registers[14] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[20__870 .GSR = "DISABLED";
    FD1S3AX \registers_14[[19__871  (.D(\registers[14] [23]), .CK(clk_c), 
            .Q(\registers[14] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[19__871 .GSR = "DISABLED";
    FD1S3AX \registers_14[[18__872  (.D(\registers[14] [22]), .CK(clk_c), 
            .Q(\registers[14] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[18__872 .GSR = "DISABLED";
    FD1S3AX \registers_14[[17__873  (.D(\registers[14] [21]), .CK(clk_c), 
            .Q(\registers[14] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[17__873 .GSR = "DISABLED";
    FD1S3AX \registers_14[[16__874  (.D(\registers[14] [20]), .CK(clk_c), 
            .Q(\registers[14] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[16__874 .GSR = "DISABLED";
    FD1S3AX \registers_14[[15__875  (.D(\registers[14] [19]), .CK(clk_c), 
            .Q(\registers[14] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[15__875 .GSR = "DISABLED";
    FD1S3AX \registers_14[[14__876  (.D(\registers[14] [18]), .CK(clk_c), 
            .Q(\registers[14] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[14__876 .GSR = "DISABLED";
    FD1S3AX \registers_14[[13__877  (.D(\registers[14] [17]), .CK(clk_c), 
            .Q(\registers[14] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[13__877 .GSR = "DISABLED";
    FD1S3AX \registers_14[[12__878  (.D(\registers[14] [16]), .CK(clk_c), 
            .Q(\registers[14] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[12__878 .GSR = "DISABLED";
    FD1S3AX \registers_14[[11__879  (.D(\registers[14] [15]), .CK(clk_c), 
            .Q(\registers[14] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[11__879 .GSR = "DISABLED";
    FD1S3AX \registers_14[[10__880  (.D(\registers[14] [14]), .CK(clk_c), 
            .Q(\registers[14] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[10__880 .GSR = "DISABLED";
    FD1S3AX \registers_14[[9__881  (.D(\registers[14] [13]), .CK(clk_c), 
            .Q(\registers[14] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[9__881 .GSR = "DISABLED";
    FD1S3AX \registers_14[[8__882  (.D(\registers[14] [12]), .CK(clk_c), 
            .Q(\registers[14] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[8__882 .GSR = "DISABLED";
    FD1S3AX \registers_14[[7__883  (.D(\registers[14] [11]), .CK(clk_c), 
            .Q(\registers[14] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[7__883 .GSR = "DISABLED";
    FD1S3AX \registers_14[[6__884  (.D(\registers[14] [10]), .CK(clk_c), 
            .Q(\registers[14] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[6__884 .GSR = "DISABLED";
    FD1S3AX \registers_14[[5__885  (.D(\registers[14] [9]), .CK(clk_c), 
            .Q(\registers[14] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[5__885 .GSR = "DISABLED";
    FD1S3AX \registers_14[[4__886  (.D(\registers[14] [8]), .CK(clk_c), 
            .Q(\registers[14] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[4__886 .GSR = "DISABLED";
    FD1S3AX \registers_15[[3__887  (.D(registers_15__3__N_1825), .CK(clk_c), 
            .Q(\registers[15] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[3__887 .GSR = "DISABLED";
    FD1S3AX \registers_15[[2__888  (.D(registers_15__2__N_1828), .CK(clk_c), 
            .Q(\registers[15] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[2__888 .GSR = "DISABLED";
    FD1S3AX \registers_15[[1__889  (.D(registers_15__1__N_1829), .CK(clk_c), 
            .Q(\registers[15] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[1__889 .GSR = "DISABLED";
    FD1S3AX \registers_15[[0__890  (.D(registers_15__0__N_1830), .CK(clk_c), 
            .Q(\registers[15] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[0__890 .GSR = "DISABLED";
    FD1S3AX \registers_15[[31__891  (.D(\registers[15] [3]), .CK(clk_c), 
            .Q(\registers[15] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[31__891 .GSR = "DISABLED";
    FD1S3AX \registers_15[[30__892  (.D(\registers[15] [2]), .CK(clk_c), 
            .Q(\registers[15] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[30__892 .GSR = "DISABLED";
    FD1S3AX \registers_15[[29__893  (.D(\registers[15] [1]), .CK(clk_c), 
            .Q(\registers[15] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[29__893 .GSR = "DISABLED";
    FD1S3AX \registers_15[[28__894  (.D(\registers[15] [0]), .CK(clk_c), 
            .Q(\registers[15] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[28__894 .GSR = "DISABLED";
    FD1S3AX \registers_15[[27__895  (.D(\registers[15] [31]), .CK(clk_c), 
            .Q(\registers[15] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[27__895 .GSR = "DISABLED";
    FD1S3AX \registers_15[[26__896  (.D(\registers[15] [30]), .CK(clk_c), 
            .Q(\registers[15] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[26__896 .GSR = "DISABLED";
    FD1S3AX \registers_15[[25__897  (.D(\registers[15] [29]), .CK(clk_c), 
            .Q(\registers[15] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[25__897 .GSR = "DISABLED";
    FD1S3AX \registers_15[[24__898  (.D(\registers[15] [28]), .CK(clk_c), 
            .Q(\registers[15] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[24__898 .GSR = "DISABLED";
    FD1S3AX \registers_15[[23__899  (.D(\registers[15] [27]), .CK(clk_c), 
            .Q(\registers[15] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[23__899 .GSR = "DISABLED";
    FD1S3AX \registers_15[[22__900  (.D(\registers[15] [26]), .CK(clk_c), 
            .Q(\registers[15] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[22__900 .GSR = "DISABLED";
    FD1S3AX \registers_15[[21__901  (.D(\registers[15] [25]), .CK(clk_c), 
            .Q(\registers[15] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[21__901 .GSR = "DISABLED";
    FD1S3AX \registers_15[[20__902  (.D(\registers[15] [24]), .CK(clk_c), 
            .Q(\registers[15] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[20__902 .GSR = "DISABLED";
    FD1S3AX \registers_15[[19__903  (.D(\registers[15] [23]), .CK(clk_c), 
            .Q(\registers[15] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[19__903 .GSR = "DISABLED";
    FD1S3AX \registers_15[[18__904  (.D(\registers[15] [22]), .CK(clk_c), 
            .Q(\registers[15] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[18__904 .GSR = "DISABLED";
    FD1S3AX \registers_15[[17__905  (.D(\registers[15] [21]), .CK(clk_c), 
            .Q(\registers[15] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[17__905 .GSR = "DISABLED";
    FD1S3AX \registers_15[[16__906  (.D(\registers[15] [20]), .CK(clk_c), 
            .Q(\registers[15] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[16__906 .GSR = "DISABLED";
    FD1S3AX \registers_15[[15__907  (.D(\registers[15] [19]), .CK(clk_c), 
            .Q(\registers[15] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[15__907 .GSR = "DISABLED";
    FD1S3AX \registers_15[[14__908  (.D(\registers[15] [18]), .CK(clk_c), 
            .Q(\registers[15] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[14__908 .GSR = "DISABLED";
    FD1S3AX \registers_15[[13__909  (.D(\registers[15] [17]), .CK(clk_c), 
            .Q(\registers[15] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[13__909 .GSR = "DISABLED";
    FD1S3AX \registers_15[[12__910  (.D(\registers[15] [16]), .CK(clk_c), 
            .Q(\registers[15] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[12__910 .GSR = "DISABLED";
    FD1S3AX \registers_15[[11__911  (.D(\registers[15] [15]), .CK(clk_c), 
            .Q(\registers[15] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[11__911 .GSR = "DISABLED";
    FD1S3AX \registers_15[[10__912  (.D(\registers[15] [14]), .CK(clk_c), 
            .Q(\registers[15] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[10__912 .GSR = "DISABLED";
    FD1S3AX \registers_15[[9__913  (.D(\registers[15] [13]), .CK(clk_c), 
            .Q(\registers[15] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[9__913 .GSR = "DISABLED";
    FD1S3AX \registers_15[[8__914  (.D(\registers[15] [12]), .CK(clk_c), 
            .Q(\registers[15] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[8__914 .GSR = "DISABLED";
    FD1S3AX \registers_15[[7__915  (.D(\registers[15] [11]), .CK(clk_c), 
            .Q(\registers[15] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[7__915 .GSR = "DISABLED";
    FD1S3AX \registers_15[[6__916  (.D(\registers[15] [10]), .CK(clk_c), 
            .Q(\registers[15] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[6__916 .GSR = "DISABLED";
    FD1S3AX \registers_15[[5__917  (.D(\registers[15] [9]), .CK(clk_c), 
            .Q(\registers[15] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[5__917 .GSR = "DISABLED";
    FD1S3AX \registers_15[[4__918  (.D(\registers[15] [8]), .CK(clk_c), 
            .Q(\registers[15] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[4__918 .GSR = "DISABLED";
    FD1S3AX \registers_1[[3__503  (.D(registers_1__3__N_1753), .CK(clk_c), 
            .Q(\registers[1] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[3__503 .GSR = "DISABLED";
    L6MUX21 i27670 (.D0(n30375), .D1(n30376), .SD(rs1[2]), .Z(n30379));
    L6MUX21 i27685 (.D0(n30390), .D1(n30391), .SD(rs2[2]), .Z(n30394));
    PFUMX i27721 (.BLUT(n30426), .ALUT(n30427), .C0(rs1[2]), .Z(n30430));
    PFUMX i27728 (.BLUT(n30433), .ALUT(n30434), .C0(rs2[2]), .Z(n30437));
    PFUMX i27585 (.BLUT(n30286), .ALUT(n30287), .C0(rs2[1]), .Z(n30294));
    PFUMX i27600 (.BLUT(n30301), .ALUT(n30302), .C0(rs1[1]), .Z(n30309));
    LUT4 i27659_3_lut (.A(\registers[2] [6]), .B(\reg_access[3][2] ), .C(rs1[0]), 
         .Z(n30368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27659_3_lut.init = 16'hcaca;
    LUT4 i27658_3_lut (.A(\registers[1] [6]), .B(rs1[0]), .Z(n30367)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27658_3_lut.init = 16'h8888;
    LUT4 i27599_3_lut (.A(\registers[14] [4]), .B(\registers[15] [4]), .C(rs1[0]), 
         .Z(n30308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27599_3_lut.init = 16'hcaca;
    LUT4 i27598_3_lut (.A(\registers[12] [4]), .B(\registers[13] [4]), .C(rs1[0]), 
         .Z(n30307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27598_3_lut.init = 16'hcaca;
    LUT4 i27597_3_lut (.A(\registers[10] [4]), .B(\registers[11] [4]), .C(rs1[0]), 
         .Z(n30306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27597_3_lut.init = 16'hcaca;
    LUT4 i27596_3_lut (.A(\registers[8] [4]), .B(\registers[9] [4]), .C(rs1[0]), 
         .Z(n30305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27596_3_lut.init = 16'hcaca;
    LUT4 i27738_4_lut_4_lut (.A(\registers[2] [5]), .B(rs1[0]), .C(rs1[1]), 
         .D(\registers[1] [5]), .Z(n30447)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i27738_4_lut_4_lut.init = 16'h2c20;
    LUT4 i27731_4_lut_4_lut (.A(\registers[2] [5]), .B(rs2[0]), .C(rs2[1]), 
         .D(\registers[1] [5]), .Z(n30440)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i27731_4_lut_4_lut.init = 16'h2c20;
    LUT4 i27595_3_lut (.A(\registers[6] [4]), .B(\registers[7] [4]), .C(rs1[0]), 
         .Z(n30304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27595_3_lut.init = 16'hcaca;
    LUT4 i27594_3_lut (.A(\registers[5] [4]), .B(rs1[0]), .Z(n30303)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27594_3_lut.init = 16'h8888;
    LUT4 i27606_3_lut (.A(n30313), .B(n30314), .C(rs1[3]), .Z(data_rs1[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27606_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(n32676), .B(data_rs1[1]), .C(n57), .D(\mie[13] ), 
         .Z(n927)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_293 (.A(n32676), .B(data_rs1[1]), .C(n57), 
         .D(\mie[9] ), .Z(n894)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_293.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_294 (.A(n32676), .B(data_rs1[1]), .C(n57), 
         .D(\mie[5] ), .Z(n861)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_294.init = 16'hf888;
    LUT4 i1_3_lut_4_lut_adj_295 (.A(n32676), .B(data_rs1[1]), .C(n57), 
         .D(\mie[1] ), .Z(n794)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_295.init = 16'hf888;
    LUT4 i27584_3_lut (.A(\registers[14] [4]), .B(\registers[15] [4]), .C(rs2[0]), 
         .Z(n30293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27584_3_lut.init = 16'hcaca;
    LUT4 i27583_3_lut (.A(\registers[12] [4]), .B(\registers[13] [4]), .C(rs2[0]), 
         .Z(n30292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27583_3_lut.init = 16'hcaca;
    LUT4 i27582_3_lut (.A(\registers[10] [4]), .B(\registers[11] [4]), .C(rs2[0]), 
         .Z(n30291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27582_3_lut.init = 16'hcaca;
    LUT4 i27581_3_lut (.A(\registers[8] [4]), .B(\registers[9] [4]), .C(rs2[0]), 
         .Z(n30290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27581_3_lut.init = 16'hcaca;
    LUT4 i27580_3_lut (.A(\registers[6] [4]), .B(\registers[7] [4]), .C(rs2[0]), 
         .Z(n30289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27580_3_lut.init = 16'hcaca;
    LUT4 i27579_3_lut (.A(\registers[5] [4]), .B(rs2[0]), .Z(n30288)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27579_3_lut.init = 16'h8888;
    L6MUX21 i27590 (.D0(n30296), .D1(n30297), .SD(rs2[2]), .Z(n30299));
    L6MUX21 i27605 (.D0(n30311), .D1(n30312), .SD(rs1[2]), .Z(n30314));
    LUT4 i27724_4_lut_4_lut (.A(\registers[2] [7]), .B(rs2[0]), .C(rs2[1]), 
         .D(\registers[1] [7]), .Z(n30433)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i27724_4_lut_4_lut.init = 16'h2c20;
    L6MUX21 i27671 (.D0(n30377), .D1(n30378), .SD(rs1[2]), .Z(n30380));
    L6MUX21 i27686 (.D0(n30392), .D1(n30393), .SD(rs2[2]), .Z(n30395));
    L6MUX21 i27722 (.D0(n30428), .D1(n30429), .SD(rs1[2]), .Z(n30431));
    L6MUX21 i27729 (.D0(n30435), .D1(n30436), .SD(rs2[2]), .Z(n30438));
    PFUMX i27735 (.BLUT(n30440), .ALUT(n30441), .C0(rs2[2]), .Z(n30444));
    L6MUX21 i27736 (.D0(n30442), .D1(n30443), .SD(rs2[2]), .Z(n30445));
    PFUMX i27742 (.BLUT(n30447), .ALUT(n30448), .C0(rs1[2]), .Z(n30451));
    L6MUX21 i27743 (.D0(n30449), .D1(n30450), .SD(rs1[2]), .Z(n30452));
    LUT4 i1_3_lut_4_lut_adj_296 (.A(n32676), .B(data_rs1[0]), .C(n29683), 
         .D(\mie[12] ), .Z(n928)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_296.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_297 (.A(n32676), .B(data_rs1[0]), .C(n29683), 
         .D(\mie[8] ), .Z(n895)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_297.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_298 (.A(n32676), .B(data_rs1[0]), .C(n29683), 
         .D(\mie[4] ), .Z(n862)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_298.init = 16'h8f88;
    LUT4 i27821_3_lut_4_lut (.A(\registers[5] [5]), .B(rs2[0]), .C(rs2[1]), 
         .D(n5_adj_3134), .Z(n30441)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i27821_3_lut_4_lut.init = 16'hf808;
    LUT4 i27818_3_lut_4_lut (.A(\registers[5] [5]), .B(rs1[0]), .C(rs1[1]), 
         .D(n5), .Z(n30448)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i27818_3_lut_4_lut.init = 16'hf808;
    LUT4 i27723_3_lut (.A(n30430), .B(n30431), .C(rs1[3]), .Z(data_rs1[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27723_3_lut.init = 16'hcaca;
    PFUMX i27586 (.BLUT(n30288), .ALUT(n30289), .C0(rs2[1]), .Z(n30295));
    PFUMX i27587 (.BLUT(n30290), .ALUT(n30291), .C0(rs2[1]), .Z(n30296));
    PFUMX i27588 (.BLUT(n30292), .ALUT(n30293), .C0(rs2[1]), .Z(n30297));
    LUT4 i27744_3_lut (.A(n30451), .B(n30452), .C(rs1[3]), .Z(data_rs1[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27744_3_lut.init = 16'hcaca;
    LUT4 i27737_3_lut (.A(n30444), .B(n30445), .C(rs2[3]), .Z(data_rs2[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27737_3_lut.init = 16'hcaca;
    LUT4 i27730_3_lut (.A(n30437), .B(n30438), .C(rs2[3]), .Z(data_rs2[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27730_3_lut.init = 16'hcaca;
    PFUMX i27601 (.BLUT(n30303), .ALUT(n30304), .C0(rs1[1]), .Z(n30310));
    LUT4 i28351_3_lut (.A(n34281), .B(n34283), .C(\counter_hi[2] ), .Z(\reg_access[4][3] )) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(40[41:55])
    defparam i28351_3_lut.init = 16'h0808;
    LUT4 i28354_3_lut (.A(\counter_hi[2] ), .B(n34283), .C(n34281), .Z(\reg_access[3][2] )) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(38[47:61])
    defparam i28354_3_lut.init = 16'h0404;
    PFUMX i27602 (.BLUT(n30305), .ALUT(n30306), .C0(rs1[1]), .Z(n30311));
    PFUMX i27603 (.BLUT(n30307), .ALUT(n30308), .C0(rs1[1]), .Z(n30312));
    LUT4 i27593_3_lut (.A(\registers[2] [4]), .B(\reg_access[4][3] ), .C(rs1[0]), 
         .Z(n30302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27593_3_lut.init = 16'hcaca;
    LUT4 i27592_3_lut (.A(\registers[1] [4]), .B(rs1[0]), .Z(n30301)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27592_3_lut.init = 16'h8888;
    LUT4 i27578_3_lut (.A(\registers[2] [4]), .B(\reg_access[4][3] ), .C(rs2[0]), 
         .Z(n30287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27578_3_lut.init = 16'hcaca;
    LUT4 i27577_3_lut (.A(\registers[1] [4]), .B(rs2[0]), .Z(n30286)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27577_3_lut.init = 16'h8888;
    LUT4 i21404_3_lut (.A(\mie[5] ), .B(\mie[13] ), .C(\counter_hi[3] ), 
         .Z(n4829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(139[15:25])
    defparam i21404_3_lut.init = 16'hcaca;
    PFUMX i27666 (.BLUT(n30367), .ALUT(n30368), .C0(rs1[1]), .Z(n30375));
    LUT4 i27606_3_lut_rep_852 (.A(n30313), .B(n30314), .C(rs1[3]), .Z(n34292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27606_3_lut_rep_852.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i5_3_lut (.A(\registers[6] [7]), .B(\registers[7] [7]), 
         .C(rs2[0]), .Z(n5_adj_3143)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i4_3_lut (.A(\reg_access[4][3] ), .B(\registers[5] [7]), 
         .C(rs2[0]), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i4_3_lut.init = 16'hcaca;
    LUT4 i27889_3_lut (.A(n4), .B(n5_adj_3143), .C(rs2[1]), .Z(n30434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27889_3_lut.init = 16'hcaca;
    PFUMX i27667 (.BLUT(n30369), .ALUT(n30370), .C0(rs1[1]), .Z(n30376));
    PFUMX i27668 (.BLUT(n30371), .ALUT(n30372), .C0(rs1[1]), .Z(n30377));
    PFUMX i27669 (.BLUT(n30373), .ALUT(n30374), .C0(rs1[1]), .Z(n30378));
    LUT4 rs1_3__I_0_Mux_3_i5_3_lut (.A(\registers[6] [7]), .B(\registers[7] [7]), 
         .C(rs1[0]), .Z(n5_adj_3144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i4_3_lut (.A(\reg_access[4][3] ), .B(\registers[5] [7]), 
         .C(rs1[0]), .Z(n4_adj_3145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i4_3_lut.init = 16'hcaca;
    LUT4 i27891_3_lut (.A(n4_adj_3145), .B(n5_adj_3144), .C(rs1[1]), .Z(n30427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27891_3_lut.init = 16'hcaca;
    PFUMX i27682 (.BLUT(n30384), .ALUT(n30385), .C0(rs2[1]), .Z(n30391));
    PFUMX i27683 (.BLUT(n30386), .ALUT(n30387), .C0(rs2[1]), .Z(n30392));
    PFUMX i27681 (.BLUT(n30382), .ALUT(n30383), .C0(rs2[1]), .Z(n30390));
    PFUMX i27684 (.BLUT(n30388), .ALUT(n30389), .C0(rs2[1]), .Z(n30393));
    PFUMX i27719 (.BLUT(n8_adj_3142), .ALUT(n9_adj_3141), .C0(rs1[1]), 
          .Z(n30428));
    PFUMX i27720 (.BLUT(n11_adj_3140), .ALUT(n12_adj_3139), .C0(rs1[1]), 
          .Z(n30429));
    PFUMX i27726 (.BLUT(n8_adj_3138), .ALUT(n9_adj_3137), .C0(rs2[1]), 
          .Z(n30435));
    PFUMX i27727 (.BLUT(n11_adj_3136), .ALUT(n12_adj_3135), .C0(rs2[1]), 
          .Z(n30436));
    PFUMX i27733 (.BLUT(n8_adj_3133), .ALUT(n9_adj_3132), .C0(rs2[1]), 
          .Z(n30442));
    PFUMX i27734 (.BLUT(n11_adj_3131), .ALUT(n12_adj_3130), .C0(rs2[1]), 
          .Z(n30443));
    PFUMX i27740 (.BLUT(n8), .ALUT(n9), .C0(rs1[1]), .Z(n30449));
    PFUMX i27741 (.BLUT(n11), .ALUT(n12), .C0(rs1[1]), .Z(n30450));
    
endmodule
//
// Verilog Description of module tinyqv_counter_U0
//

module tinyqv_counter_U0 (cy, clk_c, n32840, \increment_result_3__N_1925[0] , 
            instrret_count, n32665, n32683) /* synthesis syn_module_defined=1 */ ;
    output cy;
    input clk_c;
    input n32840;
    input \increment_result_3__N_1925[0] ;
    output [3:0]instrret_count;
    input n32665;
    input n32683;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [4:0]increment_result_3__N_1925;
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    
    FD1S3IX cy_51 (.D(increment_result_3__N_1925[4]), .CK(clk_c), .CD(n32840), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3IX register_2__48 (.D(increment_result_3__N_1925[2]), .CK(clk_c), 
            .CD(n32840), .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result_3__N_1925[1]), .CK(clk_c), 
            .CD(n32840), .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(\increment_result_3__N_1925[0] ), .CK(clk_c), 
            .CD(n32840), .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(register[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(register[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(register[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(instrret_count[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(register[10]), .CK(clk_c), .Q(instrret_count[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(register[9]), .CK(clk_c), .Q(instrret_count[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(register[8]), .CK(clk_c), .Q(instrret_count[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result_3__N_1925[3]), .CK(clk_c), 
            .CD(n32840), .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 i4775_2_lut_3_lut_4_lut (.A(instrret_count[1]), .B(n32665), .C(instrret_count[3]), 
         .D(instrret_count[2]), .Z(increment_result_3__N_1925[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4775_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4777_2_lut_3_lut_4_lut (.A(instrret_count[1]), .B(n32665), .C(instrret_count[3]), 
         .D(instrret_count[2]), .Z(increment_result_3__N_1925[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4777_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4761_2_lut_3_lut (.A(instrret_count[0]), .B(n32683), .C(instrret_count[1]), 
         .Z(increment_result_3__N_1925[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4761_2_lut_3_lut.init = 16'h7878;
    LUT4 i4768_2_lut_3_lut_4_lut (.A(instrret_count[0]), .B(n32683), .C(instrret_count[2]), 
         .D(instrret_count[1]), .Z(increment_result_3__N_1925[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4768_2_lut_3_lut_4_lut.init = 16'h78f0;
    
endmodule
//
// Verilog Description of module \tinyqv_counter(OUTPUT_WIDTH=7) 
//

module \tinyqv_counter(OUTPUT_WIDTH=7)  (cy, clk_c, n32840, \increment_result_3__N_1911[0] , 
            cycle_count_wide, n32701, n32731, n32652, n32765) /* synthesis syn_module_defined=1 */ ;
    output cy;
    input clk_c;
    input n32840;
    input \increment_result_3__N_1911[0] ;
    output [6:0]cycle_count_wide;
    input n32701;
    input n32731;
    output n32652;
    input n32765;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [4:0]increment_result_3__N_1911;
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    
    FD1S3IX cy_51 (.D(increment_result_3__N_1911[4]), .CK(clk_c), .CD(n32840), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3IX register_2__48 (.D(increment_result_3__N_1911[2]), .CK(clk_c), 
            .CD(n32840), .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result_3__N_1911[1]), .CK(clk_c), 
            .CD(n32840), .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(\increment_result_3__N_1911[0] ), .CK(clk_c), 
            .CD(n32840), .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(cycle_count_wide[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(cycle_count_wide[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(cycle_count_wide[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(cycle_count_wide[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(cycle_count_wide[6]), .CK(clk_c), .Q(cycle_count_wide[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(cycle_count_wide[5]), .CK(clk_c), .Q(cycle_count_wide[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(cycle_count_wide[4]), .CK(clk_c), .Q(cycle_count_wide[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result_3__N_1911[3]), .CK(clk_c), 
            .CD(n32840), .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 i4749_2_lut_3_lut_4_lut (.A(cycle_count_wide[1]), .B(n32701), .C(cycle_count_wide[3]), 
         .D(cycle_count_wide[2]), .Z(increment_result_3__N_1911[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4749_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4747_2_lut_3_lut_4_lut (.A(cycle_count_wide[1]), .B(n32701), .C(cycle_count_wide[3]), 
         .D(cycle_count_wide[2]), .Z(increment_result_3__N_1911[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4747_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4742_2_lut_rep_637_3_lut_4_lut (.A(cycle_count_wide[0]), .B(n32731), 
         .C(cycle_count_wide[2]), .D(cycle_count_wide[1]), .Z(n32652)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4742_2_lut_rep_637_3_lut_4_lut.init = 16'h8000;
    LUT4 i4740_2_lut_3_lut_4_lut (.A(cycle_count_wide[0]), .B(n32731), .C(cycle_count_wide[2]), 
         .D(cycle_count_wide[1]), .Z(increment_result_3__N_1911[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4740_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4733_2_lut_3_lut_4_lut (.A(cy), .B(n32765), .C(cycle_count_wide[1]), 
         .D(cycle_count_wide[0]), .Z(increment_result_3__N_1911[1])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[93:118])
    defparam i4733_2_lut_3_lut_4_lut.init = 16'h4bf0;
    
endmodule
//
// Verilog Description of module tinyqv_alu
//

module tinyqv_alu (alu_a_in, n32625, n29121, alu_b_in, \alu_op_in[2] , 
            n32748, n32688, n32592, n32646, n32626, cy_out, n28225, 
            n31758, n32738, n31760, n32624, n32749, alu_out, n4901) /* synthesis syn_module_defined=1 */ ;
    input [3:0]alu_a_in;
    input n32625;
    input n29121;
    input [3:0]alu_b_in;
    input \alu_op_in[2] ;
    input n32748;
    input n32688;
    input n32592;
    input n32646;
    input n32626;
    output cy_out;
    input n28225;
    output n31758;
    input n32738;
    output n31760;
    input n32624;
    input n32749;
    output [3:0]alu_out;
    input [3:0]n4901;
    
    
    wire n34274, n32562, n6, n29598, n29055, n32662, n32574;
    wire [3:0]n4911;
    wire [3:0]a_xor_b;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[16:23])
    
    wire n32591, n29037, n32558, n28989, n32557, n34273, cmp_res_N_1855, 
        n31759;
    wire [3:0]n4920;
    
    LUT4 i4717_2_lut_3_lut_4_lut_4_lut (.A(alu_a_in[2]), .B(n34274), .C(n32562), 
         .D(n32625), .Z(n6)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4717_2_lut_3_lut_4_lut_4_lut.init = 16'hfea8;
    LUT4 i26958_4_lut (.A(alu_a_in[0]), .B(n29121), .C(alu_b_in[0]), .D(\alu_op_in[2] ), 
         .Z(n29598)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam i26958_4_lut.init = 16'h5a66;
    LUT4 mux_3030_i2_4_lut (.A(n29055), .B(n32662), .C(\alu_op_in[2] ), 
         .D(n32574), .Z(n4911[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_3030_i2_4_lut.init = 16'hc5ca;
    LUT4 a_3__I_0_29_i3_2_lut (.A(alu_a_in[2]), .B(alu_b_in[2]), .Z(a_xor_b[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i3_2_lut.init = 16'h6666;
    LUT4 a_3__I_0_29_i4_2_lut (.A(alu_a_in[3]), .B(alu_b_in[3]), .Z(a_xor_b[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i4_2_lut.init = 16'h6666;
    LUT4 a_3__I_0_29_i1_2_lut (.A(alu_a_in[0]), .B(alu_b_in[0]), .Z(a_xor_b[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i1_2_lut.init = 16'h6666;
    LUT4 i5464_3_lut_rep_576_4_lut (.A(alu_b_in[0]), .B(n32748), .C(n32688), 
         .D(alu_a_in[0]), .Z(n32591)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i5464_3_lut_rep_576_4_lut.init = 16'hf600;
    LUT4 i5459_4_lut_rep_842 (.A(alu_a_in[1]), .B(n32592), .C(n32591), 
         .D(n32646), .Z(n34274)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i5459_4_lut_rep_842.init = 16'haaa8;
    LUT4 i4703_2_lut_rep_559_4_lut_3_lut_4_lut (.A(alu_b_in[0]), .B(n32748), 
         .C(alu_a_in[0]), .D(n32688), .Z(n32574)) /* synthesis lut_function=(A (B (C (D))+!B (C+(D)))+!A (B (C+(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i4703_2_lut_rep_559_4_lut_3_lut_4_lut.init = 16'hf660;
    LUT4 i1_2_lut_3_lut (.A(alu_b_in[2]), .B(n32748), .C(alu_a_in[2]), 
         .Z(n29037)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut.init = 16'h9696;
    LUT4 mux_3030_i3_4_lut (.A(n29037), .B(a_xor_b[2]), .C(\alu_op_in[2] ), 
         .D(n32558), .Z(n4911[2])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_3030_i3_4_lut.init = 16'hc5ca;
    LUT4 i1_2_lut_3_lut_adj_291 (.A(alu_b_in[3]), .B(n32748), .C(alu_a_in[3]), 
         .Z(n28989)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut_adj_291.init = 16'h9696;
    LUT4 i4724_4_lut_4_lut (.A(alu_a_in[3]), .B(n32557), .C(n34273), .D(n32626), 
         .Z(cy_out)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4724_4_lut_4_lut.init = 16'hfea8;
    LUT4 i4710_2_lut_rep_543_3_lut_4_lut_4_lut (.A(alu_a_in[1]), .B(n32592), 
         .C(n32591), .D(n32646), .Z(n32558)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4710_2_lut_rep_543_3_lut_4_lut_4_lut.init = 16'hfea8;
    LUT4 mux_3030_i4_4_lut (.A(n28989), .B(a_xor_b[3]), .C(\alu_op_in[2] ), 
         .D(n6), .Z(n4911[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_3030_i4_4_lut.init = 16'hc5ca;
    LUT4 i1_4_lut (.A(a_xor_b[2]), .B(a_xor_b[3]), .C(a_xor_b[0]), .D(n28225), 
         .Z(cmp_res_N_1855)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    LUT4 i4715_2_lut_rep_542_3_lut_4_lut (.A(n32646), .B(n32574), .C(n32625), 
         .D(n34274), .Z(n32557)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4715_2_lut_rep_542_3_lut_4_lut.init = 16'hf080;
    LUT4 i1_2_lut_3_lut_adj_292 (.A(alu_b_in[1]), .B(n32748), .C(alu_a_in[1]), 
         .Z(n29055)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut_adj_292.init = 16'h9696;
    LUT4 n6997_bdd_4_lut (.A(n32557), .B(n34273), .C(n32626), .D(alu_a_in[3]), 
         .Z(n31759)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+(D)))) */ ;
    defparam n6997_bdd_4_lut.init = 16'hf110;
    LUT4 alu_op_in_0__bdd_4_lut (.A(n32557), .B(n34273), .C(n32626), .D(alu_a_in[3]), 
         .Z(n31758)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C (D))))) */ ;
    defparam alu_op_in_0__bdd_4_lut.init = 16'h011f;
    LUT4 a_3__I_0_29_i2_2_lut_rep_647 (.A(alu_a_in[1]), .B(alu_b_in[1]), 
         .Z(n32662)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i2_2_lut_rep_647.init = 16'h6666;
    PFUMX i28887 (.BLUT(cmp_res_N_1855), .ALUT(n31759), .C0(n32738), .Z(n31760));
    LUT4 i4708_2_lut_rep_547_3_lut_4_lut (.A(n32624), .B(n32688), .C(n32646), 
         .D(n32591), .Z(n32562)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4708_2_lut_rep_547_3_lut_4_lut.init = 16'hf080;
    LUT4 i15202_2_lut_4_lut (.A(n32749), .B(\alu_op_in[2] ), .C(n32738), 
         .D(n4920[1]), .Z(alu_out[1])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i15202_2_lut_4_lut.init = 16'hc500;
    LUT4 i14910_2_lut_4_lut (.A(n32749), .B(\alu_op_in[2] ), .C(n32738), 
         .D(n4920[0]), .Z(alu_out[0])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i14910_2_lut_4_lut.init = 16'hc500;
    LUT4 i15200_2_lut_4_lut (.A(n32749), .B(\alu_op_in[2] ), .C(n32738), 
         .D(n4920[3]), .Z(alu_out[3])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i15200_2_lut_4_lut.init = 16'hc500;
    LUT4 i15201_2_lut_4_lut (.A(n32749), .B(\alu_op_in[2] ), .C(n32738), 
         .D(n4920[2]), .Z(alu_out[2])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i15201_2_lut_4_lut.init = 16'hc500;
    PFUMX mux_3035_i4 (.BLUT(n4911[3]), .ALUT(n4901[3]), .C0(n32738), 
          .Z(n4920[3]));
    PFUMX mux_3035_i3 (.BLUT(n4911[2]), .ALUT(n4901[2]), .C0(n32738), 
          .Z(n4920[2]));
    PFUMX mux_3035_i2 (.BLUT(n4911[1]), .ALUT(n4901[1]), .C0(n32738), 
          .Z(n4920[1]));
    PFUMX mux_3035_i1 (.BLUT(n29598), .ALUT(n4901[0]), .C0(n32738), .Z(n4920[0]));
    LUT4 i5450_4_lut_rep_841 (.A(alu_a_in[2]), .B(n34274), .C(n32562), 
         .D(n32625), .Z(n34273)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i5450_4_lut_rep_841.init = 16'haaa8;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module tqvp_uart_tx_U1
//

module tqvp_uart_tx_U1 (debug_uart_txd, clk_c, clk_c_enable_432, cycle_counter, 
            clk_c_enable_143, n6142, n72, \fsm_state[0] , next_bit, 
            n32756, debug_uart_tx_start, \data_to_write[6] , \data_to_write[0] , 
            \data_to_write[5] , \data_to_write[4] , \data_to_write[3] , 
            \data_to_write[2] , \data_to_write[1] , clk_c_enable_495, 
            n32832, uart_txd_N_3005, rst_reg_n, \data_to_write[7] , 
            n26870, n32622) /* synthesis syn_module_defined=1 */ ;
    output debug_uart_txd;
    input clk_c;
    input clk_c_enable_432;
    output [12:0]cycle_counter;
    input clk_c_enable_143;
    input n6142;
    input [12:0]n72;
    output \fsm_state[0] ;
    output next_bit;
    output n32756;
    input debug_uart_tx_start;
    input \data_to_write[6] ;
    input \data_to_write[0] ;
    input \data_to_write[5] ;
    input \data_to_write[4] ;
    input \data_to_write[3] ;
    input \data_to_write[2] ;
    input \data_to_write[1] ;
    input clk_c_enable_495;
    output n32832;
    output uart_txd_N_3005;
    input rst_reg_n;
    input \data_to_write[7] ;
    output n26870;
    output n32622;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire uart_txd_N_3003;
    wire [3:0]fsm_state;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(47[11:20])
    
    wire n31642, n31654, n32861, n9507;
    wire [7:0]data_to_send;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(39[24:36])
    wire [7:0]data_to_send_7__N_2975;
    
    wire n32621, clk_c_enable_211;
    wire [3:0]n162;
    
    wire n26871, n29517, n27946, n29523, n29519, n29513;
    
    FD1S3JX txd_reg_46 (.D(uart_txd_N_3003), .CK(clk_c), .PD(clk_c_enable_432), 
            .Q(debug_uart_txd)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(123[8] 133[4])
    defparam txd_reg_46.GSR = "DISABLED";
    FD1P3IX cycle_counter__i0 (.D(n72[0]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i0.GSR = "DISABLED";
    LUT4 fsm_state_2__bdd_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(\fsm_state[0] ), 
         .Z(n31642)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam fsm_state_2__bdd_3_lut.init = 16'h6a6a;
    FD1P3IX cycle_counter__i12 (.D(n72[12]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i12.GSR = "DISABLED";
    FD1P3IX cycle_counter__i11 (.D(n72[11]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i11.GSR = "DISABLED";
    FD1P3IX cycle_counter__i10 (.D(n72[10]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i10.GSR = "DISABLED";
    FD1P3IX cycle_counter__i9 (.D(n72[9]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i9.GSR = "DISABLED";
    FD1P3IX cycle_counter__i8 (.D(n72[8]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i8.GSR = "DISABLED";
    FD1P3IX cycle_counter__i7 (.D(n72[7]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i7.GSR = "DISABLED";
    FD1P3IX cycle_counter__i6 (.D(n72[6]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i6.GSR = "DISABLED";
    FD1P3IX cycle_counter__i5 (.D(n72[5]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i5.GSR = "DISABLED";
    FD1P3IX cycle_counter__i4 (.D(n72[4]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i4.GSR = "DISABLED";
    FD1P3IX cycle_counter__i3 (.D(n72[3]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i3.GSR = "DISABLED";
    FD1P3IX cycle_counter__i2 (.D(n72[2]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i2.GSR = "DISABLED";
    FD1P3IX cycle_counter__i1 (.D(n72[1]), .SP(clk_c_enable_143), .CD(n6142), 
            .CK(clk_c), .Q(cycle_counter[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i1.GSR = "DISABLED";
    LUT4 fsm_state_3__bdd_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(\fsm_state[0] ), .Z(n31654)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B (C (D))))) */ ;
    defparam fsm_state_3__bdd_4_lut.init = 16'h6aa2;
    LUT4 fsm_state_0__bdd_4_lut (.A(\fsm_state[0] ), .B(fsm_state[2]), .C(fsm_state[1]), 
         .D(fsm_state[3]), .Z(n32861)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;
    defparam fsm_state_0__bdd_4_lut.init = 16'h4555;
    FD1P3IX fsm_state__i3 (.D(n31654), .SP(next_bit), .CD(n9507), .CK(clk_c), 
            .Q(fsm_state[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i3.GSR = "DISABLED";
    FD1P3IX fsm_state__i2 (.D(n31642), .SP(next_bit), .CD(n9507), .CK(clk_c), 
            .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i2.GSR = "DISABLED";
    LUT4 mux_13_i7_3_lut_4_lut (.A(n32756), .B(debug_uart_tx_start), .C(\data_to_write[6] ), 
         .D(data_to_send[7]), .Z(data_to_send_7__N_2975[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut (.A(n32756), .B(debug_uart_tx_start), .C(next_bit), 
         .D(n32621), .Z(clk_c_enable_211)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam i1_3_lut_4_lut.init = 16'hfff4;
    LUT4 mux_13_i1_3_lut_4_lut (.A(n32756), .B(debug_uart_tx_start), .C(\data_to_write[0] ), 
         .D(data_to_send[1]), .Z(data_to_send_7__N_2975[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i6_3_lut_4_lut (.A(n32756), .B(debug_uart_tx_start), .C(\data_to_write[5] ), 
         .D(data_to_send[6]), .Z(data_to_send_7__N_2975[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i5_3_lut_4_lut (.A(n32756), .B(debug_uart_tx_start), .C(\data_to_write[4] ), 
         .D(data_to_send[5]), .Z(data_to_send_7__N_2975[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i4_3_lut_4_lut (.A(n32756), .B(debug_uart_tx_start), .C(\data_to_write[3] ), 
         .D(data_to_send[4]), .Z(data_to_send_7__N_2975[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i4_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX fsm_state__i1 (.D(n162[1]), .SP(next_bit), .CD(n9507), .CK(clk_c), 
            .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i1.GSR = "DISABLED";
    LUT4 mux_13_i3_3_lut_4_lut (.A(n32756), .B(debug_uart_tx_start), .C(\data_to_write[2] ), 
         .D(data_to_send[3]), .Z(data_to_send_7__N_2975[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i2_3_lut_4_lut (.A(n32756), .B(debug_uart_tx_start), .C(\data_to_write[1] ), 
         .D(data_to_send[2]), .Z(data_to_send_7__N_2975[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i2_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX fsm_state__i0 (.D(n32861), .SP(clk_c_enable_211), .CD(n32621), 
            .CK(clk_c), .Q(\fsm_state[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i0.GSR = "DISABLED";
    LUT4 i15177_3_lut_3_lut_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(\fsm_state[0] ), .Z(n162[1])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(D)))) */ ;
    defparam i15177_3_lut_3_lut_4_lut.init = 16'h33c4;
    FD1P3IX data_to_send__i0 (.D(data_to_send_7__N_2975[0]), .SP(clk_c_enable_495), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i0.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_817 (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[3]), 
         .Z(n32832)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_817.init = 16'hfefe;
    LUT4 i1_2_lut_rep_741_4_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[3]), 
         .D(\fsm_state[0] ), .Z(n32756)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_741_4_lut.init = 16'hfffe;
    LUT4 uart_txd_I_270_4_lut_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(fsm_state[3]), .Z(uart_txd_N_3005)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam uart_txd_I_270_4_lut_3_lut.init = 16'h1e1e;
    FD1P3AX data_to_send__i7 (.D(n26871), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(data_to_send[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i7.GSR = "DISABLED";
    FD1P3IX data_to_send__i6 (.D(data_to_send_7__N_2975[6]), .SP(clk_c_enable_495), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i6.GSR = "DISABLED";
    FD1P3IX data_to_send__i5 (.D(data_to_send_7__N_2975[5]), .SP(clk_c_enable_495), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i5.GSR = "DISABLED";
    FD1P3IX data_to_send__i4 (.D(data_to_send_7__N_2975[4]), .SP(clk_c_enable_495), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i4.GSR = "DISABLED";
    FD1P3IX data_to_send__i3 (.D(data_to_send_7__N_2975[3]), .SP(clk_c_enable_495), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i3.GSR = "DISABLED";
    FD1P3IX data_to_send__i2 (.D(data_to_send_7__N_2975[2]), .SP(clk_c_enable_495), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i2.GSR = "DISABLED";
    FD1P3IX data_to_send__i1 (.D(data_to_send_7__N_2975[1]), .SP(clk_c_enable_495), 
            .CD(clk_c_enable_432), .CK(clk_c), .Q(data_to_send[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i1.GSR = "DISABLED";
    LUT4 i14880_4_lut (.A(data_to_send[0]), .B(\fsm_state[0] ), .C(uart_txd_N_3005), 
         .D(n32832), .Z(uart_txd_N_3003)) /* synthesis lut_function=(A ((D)+!B)+!A !(B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(128[14] 132[8])
    defparam i14880_4_lut.init = 16'haf23;
    LUT4 i1_4_lut (.A(n29517), .B(n27946), .C(n29523), .D(n29519), .Z(next_bit)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(cycle_counter[8]), .B(cycle_counter[6]), .Z(n29517)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_286 (.A(n29513), .B(cycle_counter[2]), .C(cycle_counter[0]), 
         .D(cycle_counter[1]), .Z(n27946)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_286.init = 16'haaa8;
    LUT4 i1_4_lut_adj_287 (.A(cycle_counter[5]), .B(cycle_counter[11]), 
         .C(cycle_counter[12]), .D(cycle_counter[9]), .Z(n29523)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_287.init = 16'hfffe;
    LUT4 i1_2_lut_adj_288 (.A(cycle_counter[7]), .B(cycle_counter[10]), 
         .Z(n29519)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_288.init = 16'heeee;
    LUT4 i1_2_lut_adj_289 (.A(cycle_counter[4]), .B(cycle_counter[3]), .Z(n29513)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_289.init = 16'h8888;
    LUT4 i1_2_lut_adj_290 (.A(rst_reg_n), .B(\data_to_write[7] ), .Z(n26870)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_290.init = 16'h8888;
    LUT4 i28400_3_lut_rep_606_4_lut (.A(\fsm_state[0] ), .B(n32832), .C(debug_uart_tx_start), 
         .D(rst_reg_n), .Z(n32621)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i28400_3_lut_rep_606_4_lut.init = 16'h01ff;
    LUT4 i202_2_lut_rep_607_3_lut (.A(\fsm_state[0] ), .B(n32832), .C(debug_uart_tx_start), 
         .Z(n32622)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i202_2_lut_rep_607_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\fsm_state[0] ), .B(n32832), .C(n26870), 
         .D(debug_uart_tx_start), .Z(n26871)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i6825_2_lut_4_lut_2_lut_3_lut (.A(\fsm_state[0] ), .B(n32832), 
         .C(rst_reg_n), .Z(n9507)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i6825_2_lut_4_lut_2_lut_3_lut.init = 16'h1f1f;
    
endmodule
//
// Verilog Description of module sim_qspi_pmod
//

module sim_qspi_pmod (qspi_data_in, qspi_clk_N_56, \addr[14] , \addr_24__N_228[14] , 
            \addr[13] , \addr[12] , \addr[11] , \addr[10] , \addr[9] , 
            GND_net, VCC_net, \addr[8] , \addr[7] , \addr[6] , \addr[5] , 
            \addr[4] , \addr[3] , \addr[0] , \addr[2] , \addr[1] , 
            spi_clk_pos_derived_59, qspi_data_in_3__N_1, \writing_N_164[3] , 
            qspi_ram_a_select, qspi_ram_b_select, n32802, \addr_24__N_228[0] , 
            \addr_24__N_228[1] , \addr_24__N_228[11] , \addr_24__N_228[13] , 
            \addr_24__N_228[12] , \addr_24__N_228[2] , \addr_24__N_228[3] , 
            \addr_24__N_228[4] , \addr_24__N_228[5] , \addr_24__N_228[6] , 
            \addr_24__N_228[7] , \addr_24__N_228[8] , \addr_24__N_228[9] , 
            \addr_24__N_228[10] ) /* synthesis syn_module_defined=1 */ ;
    output [3:0]qspi_data_in;
    input qspi_clk_N_56;
    output \addr[14] ;
    input \addr_24__N_228[14] ;
    output \addr[13] ;
    output \addr[12] ;
    output \addr[11] ;
    output \addr[10] ;
    output \addr[9] ;
    input GND_net;
    input VCC_net;
    output \addr[8] ;
    output \addr[7] ;
    output \addr[6] ;
    output \addr[5] ;
    output \addr[4] ;
    output \addr[3] ;
    output \addr[0] ;
    output \addr[2] ;
    output \addr[1] ;
    input spi_clk_pos_derived_59;
    input [3:0]qspi_data_in_3__N_1;
    input \writing_N_164[3] ;
    input qspi_ram_a_select;
    input qspi_ram_b_select;
    output n32802;
    input \addr_24__N_228[0] ;
    input \addr_24__N_228[1] ;
    input \addr_24__N_228[11] ;
    input \addr_24__N_228[13] ;
    input \addr_24__N_228[12] ;
    input \addr_24__N_228[2] ;
    input \addr_24__N_228[3] ;
    input \addr_24__N_228[4] ;
    input \addr_24__N_228[5] ;
    input \addr_24__N_228[6] ;
    input \addr_24__N_228[7] ;
    input \addr_24__N_228[8] ;
    input \addr_24__N_228[9] ;
    input \addr_24__N_228[10] ;
    
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire [3:0]qspi_data_out_3__N_51;
    
    wire qspi_clk_N_56_enable_1;
    wire [24:0]addr_24__N_89;
    
    wire n24227;
    wire [5:0]start_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(24[15:26])
    wire [5:0]n29;
    
    wire n24226, n24225, n6569, n6577, n6584, n29822, n6573, n6581, 
        n29821, n6570, n6578, n29819, n6574, n6582, n29818, n6571, 
        n6579, n29816, n6575, n6583, n29815;
    wire [7:0]ram_b_buff_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(32[16:30])
    
    wire n29878, n29872, n29854, n29848;
    wire [31:0]cmd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(22[16:19])
    
    wire cmd_31__N_132, rom_buff_out_7__N_118;
    wire [3:0]data_buff_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(29[15:27])
    
    wire spi_clk_pos_derived_59_enable_4, n29873;
    wire [3:0]qspi_data_out_3__N_253;
    
    wire n30131, reading_dummy, qspi_clk_N_56_enable_2, reading_dummy_N_262, 
        n29855, n6548, n6563, n6556, n31680, n6528, n6536, n31681, 
        n6547, n6555, n31683;
    wire [12:0]n6470;
    wire [3:0]qspi_data_out_3__N_257;
    wire [7:0]rom_buff_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(30[16:28])
    
    wire n29849, n29879, n6527, n6535, n31684, reading, writing, 
        error_N_160, reading_N_139, n32870, n6550, n6558, n31702, 
        n29885, n17497, writing_N_151, n32869, qspi_clk_N_56_enable_3, 
        n29886, n6530, n6538, n31703, n29463, n29325, n29321, 
        error, ram_a_buff_out_7__N_127, n26822, n26821, qspi_clk_N_56_enable_4, 
        n11678, qspi_clk_N_56_enable_5, ram_b_buff_out_7__N_128;
    wire [11:0]n6486;
    
    wire ram_b_buff_out_7__N_131, n10665, addr_24__N_224, addr_24__N_204, 
        addr_24__N_200, addr_24__N_202, addr_24__N_222, addr_24__N_220, 
        addr_24__N_218, addr_24__N_216, addr_24__N_214, addr_24__N_212, 
        addr_24__N_210, addr_24__N_208, addr_24__N_206, n29779, n29780, 
        n6549, n6557, n31853, n31854, n6521, n6529, n6537, n6568, 
        n6576, n6572, n6580, n26686, n27878, n29465, n29387, n29251, 
        n29253;
    
    FD1S3AX qspi_data_out_i0 (.D(qspi_data_out_3__N_51[0]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i0.GSR = "DISABLED";
    FD1P3AX addr_i14 (.D(\addr_24__N_228[14] ), .SP(qspi_clk_N_56_enable_1), 
            .CK(qspi_clk_N_56), .Q(\addr[14] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i14.GSR = "ENABLED";
    FD1S3AX addr_i13 (.D(addr_24__N_89[13]), .CK(qspi_clk_N_56), .Q(\addr[13] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i13.GSR = "ENABLED";
    FD1S3AX addr_i12 (.D(addr_24__N_89[12]), .CK(qspi_clk_N_56), .Q(\addr[12] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i12.GSR = "ENABLED";
    FD1S3AX addr_i11 (.D(addr_24__N_89[11]), .CK(qspi_clk_N_56), .Q(\addr[11] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i11.GSR = "ENABLED";
    FD1S3AX addr_i10 (.D(addr_24__N_89[10]), .CK(qspi_clk_N_56), .Q(\addr[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i10.GSR = "ENABLED";
    FD1S3AX addr_i9 (.D(addr_24__N_89[9]), .CK(qspi_clk_N_56), .Q(\addr[9] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i9.GSR = "ENABLED";
    CCU2C start_count_3543_add_4_7 (.A0(start_count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24227), .S0(n29[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543_add_4_7.INIT0 = 16'haaa0;
    defparam start_count_3543_add_4_7.INIT1 = 16'h0000;
    defparam start_count_3543_add_4_7.INJECT1_0 = "NO";
    defparam start_count_3543_add_4_7.INJECT1_1 = "NO";
    CCU2C start_count_3543_add_4_5 (.A0(start_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(start_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24226), .COUT(n24227), .S0(n29[3]), .S1(n29[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543_add_4_5.INIT0 = 16'haaa0;
    defparam start_count_3543_add_4_5.INIT1 = 16'haaa0;
    defparam start_count_3543_add_4_5.INJECT1_0 = "NO";
    defparam start_count_3543_add_4_5.INJECT1_1 = "NO";
    CCU2C start_count_3543_add_4_3 (.A0(start_count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(start_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n24225), .COUT(n24226), .S0(n29[1]), .S1(n29[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543_add_4_3.INIT0 = 16'haaa0;
    defparam start_count_3543_add_4_3.INIT1 = 16'haaa0;
    defparam start_count_3543_add_4_3.INJECT1_0 = "NO";
    defparam start_count_3543_add_4_3.INJECT1_1 = "NO";
    CCU2C start_count_3543_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n24225), .S1(n29[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543_add_4_1.INIT0 = 16'h0000;
    defparam start_count_3543_add_4_1.INIT1 = 16'h555f;
    defparam start_count_3543_add_4_1.INJECT1_0 = "NO";
    defparam start_count_3543_add_4_1.INJECT1_1 = "NO";
    FD1S3AX addr_i8 (.D(addr_24__N_89[8]), .CK(qspi_clk_N_56), .Q(\addr[8] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i8.GSR = "ENABLED";
    LUT4 i27113_3_lut (.A(n6569), .B(n6577), .C(n6584), .Z(n29822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27113_3_lut.init = 16'hcaca;
    LUT4 i27112_3_lut (.A(n6573), .B(n6581), .C(n6584), .Z(n29821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27112_3_lut.init = 16'hcaca;
    LUT4 i27110_3_lut (.A(n6570), .B(n6578), .C(n6584), .Z(n29819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27110_3_lut.init = 16'hcaca;
    LUT4 i27109_3_lut (.A(n6574), .B(n6582), .C(n6584), .Z(n29818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27109_3_lut.init = 16'hcaca;
    LUT4 i27107_3_lut (.A(n6571), .B(n6579), .C(n6584), .Z(n29816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27107_3_lut.init = 16'hcaca;
    LUT4 i27106_3_lut (.A(n6575), .B(n6583), .C(n6584), .Z(n29815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27106_3_lut.init = 16'hcaca;
    FD1S3AX addr_i7 (.D(addr_24__N_89[7]), .CK(qspi_clk_N_56), .Q(\addr[7] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i7.GSR = "ENABLED";
    FD1S3AX addr_i6 (.D(addr_24__N_89[6]), .CK(qspi_clk_N_56), .Q(\addr[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i6.GSR = "ENABLED";
    FD1S3AX addr_i5 (.D(addr_24__N_89[5]), .CK(qspi_clk_N_56), .Q(\addr[5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i5.GSR = "ENABLED";
    FD1S3AX addr_i4 (.D(addr_24__N_89[4]), .CK(qspi_clk_N_56), .Q(\addr[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i4.GSR = "ENABLED";
    FD1S3AX addr_i3 (.D(addr_24__N_89[3]), .CK(qspi_clk_N_56), .Q(\addr[3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i3.GSR = "ENABLED";
    LUT4 i27169_3_lut (.A(ram_b_buff_out[4]), .B(ram_b_buff_out[0]), .C(\addr[0] ), 
         .Z(n29878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27169_3_lut.init = 16'hcaca;
    FD1S3AX addr_i2 (.D(addr_24__N_89[2]), .CK(qspi_clk_N_56), .Q(\addr[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i2.GSR = "ENABLED";
    LUT4 i27163_3_lut (.A(ram_b_buff_out[5]), .B(ram_b_buff_out[1]), .C(\addr[0] ), 
         .Z(n29872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27163_3_lut.init = 16'hcaca;
    LUT4 i27145_3_lut (.A(ram_b_buff_out[6]), .B(ram_b_buff_out[2]), .C(\addr[0] ), 
         .Z(n29854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27145_3_lut.init = 16'hcaca;
    FD1S3AX addr_i1 (.D(addr_24__N_89[1]), .CK(qspi_clk_N_56), .Q(\addr[1] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i1.GSR = "ENABLED";
    LUT4 i27139_3_lut (.A(ram_b_buff_out[7]), .B(ram_b_buff_out[3]), .C(\addr[0] ), 
         .Z(n29848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27139_3_lut.init = 16'hcaca;
    FD1S3AX start_count_3543__i0 (.D(n29[0]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543__i0.GSR = "ENABLED";
    FD1P3AX cmd_i0_i0 (.D(qspi_data_in_3__N_1[0]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i0.GSR = "ENABLED";
    LUT4 i28245_2_lut (.A(\addr[0] ), .B(\writing_N_164[3] ), .Z(rom_buff_out_7__N_118)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i28245_2_lut.init = 16'h1111;
    FD1P3AX data_buff_in_i0_i0 (.D(qspi_data_in_3__N_1[0]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i0.GSR = "DISABLED";
    PFUMX qspi_data_out_3__I_0_i2 (.BLUT(n29873), .ALUT(qspi_data_out_3__N_253[1]), 
          .C0(n30131), .Z(qspi_data_out_3__N_51[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    FD1P3AX reading_dummy_116 (.D(reading_dummy_N_262), .SP(qspi_clk_N_56_enable_2), 
            .CK(qspi_clk_N_56), .Q(reading_dummy)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam reading_dummy_116.GSR = "ENABLED";
    PFUMX qspi_data_out_3__I_0_i3 (.BLUT(n29855), .ALUT(qspi_data_out_3__N_253[2]), 
          .C0(n30131), .Z(qspi_data_out_3__N_51[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    LUT4 n6548_bdd_3_lut_28825 (.A(n6548), .B(n6563), .C(n6556), .Z(n31680)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6548_bdd_3_lut_28825.init = 16'he2e2;
    LUT4 n6548_bdd_3_lut (.A(n6528), .B(n6536), .C(n6563), .Z(n31681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n6548_bdd_3_lut.init = 16'hcaca;
    LUT4 n6547_bdd_3_lut_28828 (.A(n6547), .B(n6563), .C(n6555), .Z(n31683)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6547_bdd_3_lut_28828.init = 16'he2e2;
    FD1S3AX addr_res1_i0_i0 (.D(addr_24__N_89[1]), .CK(qspi_clk_N_56), .Q(n6470[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i0.GSR = "ENABLED";
    LUT4 i27171_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[0]), 
         .C(rom_buff_out[4]), .Z(qspi_data_out_3__N_253[0])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i27171_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27141_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[3]), 
         .C(rom_buff_out[7]), .Z(qspi_data_out_3__N_253[3])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i27141_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27147_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[2]), 
         .C(rom_buff_out[6]), .Z(qspi_data_out_3__N_253[2])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i27147_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27165_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[1]), 
         .C(rom_buff_out[5]), .Z(qspi_data_out_3__N_253[1])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i27165_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27854_3_lut_3_lut (.A(qspi_ram_b_select), .B(n29848), .C(rom_buff_out[3]), 
         .Z(n29849)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i27854_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27844_3_lut_3_lut (.A(qspi_ram_b_select), .B(n29878), .C(rom_buff_out[0]), 
         .Z(n29879)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i27844_3_lut_3_lut.init = 16'he4e4;
    LUT4 n6547_bdd_3_lut (.A(n6527), .B(n6535), .C(n6563), .Z(n31684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n6547_bdd_3_lut.init = 16'hcaca;
    LUT4 i27856_3_lut_3_lut (.A(qspi_ram_b_select), .B(n29854), .C(rom_buff_out[2]), 
         .Z(n29855)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i27856_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27858_3_lut_3_lut (.A(qspi_ram_b_select), .B(n29872), .C(rom_buff_out[1]), 
         .Z(n29873)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i27858_3_lut_3_lut.init = 16'he4e4;
    LUT4 reading_I_0_126_2_lut_rep_843 (.A(reading), .B(writing), .Z(qspi_clk_N_56_enable_1)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam reading_I_0_126_2_lut_rep_843.init = 16'heeee;
    PFUMX qspi_data_out_3__I_0_i4 (.BLUT(n29849), .ALUT(qspi_data_out_3__N_253[3]), 
          .C0(n30131), .Z(qspi_data_out_3__N_51[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    LUT4 i28413_3_lut_rep_787 (.A(\writing_N_164[3] ), .B(qspi_ram_b_select), 
         .C(qspi_ram_a_select), .Z(n32802)) /* synthesis lut_function=(!(A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(34[23:82])
    defparam i28413_3_lut_rep_787.init = 16'h7f7f;
    LUT4 i28409_2_lut_4_lut (.A(\writing_N_164[3] ), .B(qspi_ram_b_select), 
         .C(qspi_ram_a_select), .D(\addr[0] ), .Z(spi_clk_pos_derived_59_enable_4)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(34[23:82])
    defparam i28409_2_lut_4_lut.init = 16'h007f;
    LUT4 i28386_4_lut_then_3_lut_4_lut (.A(reading), .B(writing), .C(error_N_160), 
         .D(reading_N_139), .Z(n32870)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i28386_4_lut_then_3_lut_4_lut.init = 16'h1110;
    PFUMX qspi_data_out_3__I_0_i1 (.BLUT(n29879), .ALUT(qspi_data_out_3__N_253[0]), 
          .C0(n30131), .Z(qspi_data_out_3__N_51[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    FD1S3AX qspi_data_out_i3 (.D(qspi_data_out_3__N_51[3]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i3.GSR = "DISABLED";
    FD1S3AX qspi_data_out_i2 (.D(qspi_data_out_3__N_51[2]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i2.GSR = "DISABLED";
    LUT4 n6550_bdd_3_lut_28842 (.A(n6550), .B(n6563), .C(n6558), .Z(n31702)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6550_bdd_3_lut_28842.init = 16'he2e2;
    FD1S3AX qspi_data_out_i1 (.D(qspi_data_out_3__N_51[1]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i1.GSR = "DISABLED";
    FD1P3AX reading_115 (.D(n29885), .SP(reading_N_139), .CK(qspi_clk_N_56), 
            .Q(reading)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam reading_115.GSR = "ENABLED";
    LUT4 i28386_4_lut_else_3_lut_4_lut (.A(reading), .B(writing), .C(n17497), 
         .D(writing_N_151), .Z(n32869)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i28386_4_lut_else_3_lut_4_lut.init = 16'h0100;
    FD1P3AX writing_117 (.D(n29886), .SP(qspi_clk_N_56_enable_3), .CK(qspi_clk_N_56), 
            .Q(writing)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam writing_117.GSR = "ENABLED";
    LUT4 n6550_bdd_3_lut (.A(n6530), .B(n6538), .C(n6563), .Z(n31703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n6550_bdd_3_lut.init = 16'hcaca;
    FD1S3AX start_count_3543__i1 (.D(n29[1]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543__i1.GSR = "ENABLED";
    FD1S3AX start_count_3543__i2 (.D(n29[2]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543__i2.GSR = "ENABLED";
    FD1S3AX start_count_3543__i3 (.D(n29[3]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543__i3.GSR = "ENABLED";
    FD1S3AX start_count_3543__i4 (.D(n29[4]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543__i4.GSR = "ENABLED";
    FD1S3AX start_count_3543__i5 (.D(n29[5]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3543__i5.GSR = "ENABLED";
    FD1P3AX cmd_i0_i1 (.D(qspi_data_in_3__N_1[1]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i1.GSR = "ENABLED";
    FD1P3AX cmd_i0_i2 (.D(qspi_data_in_3__N_1[2]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i2.GSR = "ENABLED";
    FD1P3AX cmd_i0_i3 (.D(qspi_data_in_3__N_1[3]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i3.GSR = "ENABLED";
    FD1P3AX cmd_i0_i4 (.D(cmd[0]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i4.GSR = "ENABLED";
    FD1P3AX cmd_i0_i5 (.D(cmd[1]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i5.GSR = "ENABLED";
    FD1P3AX cmd_i0_i6 (.D(cmd[2]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i6.GSR = "ENABLED";
    FD1P3AX cmd_i0_i7 (.D(cmd[3]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i7.GSR = "ENABLED";
    FD1P3AX cmd_i0_i8 (.D(cmd[4]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i8.GSR = "ENABLED";
    FD1P3AX cmd_i0_i9 (.D(cmd[5]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i9.GSR = "ENABLED";
    FD1P3AX cmd_i0_i10 (.D(cmd[6]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i10.GSR = "ENABLED";
    FD1P3AX cmd_i0_i11 (.D(cmd[7]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i11.GSR = "ENABLED";
    FD1P3AX cmd_i0_i12 (.D(cmd[8]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i12.GSR = "ENABLED";
    FD1P3AX cmd_i0_i13 (.D(cmd[9]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i13.GSR = "ENABLED";
    FD1P3AX cmd_i0_i14 (.D(cmd[10]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i14.GSR = "ENABLED";
    FD1P3AX cmd_i0_i15 (.D(cmd[11]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i15.GSR = "ENABLED";
    FD1P3AX cmd_i0_i16 (.D(cmd[12]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i16.GSR = "ENABLED";
    FD1P3AX cmd_i0_i17 (.D(cmd[13]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i17.GSR = "ENABLED";
    FD1P3AX cmd_i0_i18 (.D(cmd[14]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i18.GSR = "ENABLED";
    FD1P3AX cmd_i0_i19 (.D(cmd[15]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i19.GSR = "ENABLED";
    FD1P3AX cmd_i0_i20 (.D(cmd[16]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i20.GSR = "ENABLED";
    FD1P3AX cmd_i0_i21 (.D(cmd[17]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i21.GSR = "ENABLED";
    FD1P3AX cmd_i0_i22 (.D(cmd[18]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i22.GSR = "ENABLED";
    FD1P3AX cmd_i0_i23 (.D(cmd[19]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i23.GSR = "ENABLED";
    FD1P3AX cmd_i0_i24 (.D(cmd[20]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i24.GSR = "ENABLED";
    FD1P3AX cmd_i0_i25 (.D(cmd[21]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i25.GSR = "ENABLED";
    FD1P3AX cmd_i0_i26 (.D(cmd[22]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i26.GSR = "ENABLED";
    FD1P3AX cmd_i0_i27 (.D(cmd[23]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i27.GSR = "ENABLED";
    FD1P3AX cmd_i0_i28 (.D(cmd[24]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i28.GSR = "ENABLED";
    FD1P3AX cmd_i0_i29 (.D(cmd[25]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i29.GSR = "ENABLED";
    FD1P3AX cmd_i0_i30 (.D(cmd[26]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i30.GSR = "ENABLED";
    FD1P3AX cmd_i0_i31 (.D(cmd[27]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i31.GSR = "ENABLED";
    FD1P3AX data_buff_in_i0_i1 (.D(qspi_data_in_3__N_1[1]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i1.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(start_count[3]), .B(n29463), .C(n29325), .D(\writing_N_164[3] ), 
         .Z(writing_N_151)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h2010;
    FD1P3AX data_buff_in_i0_i2 (.D(qspi_data_in_3__N_1[2]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i2.GSR = "DISABLED";
    FD1P3AX data_buff_in_i0_i3 (.D(qspi_data_in_3__N_1[3]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i3.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_275 (.A(start_count[0]), .B(n29321), .C(start_count[1]), 
         .D(\writing_N_164[3] ), .Z(n29325)) /* synthesis lut_function=(!(A+((C (D)+!C !(D))+!B))) */ ;
    defparam i1_4_lut_adj_275.init = 16'h0440;
    LUT4 i1_3_lut (.A(start_count[2]), .B(error), .C(\writing_N_164[3] ), 
         .Z(n29321)) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(C)))) */ ;
    defparam i1_3_lut.init = 16'h1212;
    LUT4 i1_2_lut (.A(start_count[4]), .B(start_count[5]), .Z(n29463)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(93[21:38])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i28248_2_lut (.A(\addr[0] ), .B(qspi_ram_a_select), .Z(ram_a_buff_out_7__N_127)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i28248_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_4_lut (.A(writing), .B(\addr[0] ), .C(\addr[12] ), 
         .D(qspi_ram_a_select), .Z(n26822)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(49[14:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_276 (.A(writing), .B(\addr[0] ), .C(\addr[12] ), 
         .D(qspi_ram_a_select), .Z(n26821)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(49[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_276.init = 16'h0008;
    FD1P3IX addr_i0 (.D(\addr_24__N_228[0] ), .SP(qspi_clk_N_56_enable_4), 
            .CD(n11678), .CK(qspi_clk_N_56), .Q(\addr[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i0.GSR = "ENABLED";
    FD1P3AX error_118 (.D(VCC_net), .SP(qspi_clk_N_56_enable_5), .CK(qspi_clk_N_56), 
            .Q(error)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam error_118.GSR = "ENABLED";
    LUT4 ram_a_buff_out_7__N_124_I_0_2_lut_3_lut (.A(writing), .B(\addr[0] ), 
         .C(qspi_ram_b_select), .Z(ram_b_buff_out_7__N_128)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(49[14:31])
    defparam ram_a_buff_out_7__N_124_I_0_2_lut_3_lut.init = 16'h0808;
    FD1S3AX addr_res2_i0_i11 (.D(addr_24__N_89[12]), .CK(qspi_clk_N_56), 
            .Q(n6486[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res2_i0_i11.GSR = "ENABLED";
    LUT4 i28253_2_lut (.A(\addr[0] ), .B(qspi_ram_b_select), .Z(ram_b_buff_out_7__N_131)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i28253_2_lut.init = 16'h1111;
    LUT4 i27177_4_lut_4_lut_4_lut (.A(reading), .B(writing), .C(n10665), 
         .D(n17497), .Z(n29886)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i27177_4_lut_4_lut_4_lut.init = 16'hcdcc;
    LUT4 i1_2_lut_3_lut_4_lut_adj_277 (.A(reading), .B(writing), .C(reading_dummy), 
         .D(writing_N_151), .Z(qspi_clk_N_56_enable_4)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i1_2_lut_3_lut_4_lut_adj_277.init = 16'hefee;
    LUT4 addr_24__I_0_i2_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[1] ), 
         .D(addr_24__N_224), .Z(addr_24__N_89[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i12_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[11] ), 
         .D(addr_24__N_204), .Z(addr_24__N_89[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i8970_2_lut_3_lut_4_lut (.A(reading), .B(writing), .C(reading_dummy), 
         .D(writing_N_151), .Z(n11678)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i8970_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 addr_24__I_0_i14_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[13] ), 
         .D(addr_24__N_200), .Z(addr_24__N_89[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i13_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[12] ), 
         .D(addr_24__N_202), .Z(addr_24__N_89[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i3_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[2] ), 
         .D(addr_24__N_222), .Z(addr_24__N_89[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i3_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX addr_res1_i0_i1 (.D(addr_24__N_89[2]), .CK(qspi_clk_N_56), .Q(n6470[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i1.GSR = "ENABLED";
    PFUMX i29313 (.BLUT(n32869), .ALUT(n32870), .C0(reading_dummy), .Z(qspi_clk_N_56_enable_2));
    LUT4 addr_24__I_0_i4_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[3] ), 
         .D(addr_24__N_220), .Z(addr_24__N_89[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i5_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[4] ), 
         .D(addr_24__N_218), .Z(addr_24__N_89[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i6_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[5] ), 
         .D(addr_24__N_216), .Z(addr_24__N_89[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i6_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX addr_res1_i0_i2 (.D(addr_24__N_89[3]), .CK(qspi_clk_N_56), .Q(n6470[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i2.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i3 (.D(addr_24__N_89[4]), .CK(qspi_clk_N_56), .Q(n6470[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i3.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i4 (.D(addr_24__N_89[5]), .CK(qspi_clk_N_56), .Q(n6470[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i4.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i5 (.D(addr_24__N_89[6]), .CK(qspi_clk_N_56), .Q(n6470[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i5.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i6 (.D(addr_24__N_89[7]), .CK(qspi_clk_N_56), .Q(n6470[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i6.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i7 (.D(addr_24__N_89[8]), .CK(qspi_clk_N_56), .Q(n6470[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i7.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i8 (.D(addr_24__N_89[9]), .CK(qspi_clk_N_56), .Q(n6470[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i8.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i9 (.D(addr_24__N_89[10]), .CK(qspi_clk_N_56), 
            .Q(n6470[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i9.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i10 (.D(addr_24__N_89[11]), .CK(qspi_clk_N_56), 
            .Q(n6470[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i10.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i12 (.D(addr_24__N_89[13]), .CK(qspi_clk_N_56), 
            .Q(n6470[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i12.GSR = "ENABLED";
    LUT4 addr_24__I_0_i7_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[6] ), 
         .D(addr_24__N_214), .Z(addr_24__N_89[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i8_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[7] ), 
         .D(addr_24__N_212), .Z(addr_24__N_89[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i9_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[8] ), 
         .D(addr_24__N_210), .Z(addr_24__N_89[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i10_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[9] ), 
         .D(addr_24__N_208), .Z(addr_24__N_89[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i11_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[10] ), 
         .D(addr_24__N_206), .Z(addr_24__N_89[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i11_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i27072 (.BLUT(n29779), .ALUT(n29780), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[0]));
    LUT4 i27176_4_lut_3_lut (.A(reading), .B(writing), .C(reading_dummy), 
         .Z(n29885)) /* synthesis lut_function=(A+!(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i27176_4_lut_3_lut.init = 16'hbaba;
    LUT4 n6549_bdd_3_lut_28944 (.A(n6549), .B(n6563), .C(n6557), .Z(n31853)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6549_bdd_3_lut_28944.init = 16'he2e2;
    PFUMX i28945 (.BLUT(n31854), .ALUT(n31853), .C0(n6521), .Z(rom_buff_out[2]));
    LUT4 n6549_bdd_3_lut (.A(n6529), .B(n6537), .C(n6563), .Z(n31854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n6549_bdd_3_lut.init = 16'hcaca;
    LUT4 i27071_3_lut (.A(n6568), .B(n6576), .C(n6584), .Z(n29780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27071_3_lut.init = 16'hcaca;
    LUT4 i27070_3_lut (.A(n6572), .B(n6580), .C(n6584), .Z(n29779)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27070_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_278 (.A(cmd[27]), .B(n26686), .C(cmd[24]), .Z(n10665)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(102[26:45])
    defparam i1_3_lut_adj_278.init = 16'hfefe;
    LUT4 i8883_2_lut_3_lut (.A(n17497), .B(writing_N_151), .C(reading_dummy), 
         .Z(reading_dummy_N_262)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i8883_2_lut_3_lut.init = 16'h0404;
    PFUMX i28843 (.BLUT(n31703), .ALUT(n31702), .C0(n6521), .Z(rom_buff_out[3]));
    LUT4 i28520_3_lut (.A(reading), .B(writing), .C(error), .Z(cmd_31__N_132)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i28520_3_lut.init = 16'h0101;
    LUT4 i5269_2_lut_rep_683 (.A(writing_N_151), .B(reading_dummy), .Z(qspi_clk_N_56_enable_3)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5269_2_lut_rep_683.init = 16'h2222;
    LUT4 i5270_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[12]), 
         .D(\addr[13] ), .Z(addr_24__N_200)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5270_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5272_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[11]), 
         .D(\addr[12] ), .Z(addr_24__N_202)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5272_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5274_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[10]), 
         .D(\addr[11] ), .Z(addr_24__N_204)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5274_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5276_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[9]), 
         .D(\addr[10] ), .Z(addr_24__N_206)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5276_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5278_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[8]), 
         .D(\addr[9] ), .Z(addr_24__N_208)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5278_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5280_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[7]), 
         .D(\addr[8] ), .Z(addr_24__N_210)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5280_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5282_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[6]), 
         .D(\addr[7] ), .Z(addr_24__N_212)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5282_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5284_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[5]), 
         .D(\addr[6] ), .Z(addr_24__N_214)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5284_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5286_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[4]), 
         .D(\addr[5] ), .Z(addr_24__N_216)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5286_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5288_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[3]), 
         .D(\addr[4] ), .Z(addr_24__N_218)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5288_3_lut_4_lut.init = 16'hfd20;
    LUT4 i28250_4_lut (.A(n27878), .B(qspi_clk_N_56_enable_1), .C(error_N_160), 
         .D(reading_dummy), .Z(qspi_clk_N_56_enable_5)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i28250_4_lut.init = 16'h3022;
    LUT4 i1_3_lut_adj_279 (.A(writing_N_151), .B(n17497), .C(n10665), 
         .Z(n27878)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_279.init = 16'h8080;
    LUT4 i5290_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[2]), 
         .D(\addr[3] ), .Z(addr_24__N_220)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5290_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5292_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[1]), 
         .D(\addr[2] ), .Z(addr_24__N_222)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5292_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5294_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[0]), 
         .D(\addr[1] ), .Z(addr_24__N_224)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5294_3_lut_4_lut.init = 16'hfd20;
    PFUMX i28829 (.BLUT(n31684), .ALUT(n31683), .C0(n6521), .Z(rom_buff_out[0]));
    LUT4 i28580_3_lut (.A(qspi_ram_a_select), .B(qspi_ram_b_select), .C(\addr[0] ), 
         .Z(n30131)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26] 113[96])
    defparam i28580_3_lut.init = 16'h5d5d;
    PFUMX i28826 (.BLUT(n31681), .ALUT(n31680), .C0(n6521), .Z(rom_buff_out[1]));
    LUT4 i28327_4_lut (.A(start_count[2]), .B(start_count[3]), .C(n29465), 
         .D(n29463), .Z(reading_N_139)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(93[21:38])
    defparam i28327_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_adj_280 (.A(start_count[0]), .B(start_count[1]), .Z(n29465)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(93[21:38])
    defparam i1_2_lut_adj_280.init = 16'heeee;
    LUT4 i1_4_lut_adj_281 (.A(n29387), .B(n29463), .C(start_count[3]), 
         .D(cmd[1]), .Z(error_N_160)) /* synthesis lut_function=(!(A (B+(C))+!A (B+(C+(D))))) */ ;
    defparam i1_4_lut_adj_281.init = 16'h0203;
    LUT4 i1_3_lut_adj_282 (.A(cmd[3]), .B(cmd[0]), .C(cmd[2]), .Z(n29387)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_3_lut_adj_282.init = 16'hfdfd;
    LUT4 i14850_4_lut (.A(\writing_N_164[3] ), .B(cmd[27]), .C(n26686), 
         .D(cmd[24]), .Z(n17497)) /* synthesis lut_function=(A ((C+!(D))+!B)) */ ;
    defparam i14850_4_lut.init = 16'ha2aa;
    LUT4 i1_4_lut_adj_283 (.A(n29251), .B(cmd[25]), .C(n29253), .D(cmd[26]), 
         .Z(n26686)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(102[26:45])
    defparam i1_4_lut_adj_283.init = 16'hfffb;
    LUT4 i1_2_lut_adj_284 (.A(cmd[29]), .B(cmd[30]), .Z(n29251)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(102[26:45])
    defparam i1_2_lut_adj_284.init = 16'heeee;
    LUT4 i1_2_lut_adj_285 (.A(cmd[31]), .B(cmd[28]), .Z(n29253)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(102[26:45])
    defparam i1_2_lut_adj_285.init = 16'heeee;
    PFUMX i27108 (.BLUT(n29815), .ALUT(n29816), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[3]));
    PFUMX i27111 (.BLUT(n29818), .ALUT(n29819), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[2]));
    PFUMX i27114 (.BLUT(n29821), .ALUT(n29822), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[1]));
    \BRAM(ADDR_WIDTH=13)  rom (.n6563(n6563), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .rom_buff_out_7__N_118(rom_buff_out_7__N_118), .n6475(n6486[11]), 
            .\addr[1] (\addr[1] ), .\addr[2] (\addr[2] ), .\addr[3] (\addr[3] ), 
            .\addr[4] (\addr[4] ), .\addr[5] (\addr[5] ), .\addr[6] (\addr[6] ), 
            .\addr[7] (\addr[7] ), .\addr[8] (\addr[8] ), .\addr[9] (\addr[9] ), 
            .\addr[10] (\addr[10] ), .\addr[11] (\addr[11] ), .n6474(n6470[0]), 
            .n6469(n6470[1]), .n6468(n6470[2]), .n6467(n6470[3]), .n6466(n6470[4]), 
            .n6465(n6470[5]), .n6464(n6470[6]), .n6463(n6470[7]), .n6462(n6470[8]), 
            .n6461(n6470[9]), .n6460(n6470[10]), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .data_buff_in({data_buff_in}), .n6555(n6555), .n6556(n6556), 
            .n6557(n6557), .n6558(n6558), .GND_net(GND_net), .VCC_net(VCC_net), 
            .n6547(n6547), .n6548(n6548), .n6549(n6549), .n6550(n6550), 
            .n6527(n6527), .n6528(n6528), .n6529(n6529), .n6530(n6530), 
            .n6535(n6535), .n6536(n6536), .n6537(n6537), .n6538(n6538), 
            .n6521(n6521), .n6458(n6470[12]), .\rom_buff_out[7] (rom_buff_out[7]), 
            .\rom_buff_out[6] (rom_buff_out[6]), .\rom_buff_out[5] (rom_buff_out[5]), 
            .\rom_buff_out[4] (rom_buff_out[4])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(36[58] 43[6])
    \BRAM(ADDR_WIDTH=11)  ram_b (.\addr[1] (\addr[1] ), .\addr[2] (\addr[2] ), 
            .\addr[3] (\addr[3] ), .\addr[4] (\addr[4] ), .\addr[5] (\addr[5] ), 
            .\addr[6] (\addr[6] ), .\addr[7] (\addr[7] ), .\addr[8] (\addr[8] ), 
            .\addr[9] (\addr[9] ), .\addr[10] (\addr[10] ), .\addr[11] (\addr[11] ), 
            .n6474(n6470[0]), .n6469(n6470[1]), .n6468(n6470[2]), .n6467(n6470[3]), 
            .n6466(n6470[4]), .n6465(n6470[5]), .n6464(n6470[6]), .n6463(n6470[7]), 
            .n6462(n6470[8]), .n6461(n6470[9]), .n6460(n6470[10]), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .data_buff_in({data_buff_in}), .ram_b_buff_out({ram_b_buff_out}), 
            .spi_clk_pos_derived_59(spi_clk_pos_derived_59), .ram_b_buff_out_7__N_128(ram_b_buff_out_7__N_128), 
            .ram_b_buff_out_7__N_131(ram_b_buff_out_7__N_131), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(52[37] 59[6])
    \BRAM(ADDR_WIDTH=12)  ram_a (.\addr[1] (\addr[1] ), .\addr[2] (\addr[2] ), 
            .\addr[3] (\addr[3] ), .\addr[4] (\addr[4] ), .\addr[5] (\addr[5] ), 
            .\addr[6] (\addr[6] ), .\addr[7] (\addr[7] ), .\addr[8] (\addr[8] ), 
            .\addr[9] (\addr[9] ), .\addr[10] (\addr[10] ), .\addr[11] (\addr[11] ), 
            .n6474(n6470[0]), .n6469(n6470[1]), .n6468(n6470[2]), .n6467(n6470[3]), 
            .n6466(n6470[4]), .n6465(n6470[5]), .n6464(n6470[6]), .n6463(n6470[7]), 
            .n6462(n6470[8]), .n6461(n6470[9]), .n6460(n6470[10]), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .data_buff_in({data_buff_in}), .n6576(n6576), .n6577(n6577), 
            .n6578(n6578), .n6579(n6579), .n6580(n6580), .n6581(n6581), 
            .n6582(n6582), .n6583(n6583), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .n26822(n26822), .ram_a_buff_out_7__N_127(ram_a_buff_out_7__N_127), 
            .GND_net(GND_net), .VCC_net(VCC_net), .n6568(n6568), .n6569(n6569), 
            .n6570(n6570), .n6571(n6571), .n6572(n6572), .n6573(n6573), 
            .n6574(n6574), .n6575(n6575), .n26821(n26821), .n6584(n6584), 
            .n6475(n6486[11])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(44[37] 51[6])
    
endmodule
//
// Verilog Description of module \BRAM(ADDR_WIDTH=13) 
//

module \BRAM(ADDR_WIDTH=13)  (n6563, spi_clk_pos_derived_59, rom_buff_out_7__N_118, 
            n6475, \addr[1] , \addr[2] , \addr[3] , \addr[4] , \addr[5] , 
            \addr[6] , \addr[7] , \addr[8] , \addr[9] , \addr[10] , 
            \addr[11] , n6474, n6469, n6468, n6467, n6466, n6465, 
            n6464, n6463, n6462, n6461, n6460, qspi_data_in_3__N_1, 
            data_buff_in, n6555, n6556, n6557, n6558, GND_net, VCC_net, 
            n6547, n6548, n6549, n6550, n6527, n6528, n6529, n6530, 
            n6535, n6536, n6537, n6538, n6521, n6458, \rom_buff_out[7] , 
            \rom_buff_out[6] , \rom_buff_out[5] , \rom_buff_out[4] ) /* synthesis syn_module_defined=1 */ ;
    output n6563;
    input spi_clk_pos_derived_59;
    input rom_buff_out_7__N_118;
    input n6475;
    input \addr[1] ;
    input \addr[2] ;
    input \addr[3] ;
    input \addr[4] ;
    input \addr[5] ;
    input \addr[6] ;
    input \addr[7] ;
    input \addr[8] ;
    input \addr[9] ;
    input \addr[10] ;
    input \addr[11] ;
    input n6474;
    input n6469;
    input n6468;
    input n6467;
    input n6466;
    input n6465;
    input n6464;
    input n6463;
    input n6462;
    input n6461;
    input n6460;
    input [3:0]qspi_data_in_3__N_1;
    input [3:0]data_buff_in;
    output n6555;
    output n6556;
    output n6557;
    output n6558;
    input GND_net;
    input VCC_net;
    output n6547;
    output n6548;
    output n6549;
    output n6550;
    output n6527;
    output n6528;
    output n6529;
    output n6530;
    output n6535;
    output n6536;
    output n6537;
    output n6538;
    output n6521;
    input n6458;
    output \rom_buff_out[7] ;
    output \rom_buff_out[6] ;
    output \rom_buff_out[5] ;
    output \rom_buff_out[4] ;
    
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    wire n6551, n6559, n29801, n6531, n6539, n29800, n6560, n6561, 
        n6562, n6552, n6553, n6554, n6532, n6533, n6534, n6540, 
        n6541, n6542, n29798, n29797, n29795, n29794, n29792, 
        n29791;
    
    FD1P3AX i4295 (.D(n6475), .SP(rom_buff_out_7__N_118), .CK(spi_clk_pos_derived_59), 
            .Q(n6563));
    defparam i4295.GSR = "DISABLED";
    LUT4 i27092_3_lut (.A(n6551), .B(n6559), .C(n6563), .Z(n29801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27092_3_lut.init = 16'hcaca;
    LUT4 i27091_3_lut (.A(n6531), .B(n6539), .C(n6563), .Z(n29800)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27091_3_lut.init = 16'hcaca;
    DP16KD mem3 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6474), .ADB4(n6469), 
           .ADB5(n6468), .ADB6(n6467), .ADB7(n6466), .ADB8(n6465), .ADB9(n6464), 
           .ADB10(n6463), .ADB11(n6462), .ADB12(n6461), .ADB13(n6460), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6555), .DOB1(n6556), .DOB2(n6557), 
           .DOB3(n6558), .DOB4(n6559), .DOB5(n6560), .DOB6(n6561), .DOB7(n6562));
    defparam mem3.DATA_WIDTH_A = 9;
    defparam mem3.DATA_WIDTH_B = 9;
    defparam mem3.REGMODE_A = "NOREG";
    defparam mem3.REGMODE_B = "NOREG";
    defparam mem3.RESETMODE = "SYNC";
    defparam mem3.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem3.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem3.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem3.CSDECODE_A = "0b000";
    defparam mem3.CSDECODE_B = "0b000";
    defparam mem3.GSR = "DISABLED";
    defparam mem3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INIT_DATA = "STATIC";
    DP16KD mem1 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6474), .ADB4(n6469), 
           .ADB5(n6468), .ADB6(n6467), .ADB7(n6466), .ADB8(n6465), .ADB9(n6464), 
           .ADB10(n6463), .ADB11(n6462), .ADB12(n6461), .ADB13(n6460), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6547), .DOB1(n6548), .DOB2(n6549), 
           .DOB3(n6550), .DOB4(n6551), .DOB5(n6552), .DOB6(n6553), .DOB7(n6554));
    defparam mem1.DATA_WIDTH_A = 9;
    defparam mem1.DATA_WIDTH_B = 9;
    defparam mem1.REGMODE_A = "NOREG";
    defparam mem1.REGMODE_B = "NOREG";
    defparam mem1.RESETMODE = "SYNC";
    defparam mem1.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem1.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem1.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem1.CSDECODE_A = "0b000";
    defparam mem1.CSDECODE_B = "0b000";
    defparam mem1.GSR = "DISABLED";
    defparam mem1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INIT_DATA = "STATIC";
    DP16KD mem0 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6474), .ADB4(n6469), 
           .ADB5(n6468), .ADB6(n6467), .ADB7(n6466), .ADB8(n6465), .ADB9(n6464), 
           .ADB10(n6463), .ADB11(n6462), .ADB12(n6461), .ADB13(n6460), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6527), .DOB1(n6528), .DOB2(n6529), 
           .DOB3(n6530), .DOB4(n6531), .DOB5(n6532), .DOB6(n6533), .DOB7(n6534));
    defparam mem0.DATA_WIDTH_A = 9;
    defparam mem0.DATA_WIDTH_B = 9;
    defparam mem0.REGMODE_A = "NOREG";
    defparam mem0.REGMODE_B = "NOREG";
    defparam mem0.RESETMODE = "SYNC";
    defparam mem0.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem0.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem0.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem0.CSDECODE_A = "0b000";
    defparam mem0.CSDECODE_B = "0b000";
    defparam mem0.GSR = "DISABLED";
    defparam mem0.INITVAL_00 = "0x00000000000000000004108E7080840088A002F50E8930682004A731E02400C800006F00A000006F";
    defparam mem0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_02 = "0x00280002170100000437080011029300200002B70000000244000000008000000000700000000070";
    defparam mem0.INITVAL_03 = "0x0602000073068820684416073000A4128B30888506020000731400105079004C0000EF1F44100213";
    defparam mem0.INITVAL_04 = "0x1D80110E93000E61F2631D80110E131D80110C930602000073068820604416073000A4128B308885";
    defparam mem0.INITVAL_05 = "0x11C911FEF710C93004F60EA630008710E931800110C130020000EB71FCE71DAE300EC1000071C023";
    defparam mem0.INITVAL_06 = "0x1FCD7136E31FCC705C2300E1100E9108690036C000E9312CB21800110E1300C91036C000C13134F1";
    defparam mem0.INITVAL_07 = "0x00EC100E41000A71E023000070EA030404000E131D80110E93000670FC631D801106131D80110E13";
    defparam mem0.INITVAL_08 = "0x00E130800510A930000302CB70200000E370100000AB71A6B80100000EB708E41100821FC671D4E3";
    defparam mem0.INITVAL_09 = "0x1FCE311E910861C0861000005100231FCF61FCE311E910861C086101128808A051A6F610C931E007";
    defparam mem0.INITVAL_0A = "0x06882180A1144230009500E63188811089300A051D026102040049500263180011688316EDD1FCF6";
    defparam mem0.INITVAL_0B = "0x1607308CA11888110E1306020000730688206045060730000800A3717ECD1808110A130602000073";
    defparam mem0.INITVAL_0C = "0x1407306045140730000800AB7180B114023000B601C63000E511A6300A85112881800116A8306006";
    defparam mem0.INITVAL_0D = "0x002000000817EE106006160731FCE601CE31804114E03060061407316EDD1808110A931008206006";
    defparam mem0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000020000008";
    defparam mem0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INIT_DATA = "STATIC";
    DP16KD mem2 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6474), .ADB4(n6469), 
           .ADB5(n6468), .ADB6(n6467), .ADB7(n6466), .ADB8(n6465), .ADB9(n6464), 
           .ADB10(n6463), .ADB11(n6462), .ADB12(n6461), .ADB13(n6460), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6535), .DOB1(n6536), .DOB2(n6537), 
           .DOB3(n6538), .DOB4(n6539), .DOB5(n6540), .DOB6(n6541), .DOB7(n6542));
    defparam mem2.DATA_WIDTH_A = 9;
    defparam mem2.DATA_WIDTH_B = 9;
    defparam mem2.REGMODE_A = "NOREG";
    defparam mem2.REGMODE_B = "NOREG";
    defparam mem2.RESETMODE = "SYNC";
    defparam mem2.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem2.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem2.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem2.CSDECODE_A = "0b000";
    defparam mem2.CSDECODE_B = "0b000";
    defparam mem2.GSR = "DISABLED";
    defparam mem2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INIT_DATA = "STATIC";
    LUT4 i27089_3_lut (.A(n6552), .B(n6560), .C(n6563), .Z(n29798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27089_3_lut.init = 16'hcaca;
    LUT4 i27088_3_lut (.A(n6532), .B(n6540), .C(n6563), .Z(n29797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27088_3_lut.init = 16'hcaca;
    LUT4 i27086_3_lut (.A(n6553), .B(n6561), .C(n6563), .Z(n29795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27086_3_lut.init = 16'hcaca;
    FD1P3AX i4277 (.D(n6458), .SP(rom_buff_out_7__N_118), .CK(spi_clk_pos_derived_59), 
            .Q(n6521));
    defparam i4277.GSR = "DISABLED";
    LUT4 i27085_3_lut (.A(n6533), .B(n6541), .C(n6563), .Z(n29794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27085_3_lut.init = 16'hcaca;
    LUT4 i27083_3_lut (.A(n6554), .B(n6562), .C(n6563), .Z(n29792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27083_3_lut.init = 16'hcaca;
    LUT4 i27082_3_lut (.A(n6534), .B(n6542), .C(n6563), .Z(n29791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27082_3_lut.init = 16'hcaca;
    PFUMX i27084 (.BLUT(n29791), .ALUT(n29792), .C0(n6521), .Z(\rom_buff_out[7] ));
    PFUMX i27087 (.BLUT(n29794), .ALUT(n29795), .C0(n6521), .Z(\rom_buff_out[6] ));
    PFUMX i27090 (.BLUT(n29797), .ALUT(n29798), .C0(n6521), .Z(\rom_buff_out[5] ));
    PFUMX i27093 (.BLUT(n29800), .ALUT(n29801), .C0(n6521), .Z(\rom_buff_out[4] ));
    
endmodule
//
// Verilog Description of module \BRAM(ADDR_WIDTH=11) 
//

module \BRAM(ADDR_WIDTH=11)  (\addr[1] , \addr[2] , \addr[3] , \addr[4] , 
            \addr[5] , \addr[6] , \addr[7] , \addr[8] , \addr[9] , 
            \addr[10] , \addr[11] , n6474, n6469, n6468, n6467, 
            n6466, n6465, n6464, n6463, n6462, n6461, n6460, qspi_data_in_3__N_1, 
            data_buff_in, ram_b_buff_out, spi_clk_pos_derived_59, ram_b_buff_out_7__N_128, 
            ram_b_buff_out_7__N_131, GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input \addr[1] ;
    input \addr[2] ;
    input \addr[3] ;
    input \addr[4] ;
    input \addr[5] ;
    input \addr[6] ;
    input \addr[7] ;
    input \addr[8] ;
    input \addr[9] ;
    input \addr[10] ;
    input \addr[11] ;
    input n6474;
    input n6469;
    input n6468;
    input n6467;
    input n6466;
    input n6465;
    input n6464;
    input n6463;
    input n6462;
    input n6461;
    input n6460;
    input [3:0]qspi_data_in_3__N_1;
    input [3:0]data_buff_in;
    output [7:0]ram_b_buff_out;
    input spi_clk_pos_derived_59;
    input ram_b_buff_out_7__N_128;
    input ram_b_buff_out_7__N_131;
    input GND_net;
    input VCC_net;
    
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    DP16KD mem0 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(ram_b_buff_out_7__N_128), .CSA0(GND_net), .CSA1(GND_net), 
           .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
           .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
           .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), 
           .DIB10(GND_net), .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), 
           .DIB14(GND_net), .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), 
           .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6474), 
           .ADB4(n6469), .ADB5(n6468), .ADB6(n6467), .ADB7(n6466), .ADB8(n6465), 
           .ADB9(n6464), .ADB10(n6463), .ADB11(n6462), .ADB12(n6461), 
           .ADB13(n6460), .CEB(ram_b_buff_out_7__N_131), .OCEB(VCC_net), 
           .CLKB(spi_clk_pos_derived_59), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOB0(ram_b_buff_out[0]), 
           .DOB1(ram_b_buff_out[1]), .DOB2(ram_b_buff_out[2]), .DOB3(ram_b_buff_out[3]), 
           .DOB4(ram_b_buff_out[4]), .DOB5(ram_b_buff_out[5]), .DOB6(ram_b_buff_out[6]), 
           .DOB7(ram_b_buff_out[7]));
    defparam mem0.DATA_WIDTH_A = 9;
    defparam mem0.DATA_WIDTH_B = 9;
    defparam mem0.REGMODE_A = "NOREG";
    defparam mem0.REGMODE_B = "NOREG";
    defparam mem0.RESETMODE = "SYNC";
    defparam mem0.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem0.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem0.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem0.CSDECODE_A = "0b000";
    defparam mem0.CSDECODE_B = "0b000";
    defparam mem0.GSR = "DISABLED";
    defparam mem0.INITVAL_00 = "0x00000000000000000004108E7080840088A002F50E8930682004A731E02400C800006F00A000006F";
    defparam mem0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_02 = "0x00280002170100000437080011029300200002B70000000244000000008000000000700000000070";
    defparam mem0.INITVAL_03 = "0x0602000073068820684416073000A4128B30888506020000731400105079004C0000EF1F44100213";
    defparam mem0.INITVAL_04 = "0x1D80110E93000E61F2631D80110E131D80110C930602000073068820604416073000A4128B308885";
    defparam mem0.INITVAL_05 = "0x11C911FEF710C93004F60EA630008710E931800110C130020000EB71FCE71DAE300EC1000071C023";
    defparam mem0.INITVAL_06 = "0x1FCD7136E31FCC705C2300E1100E9108690036C000E9312CB21800110E1300C91036C000C13134F1";
    defparam mem0.INITVAL_07 = "0x00EC100E41000A71E023000070EA030404000E131D80110E93000670FC631D801106131D80110E13";
    defparam mem0.INITVAL_08 = "0x00E130800510A930000302CB70200000E370100000AB71A6B80100000EB708E41100821FC671D4E3";
    defparam mem0.INITVAL_09 = "0x1FCE311E910861C0861000005100231FCF61FCE311E910861C086101128808A051A6F610C931E007";
    defparam mem0.INITVAL_0A = "0x06882180A1144230009500E63188811089300A051D026102040049500263180011688316EDD1FCF6";
    defparam mem0.INITVAL_0B = "0x1607308CA11888110E1306020000730688206045060730000800A3717ECD1808110A130602000073";
    defparam mem0.INITVAL_0C = "0x1407306045140730000800AB7180B114023000B601C63000E511A6300A85112881800116A8306006";
    defparam mem0.INITVAL_0D = "0x002000000817EE106006160731FCE601CE31804114E03060061407316EDD1808110A931008206006";
    defparam mem0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000020000008";
    defparam mem0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INIT_DATA = "STATIC";
    
endmodule
//
// Verilog Description of module \BRAM(ADDR_WIDTH=12) 
//

module \BRAM(ADDR_WIDTH=12)  (\addr[1] , \addr[2] , \addr[3] , \addr[4] , 
            \addr[5] , \addr[6] , \addr[7] , \addr[8] , \addr[9] , 
            \addr[10] , \addr[11] , n6474, n6469, n6468, n6467, 
            n6466, n6465, n6464, n6463, n6462, n6461, n6460, qspi_data_in_3__N_1, 
            data_buff_in, n6576, n6577, n6578, n6579, n6580, n6581, 
            n6582, n6583, spi_clk_pos_derived_59, n26822, ram_a_buff_out_7__N_127, 
            GND_net, VCC_net, n6568, n6569, n6570, n6571, n6572, 
            n6573, n6574, n6575, n26821, n6584, n6475) /* synthesis syn_module_defined=1 */ ;
    input \addr[1] ;
    input \addr[2] ;
    input \addr[3] ;
    input \addr[4] ;
    input \addr[5] ;
    input \addr[6] ;
    input \addr[7] ;
    input \addr[8] ;
    input \addr[9] ;
    input \addr[10] ;
    input \addr[11] ;
    input n6474;
    input n6469;
    input n6468;
    input n6467;
    input n6466;
    input n6465;
    input n6464;
    input n6463;
    input n6462;
    input n6461;
    input n6460;
    input [3:0]qspi_data_in_3__N_1;
    input [3:0]data_buff_in;
    output n6576;
    output n6577;
    output n6578;
    output n6579;
    output n6580;
    output n6581;
    output n6582;
    output n6583;
    input spi_clk_pos_derived_59;
    input n26822;
    input ram_a_buff_out_7__N_127;
    input GND_net;
    input VCC_net;
    output n6568;
    output n6569;
    output n6570;
    output n6571;
    output n6572;
    output n6573;
    output n6574;
    output n6575;
    input n26821;
    output n6584;
    input n6475;
    
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    DP16KD mem1 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(n26822), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6474), .ADB4(n6469), 
           .ADB5(n6468), .ADB6(n6467), .ADB7(n6466), .ADB8(n6465), .ADB9(n6464), 
           .ADB10(n6463), .ADB11(n6462), .ADB12(n6461), .ADB13(n6460), 
           .CEB(ram_a_buff_out_7__N_127), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6576), .DOB1(n6577), .DOB2(n6578), 
           .DOB3(n6579), .DOB4(n6580), .DOB5(n6581), .DOB6(n6582), .DOB7(n6583));
    defparam mem1.DATA_WIDTH_A = 9;
    defparam mem1.DATA_WIDTH_B = 9;
    defparam mem1.REGMODE_A = "NOREG";
    defparam mem1.REGMODE_B = "NOREG";
    defparam mem1.RESETMODE = "SYNC";
    defparam mem1.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem1.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem1.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem1.CSDECODE_A = "0b000";
    defparam mem1.CSDECODE_B = "0b000";
    defparam mem1.GSR = "DISABLED";
    defparam mem1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INIT_DATA = "STATIC";
    DP16KD mem0 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(n26821), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6474), .ADB4(n6469), 
           .ADB5(n6468), .ADB6(n6467), .ADB7(n6466), .ADB8(n6465), .ADB9(n6464), 
           .ADB10(n6463), .ADB11(n6462), .ADB12(n6461), .ADB13(n6460), 
           .CEB(ram_a_buff_out_7__N_127), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6568), .DOB1(n6569), .DOB2(n6570), 
           .DOB3(n6571), .DOB4(n6572), .DOB5(n6573), .DOB6(n6574), .DOB7(n6575));
    defparam mem0.DATA_WIDTH_A = 9;
    defparam mem0.DATA_WIDTH_B = 9;
    defparam mem0.REGMODE_A = "NOREG";
    defparam mem0.REGMODE_B = "NOREG";
    defparam mem0.RESETMODE = "SYNC";
    defparam mem0.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem0.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem0.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem0.CSDECODE_A = "0b000";
    defparam mem0.CSDECODE_B = "0b000";
    defparam mem0.GSR = "DISABLED";
    defparam mem0.INITVAL_00 = "0x00000000000000000004108E7080840088A002F50E8930682004A731E02400C800006F00A000006F";
    defparam mem0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_02 = "0x00280002170100000437080011029300200002B70000000244000000008000000000700000000070";
    defparam mem0.INITVAL_03 = "0x0602000073068820684416073000A4128B30888506020000731400105079004C0000EF1F44100213";
    defparam mem0.INITVAL_04 = "0x1D80110E93000E61F2631D80110E131D80110C930602000073068820604416073000A4128B308885";
    defparam mem0.INITVAL_05 = "0x11C911FEF710C93004F60EA630008710E931800110C130020000EB71FCE71DAE300EC1000071C023";
    defparam mem0.INITVAL_06 = "0x1FCD7136E31FCC705C2300E1100E9108690036C000E9312CB21800110E1300C91036C000C13134F1";
    defparam mem0.INITVAL_07 = "0x00EC100E41000A71E023000070EA030404000E131D80110E93000670FC631D801106131D80110E13";
    defparam mem0.INITVAL_08 = "0x00E130800510A930000302CB70200000E370100000AB71A6B80100000EB708E41100821FC671D4E3";
    defparam mem0.INITVAL_09 = "0x1FCE311E910861C0861000005100231FCF61FCE311E910861C086101128808A051A6F610C931E007";
    defparam mem0.INITVAL_0A = "0x06882180A1144230009500E63188811089300A051D026102040049500263180011688316EDD1FCF6";
    defparam mem0.INITVAL_0B = "0x1607308CA11888110E1306020000730688206045060730000800A3717ECD1808110A130602000073";
    defparam mem0.INITVAL_0C = "0x1407306045140730000800AB7180B114023000B601C63000E511A6300A85112881800116A8306006";
    defparam mem0.INITVAL_0D = "0x002000000817EE106006160731FCE601CE31804114E03060061407316EDD1808110A931008206006";
    defparam mem0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000020000008";
    defparam mem0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INIT_DATA = "STATIC";
    FD1P3AX i4302 (.D(n6475), .SP(ram_a_buff_out_7__N_127), .CK(spi_clk_pos_derived_59), 
            .Q(n6584));
    defparam i4302.GSR = "DISABLED";
    
endmodule
