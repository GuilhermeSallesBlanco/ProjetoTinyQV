// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Mon Dec 01 20:04:53 2025
//
// Verilog Description of module tinyQV_top
//

module tinyQV_top (clk, rst_n, ui_in, uo_out) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(8[8:18])
    input clk;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    input rst_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(10[20:25])
    input [7:0]ui_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    output [7:0]uo_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    wire GND_net, VCC_net, rst_n_c, ui_in_c_1, ui_in_c_0, uo_out_c_6, 
        uo_out_c_5, uo_out_c_4, uo_out_c_3, uo_out_c_2, rst_reg_n;
    wire [3:0]qspi_data_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(34[16:28])
    wire [3:0]qspi_data_oe;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(36[16:28])
    
    wire qspi_ram_a_select, qspi_ram_b_select;
    wire [27:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    wire [31:0]data_to_write;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(56[17:30])
    wire [31:0]data_from_read;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(59[16:30])
    wire [3:0]debug_rd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(75[16:24])
    
    wire debug_uart_txd;
    wire [7:6]gpio_out_sel;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(79[16:28])
    
    wire debug_register_data;
    wire [3:0]debug_rd_r;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(85[15:25])
    
    wire debug_uart_tx_start, n19951, peri_data_ready, n45, read_en;
    wire [7:0]ui_in_sync0;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(101[15:26])
    wire [7:0]ui_in_sync;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(102[15:25])
    wire [7:0]time_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(222[15:25])
    wire [3:0]qspi_data_in_3__N_1;
    wire [3:0]qspi_data_out_3__N_5;
    wire [1:0]gpio_out_sel_7__N_13;
    
    wire n44, n24126;
    wire [24:0]addr_adj_2695;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(23[16:20])
    
    wire writing, n5505;
    wire [31:0]addr_24__N_228;
    
    wire n24118, n4319, n43;
    wire [31:0]writing_N_164;
    
    wire n24114, debug_instr_valid, n42;
    wire [23:1]instr_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(56[15:25])
    wire [1:0]qv_data_write_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(64[15:30])
    
    wire n24110, rst_reg_n_adj_2691, n41, n40, next_bit, n39, uart_txd_N_2596, 
        clk_c_enable_358, n38, mem_op_increment_reg_de;
    wire [31:0]imm;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(100[16:19])
    wire [2:1]instr_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(113[15:24])
    
    wire mem_op_increment_reg, interrupt_core;
    wire [31:0]pc;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(128[17:19])
    wire [31:0]next_pc_for_core;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(129[17:33])
    wire [27:0]addr_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(131[17:25])
    wire [4:2]counter_hi;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(139[15:25])
    
    wire is_timer_addr;
    wire [3:1]instr_write_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(152[15:33])
    
    wire was_early_branch, data_ready_sync;
    wire [23:1]early_branch_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[17:34])
    
    wire n22303, n5508, clk_c_enable_420, n19950, n27106;
    wire [22:0]instr_addr_23__N_318;
    
    wire data_stall, n19923, n19949, n24806, n24804, n24803, n7164, 
        continue_txn_N_2131, data_stall_N_2158, n22999;
    wire [31:0]next_fsm_state_3__N_2499;
    
    wire n27392, n22992, n2096, clk_c_enable_426, clk_c_enable_346, 
        n2035, n2101, n2055;
    wire [1:0]cycle;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(58[15:20])
    
    wire n27083;
    wire [3:0]mul_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(138[16:23])
    
    wire n6930, n19948, n19921, n19947, n19946, n19945, clk_c_enable_367, 
        clk_c_enable_350, n808, n19944, clk_c_enable_369, n805, n19943, 
        n4057, n19942, n4577, n19941, n19940, n23908, n19939, 
        n19920, n19980, n19979, n19978, n19938, n17432, n19977, 
        n19937, n19976, n19936, n19935, n19975, n19974, n8869, 
        n19934, n19973, n19972, n19933, n19932, n19930, clk_c_enable_273, 
        n19929, n19928, n19927, n19926, n19925, n44_adj_2692, n27082, 
        n22097, n19964, n19963;
    wire [2:0]fsm_state_adj_2808;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(82[15:24])
    
    wire is_writing;
    wire [23:0]addr_adj_2809;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(84[31:35])
    
    wire is_writing_N_2331, n24802, n27081, n24561, n27080, n27365, 
        clk_c_enable_341, n1167, n27358, n27354, n27350, n24522, 
        n27342;
    wire [15:0]accum;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(104[22:27])
    wire [19:0]next_accum;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[23:33])
    wire [19:0]d_3__N_1868;
    
    wire n27335, n4307, n4309, n19962, n19961, n27127, n19960, 
        n19959, n19958, n26802, n26801, n15210, n26793, n19924, 
        n19956, n27306, n19955, n19954, n27299, n19922, n19953, 
        n19952, n27297, n27294, n27279, n27269, n26711, n24428, 
        n24376, n24314, n24312, n27241, n27237, n23276, n27393, 
        n24260, n27224, n27223, n27220, n27218, n27210, n23252, 
        n11, n27110, n3, n24140;
    
    VHI i2 (.Z(VCC_net));
    INV i24965 (.A(clk_c), .Z(clk_N_45));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    FD1S3AX debug_rd_r_i0 (.D(debug_rd[0]), .CK(clk_c), .Q(debug_rd_r[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(241[12] 243[8])
    defparam debug_rd_r_i0.GSR = "DISABLED";
    FD1S3AX rst_reg_n_53 (.D(rst_n_c), .CK(clk_N_45), .Q(rst_reg_n));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(31[12:46])
    defparam rst_reg_n_53.GSR = "DISABLED";
    \uart_tx(BIT_RATE=1000000,CLK_HZ=14000000)  i_debug_uart_tx (.debug_uart_txd(debug_uart_txd), 
            .clk_c(clk_c), .clk_c_enable_341(clk_c_enable_341), .clk_c_enable_426(clk_c_enable_426), 
            .n27294(n27294), .debug_uart_tx_start(debug_uart_tx_start), 
            .\data_to_write[4] (data_to_write[4]), .\data_to_write[5] (data_to_write[5]), 
            .\data_to_write[6] (data_to_write[6]), .rst_reg_n(rst_reg_n), 
            .n27210(n27210), .next_bit(next_bit), .uart_txd_N_2596(uart_txd_N_2596), 
            .\data_to_write[2] (data_to_write[2]), .\data_to_write[1] (data_to_write[1]), 
            .\data_to_write[0] (data_to_write[0]), .\data_to_write[7] (data_to_write[7]), 
            .\data_to_write[3] (data_to_write[3])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(213[67] 220[6])
    \peripherals_min(CLOCK_MHZ=14)  i_peripherals (.peri_data_ready(peri_data_ready), 
            .clk_c(clk_c), .clk_c_enable_341(clk_c_enable_341), .read_en(read_en)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(161[46] 180[6])
    FD1P3AX gpio_out_sel_i7 (.D(gpio_out_sel_7__N_13[1]), .SP(clk_c_enable_420), 
            .CK(clk_c), .Q(gpio_out_sel[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(204[12] 211[8])
    defparam gpio_out_sel_i7.GSR = "DISABLED";
    GSR GSR_INST (.GSR(n27335));
    IB ui_in_pad_0 (.I(ui_in[0]), .O(ui_in_c_0));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_1 (.I(ui_in[1]), .O(ui_in_c_1));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB rst_n_pad (.I(rst_n), .O(rst_n_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(10[20:25])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    OB uo_out_pad_0 (.I(GND_net), .O(uo_out[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_1 (.I(GND_net), .O(uo_out[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    CCU2C time_count_3234_add_4_5 (.A0(time_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19944), .COUT(n19945), .S0(n42), .S1(n41));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234_add_4_5.INIT0 = 16'haaa0;
    defparam time_count_3234_add_4_5.INIT1 = 16'haaa0;
    defparam time_count_3234_add_4_5.INJECT1_0 = "NO";
    defparam time_count_3234_add_4_5.INJECT1_1 = "NO";
    OB uo_out_pad_2 (.I(uo_out_c_2), .O(uo_out[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    CCU2C time_count_3234_add_4_3 (.A0(time_count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19943), .COUT(n19944), .S0(n44), .S1(n43));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234_add_4_3.INIT0 = 16'haaa0;
    defparam time_count_3234_add_4_3.INIT1 = 16'haaa0;
    defparam time_count_3234_add_4_3.INJECT1_0 = "NO";
    defparam time_count_3234_add_4_3.INJECT1_1 = "NO";
    LUT4 i3356_4_lut_then_3_lut (.A(n27218), .B(counter_hi[4]), .C(counter_hi[3]), 
         .Z(n27393)) /* synthesis lut_function=(A+!((C)+!B)) */ ;
    defparam i3356_4_lut_then_3_lut.init = 16'haeae;
    LUT4 i3356_4_lut_else_3_lut (.A(n27218), .B(counter_hi[4]), .C(counter_hi[3]), 
         .D(counter_hi[2]), .Z(n27392)) /* synthesis lut_function=(A+!((C+!(D))+!B)) */ ;
    defparam i3356_4_lut_else_3_lut.init = 16'haeaa;
    LUT4 i12467_2_lut (.A(qspi_data_in[3]), .B(rst_reg_n), .Z(qspi_data_out_3__N_5[3])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(127[22:56])
    defparam i12467_2_lut.init = 16'h8888;
    CCU2C time_count_3234_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n19943), .S1(n45));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234_add_4_1.INIT0 = 16'h0000;
    defparam time_count_3234_add_4_1.INIT1 = 16'h555f;
    defparam time_count_3234_add_4_1.INJECT1_0 = "NO";
    defparam time_count_3234_add_4_1.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync_i2 (.D(ui_in_sync0[1]), .CK(clk_c), .Q(ui_in_sync[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i2.GSR = "DISABLED";
    LUT4 i22463_3_lut (.A(data_stall), .B(data_stall_N_2158), .C(continue_txn_N_2131), 
         .Z(n24806)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam i22463_3_lut.init = 16'hcece;
    LUT4 n5057_bdd_3_lut_24158_4_lut (.A(n27224), .B(n17432), .C(gpio_out_sel[7]), 
         .D(data_from_read[2]), .Z(n26793)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (C+(D))) */ ;
    defparam n5057_bdd_3_lut_24158_4_lut.init = 16'hffd0;
    LUT4 i23651_2_lut (.A(rst_reg_n), .B(n805), .Z(n15210)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i23651_2_lut.init = 16'h1111;
    FD1S3AX ui_in_sync0_i2 (.D(ui_in_c_1), .CK(clk_c), .Q(ui_in_sync0[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i2.GSR = "DISABLED";
    CCU2C _add_1_4407_add_4_21 (.A0(early_branch_addr[21]), .B0(was_early_branch), 
          .C0(pc[21]), .D0(VCC_net), .A1(early_branch_addr[22]), .B1(was_early_branch), 
          .C1(pc[22]), .D1(VCC_net), .CIN(n19929), .COUT(n19930), .S0(instr_addr_23__N_318[20]), 
          .S1(instr_addr_23__N_318[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_21.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_21.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_19 (.A0(early_branch_addr[19]), .B0(was_early_branch), 
          .C0(pc[19]), .D0(VCC_net), .A1(early_branch_addr[20]), .B1(was_early_branch), 
          .C1(pc[20]), .D1(VCC_net), .CIN(n19928), .COUT(n19929), .S0(instr_addr_23__N_318[18]), 
          .S1(instr_addr_23__N_318[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_19.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_19.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_17 (.A0(early_branch_addr[17]), .B0(was_early_branch), 
          .C0(pc[17]), .D0(VCC_net), .A1(early_branch_addr[18]), .B1(was_early_branch), 
          .C1(pc[18]), .D1(VCC_net), .CIN(n19927), .COUT(n19928), .S0(instr_addr_23__N_318[16]), 
          .S1(instr_addr_23__N_318[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_17.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_17.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_15 (.A0(early_branch_addr[15]), .B0(was_early_branch), 
          .C0(pc[15]), .D0(VCC_net), .A1(early_branch_addr[16]), .B1(was_early_branch), 
          .C1(pc[16]), .D1(VCC_net), .CIN(n19926), .COUT(n19927), .S0(instr_addr_23__N_318[14]), 
          .S1(instr_addr_23__N_318[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_15.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_15.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_13 (.A0(early_branch_addr[13]), .B0(was_early_branch), 
          .C0(pc[13]), .D0(VCC_net), .A1(early_branch_addr[14]), .B1(was_early_branch), 
          .C1(pc[14]), .D1(VCC_net), .CIN(n19925), .COUT(n19926), .S0(instr_addr_23__N_318[12]), 
          .S1(instr_addr_23__N_318[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_13.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_13.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_11 (.A0(early_branch_addr[11]), .B0(was_early_branch), 
          .C0(pc[11]), .D0(VCC_net), .A1(early_branch_addr[12]), .B1(was_early_branch), 
          .C1(pc[12]), .D1(VCC_net), .CIN(n19924), .COUT(n19925), .S0(instr_addr_23__N_318[10]), 
          .S1(instr_addr_23__N_318[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_11.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_11.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_9 (.A0(early_branch_addr[9]), .B0(was_early_branch), 
          .C0(pc[9]), .D0(VCC_net), .A1(early_branch_addr[10]), .B1(was_early_branch), 
          .C1(pc[10]), .D1(VCC_net), .CIN(n19923), .COUT(n19924), .S0(instr_addr_23__N_318[8]), 
          .S1(instr_addr_23__N_318[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_9.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_9.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_7 (.A0(early_branch_addr[7]), .B0(was_early_branch), 
          .C0(pc[7]), .D0(VCC_net), .A1(early_branch_addr[8]), .B1(was_early_branch), 
          .C1(pc[8]), .D1(VCC_net), .CIN(n19922), .COUT(n19923), .S0(instr_addr_23__N_318[6]), 
          .S1(instr_addr_23__N_318[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_7.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_7.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_3 (.A0(pc[3]), .B0(was_early_branch), .C0(early_branch_addr[3]), 
          .D0(instr_write_offset[3]), .A1(early_branch_addr[4]), .B1(was_early_branch), 
          .C1(pc[4]), .D1(VCC_net), .CIN(n19920), .COUT(n19921), .S0(instr_addr_23__N_318[2]), 
          .S1(instr_addr_23__N_318[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_4407_add_4_3.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_3.INJECT1_1 = "NO";
    FD1P3AX debug_register_data_58 (.D(n7164), .SP(clk_c_enable_273), .CK(clk_c), 
            .Q(debug_register_data));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(234[12] 239[8])
    defparam debug_register_data_58.GSR = "DISABLED";
    OB uo_out_pad_4 (.I(uo_out_c_4), .O(uo_out[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    FD1S3AX debug_rd_r_i3 (.D(debug_rd[3]), .CK(clk_c), .Q(debug_rd_r[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(241[12] 243[8])
    defparam debug_rd_r_i3.GSR = "DISABLED";
    tinyQV i_tinyqv (.rst_reg_n_adj_15(rst_reg_n_adj_2691), .clk_c(clk_c), 
           .rst_reg_n(rst_reg_n), .\data_from_read[2] (data_from_read[2]), 
           .n27358(n27358), .\addr[2] (addr[2]), .n22303(n22303), .read_en(read_en), 
           .n17432(n17432), .\addr[5] (addr[5]), .n24260(n24260), .n24118(n24118), 
           .n27269(n27269), .counter_hi({counter_hi}), .peri_data_ready(peri_data_ready), 
           .clk_c_enable_341(clk_c_enable_341), .\instr_addr_23__N_318[0] (instr_addr_23__N_318[0]), 
           .\instr_addr_23__N_318[18] (instr_addr_23__N_318[18]), .\instr_addr_23__N_318[14] (instr_addr_23__N_318[14]), 
           .\instr_addr_23__N_318[15] (instr_addr_23__N_318[15]), .\instr_addr_23__N_318[16] (instr_addr_23__N_318[16]), 
           .\instr_addr_23__N_318[17] (instr_addr_23__N_318[17]), .\instr_addr_23__N_318[6] (instr_addr_23__N_318[6]), 
           .\addr[7] (addr[7]), .\instr_addr_23__N_318[5] (instr_addr_23__N_318[5]), 
           .\addr[6] (addr[6]), .\instr_addr_23__N_318[7] (instr_addr_23__N_318[7]), 
           .\addr[8] (addr[8]), .\instr_addr_23__N_318[3] (instr_addr_23__N_318[3]), 
           .\addr[4] (addr[4]), .\instr_addr_23__N_318[10] (instr_addr_23__N_318[10]), 
           .data_stall(data_stall), .\instr_addr_23__N_318[9] (instr_addr_23__N_318[9]), 
           .\addr[10] (addr[10]), .\instr_addr_23__N_318[11] (instr_addr_23__N_318[11]), 
           .\instr_addr_23__N_318[8] (instr_addr_23__N_318[8]), .\addr[9] (addr[9]), 
           .\instr_addr[1] (instr_addr[1]), .\addr[1] (addr[1]), .\instr_addr_23__N_318[12] (instr_addr_23__N_318[12]), 
           .\instr_addr_23__N_318[22] (instr_addr_23__N_318[22]), .\instr_addr_23__N_318[13] (instr_addr_23__N_318[13]), 
           .\instr_addr_23__N_318[4] (instr_addr_23__N_318[4]), .\instr_addr_23__N_318[19] (instr_addr_23__N_318[19]), 
           .\instr_addr_23__N_318[20] (instr_addr_23__N_318[20]), .\instr_addr_23__N_318[21] (instr_addr_23__N_318[21]), 
           .n27081(n27081), .is_writing_N_2331(is_writing_N_2331), .n27299(n27299), 
           .\data_to_write[7] (data_to_write[7]), .\data_to_write[6] (data_to_write[6]), 
           .continue_txn_N_2131(continue_txn_N_2131), .data_stall_N_2158(data_stall_N_2158), 
           .\data_to_write[5] (data_to_write[5]), .\pc[1] (pc[1]), .\pc[2] (pc[2]), 
           .n24806(n24806), .\data_to_write[4] (data_to_write[4]), .qv_data_write_n({qv_data_write_n}), 
           .\data_to_write[0] (data_to_write[0]), .\data_to_write[3] (data_to_write[3]), 
           .\data_to_write[2] (data_to_write[2]), .\data_to_write[1] (data_to_write[1]), 
           .n27082(n27082), .\addr[0] (addr[0]), .is_writing(is_writing), 
           .\instr_addr_23__N_318[2] (instr_addr_23__N_318[2]), .\addr[3] (addr[3]), 
           .n6930(n6930), .\writing_N_164[3] (writing_N_164[3]), .n27083(n27083), 
           .qspi_ram_b_select(qspi_ram_b_select), .\qspi_data_out_3__N_5[0] (qspi_data_out_3__N_5[0]), 
           .qspi_ram_a_select(qspi_ram_a_select), .n24802(n24802), .qspi_data_in({qspi_data_in}), 
           .\fsm_state[0] (fsm_state_adj_2808[0]), .n23276(n23276), .clk_c_enable_358(clk_c_enable_358), 
           .clk_c_enable_369(clk_c_enable_369), .n23252(n23252), .clk_N_45(clk_N_45), 
           .\qspi_data_out_3__N_5[2] (qspi_data_out_3__N_5[2]), .n4319(n4319), 
           .n4307(n4307), .\qspi_data_oe[3] (qspi_data_oe[3]), .clk_c_enable_346(clk_c_enable_346), 
           .n27080(n27080), .\qspi_data_out_3__N_5[3] (qspi_data_out_3__N_5[3]), 
           .\addr[20] (addr_adj_2809[20]), .\addr[22] (addr_adj_2809[22]), 
           .spi_clk_pos_derived_59(spi_clk_pos_derived_59), .qspi_clk_N_56(qspi_clk_N_56), 
           .next_bit(next_bit), .n27210(n27210), .uart_txd_N_2596(uart_txd_N_2596), 
           .clk_c_enable_426(clk_c_enable_426), .n24376(n24376), .n44(n44_adj_2692), 
           .clk_c_enable_273(clk_c_enable_273), .n805(n805), .clk_c_enable_420(clk_c_enable_420), 
           .n27365(n27365), .n22097(n22097), .n4309(n4309), .n26711(n26711), 
           .n5508(n5508), .n5505(n5505), .n22992(n22992), .\instr_len[2] (instr_len[2]), 
           .VCC_net(VCC_net), .interrupt_core(interrupt_core), .n2055(n2055), 
           .debug_instr_valid(debug_instr_valid), .was_early_branch(was_early_branch), 
           .n2035(n2035), .\pc[10] (pc[10]), .n27106(n27106), .data_ready_sync(data_ready_sync), 
           .n2096(n2096), .n2101(n2101), .\imm[23] (imm[23]), .n4057(n4057), 
           .n26793(n26793), .\imm[22] (imm[22]), .\imm[1] (imm[1]), .\imm[10] (imm[10]), 
           .\imm[21] (imm[21]), .\imm[20] (imm[20]), .\imm[6] (imm[6]), 
           .\imm[19] (imm[19]), .\imm[18] (imm[18]), .\imm[17] (imm[17]), 
           .\imm[16] (imm[16]), .\imm[15] (imm[15]), .\imm[14] (imm[14]), 
           .\imm[13] (imm[13]), .\imm[12] (imm[12]), .\imm[11] (imm[11]), 
           .\imm[9] (imm[9]), .\imm[8] (imm[8]), .\imm[7] (imm[7]), .\imm[5] (imm[5]), 
           .\imm[4] (imm[4]), .\imm[3] (imm[3]), .\imm[2] (imm[2]), .is_timer_addr(is_timer_addr), 
           .n27354(n27354), .n27342(n27342), .\addr_out[1] (addr_out[1]), 
           .\instr_write_offset[3] (instr_write_offset[3]), .n27297(n27297), 
           .mem_op_increment_reg(mem_op_increment_reg), .n24804(n24804), 
           .\pc[23] (pc[23]), .\next_pc_for_core[6] (next_pc_for_core[6]), 
           .\next_pc_for_core[4] (next_pc_for_core[4]), .\next_pc_for_core[9] (next_pc_for_core[9]), 
           .\next_pc_for_core[13] (next_pc_for_core[13]), .\pc[8] (pc[8]), 
           .\pc[12] (pc[12]), .\next_pc_for_core[3] (next_pc_for_core[3]), 
           .\next_pc_for_core[5] (next_pc_for_core[5]), .\pc[4] (pc[4]), 
           .\next_pc_for_core[7] (next_pc_for_core[7]), .\next_pc_for_core[8] (next_pc_for_core[8]), 
           .\next_pc_for_core[10] (next_pc_for_core[10]), .\next_pc_for_core[12] (next_pc_for_core[12]), 
           .\next_pc_for_core[11] (next_pc_for_core[11]), .\next_pc_for_core[14] (next_pc_for_core[14]), 
           .\next_pc_for_core[15] (next_pc_for_core[15]), .\next_pc_for_core[16] (next_pc_for_core[16]), 
           .\next_pc_for_core[17] (next_pc_for_core[17]), .\next_pc_for_core[18] (next_pc_for_core[18]), 
           .\next_pc_for_core[19] (next_pc_for_core[19]), .\next_pc_for_core[20] (next_pc_for_core[20]), 
           .\next_pc_for_core[21] (next_pc_for_core[21]), .\next_pc_for_core[22] (next_pc_for_core[22]), 
           .\next_pc_for_core[23] (next_pc_for_core[23]), .\pc[22] (pc[22]), 
           .\pc[21] (pc[21]), .\pc[20] (pc[20]), .\pc[19] (pc[19]), .\pc[18] (pc[18]), 
           .\pc[17] (pc[17]), .\pc[16] (pc[16]), .\pc[15] (pc[15]), .\pc[14] (pc[14]), 
           .\pc[13] (pc[13]), .\pc[11] (pc[11]), .\pc[9] (pc[9]), .\pc[7] (pc[7]), 
           .\pc[6] (pc[6]), .\pc[5] (pc[5]), .\pc[3] (pc[3]), .n27127(n27127), 
           .n27110(n27110), .cycle({cycle}), .n27350(n27350), .\early_branch_addr[3] (early_branch_addr[3]), 
           .\early_branch_addr[6] (early_branch_addr[6]), .\early_branch_addr[2] (early_branch_addr[2]), 
           .\early_branch_addr[5] (early_branch_addr[5]), .\early_branch_addr[4] (early_branch_addr[4]), 
           .\early_branch_addr[7] (early_branch_addr[7]), .\early_branch_addr[8] (early_branch_addr[8]), 
           .\early_branch_addr[9] (early_branch_addr[9]), .\early_branch_addr[10] (early_branch_addr[10]), 
           .\early_branch_addr[11] (early_branch_addr[11]), .\early_branch_addr[12] (early_branch_addr[12]), 
           .\early_branch_addr[13] (early_branch_addr[13]), .\early_branch_addr[14] (early_branch_addr[14]), 
           .\early_branch_addr[15] (early_branch_addr[15]), .\early_branch_addr[16] (early_branch_addr[16]), 
           .\early_branch_addr[17] (early_branch_addr[17]), .\early_branch_addr[18] (early_branch_addr[18]), 
           .\early_branch_addr[19] (early_branch_addr[19]), .\early_branch_addr[20] (early_branch_addr[20]), 
           .\early_branch_addr[21] (early_branch_addr[21]), .\early_branch_addr[22] (early_branch_addr[22]), 
           .\early_branch_addr[23] (early_branch_addr[23]), .n27294(n27294), 
           .n27306(n27306), .\data_from_read[6] (data_from_read[6]), .n24126(n24126), 
           .n27241(n27241), .n8869(n8869), .n27279(n27279), .n23908(n23908), 
           .n27220(n27220), .mem_op_increment_reg_de(mem_op_increment_reg_de), 
           .n27218(n27218), .\next_fsm_state_3__N_2499[3] (next_fsm_state_3__N_2499[3]), 
           .clk_c_enable_350(clk_c_enable_350), .clk_c_enable_367(clk_c_enable_367), 
           .\mul_out[2] (mul_out[2]), .\mul_out[3] (mul_out[3]), .\mul_out[1] (mul_out[1]), 
           .\ui_in_sync[1] (ui_in_sync[1]), .n1167(n1167), .debug_rd({debug_rd}), 
           .accum({accum}), .d_3__N_1868({d_3__N_1868}), .n4577(n4577), 
           .n26802(n26802), .n27223(n27223), .\next_accum[5] (next_accum[5]), 
           .\next_accum[6] (next_accum[6]), .\next_accum[7] (next_accum[7]), 
           .GND_net(GND_net), .\next_accum[8] (next_accum[8]), .\next_accum[9] (next_accum[9]), 
           .\next_accum[10] (next_accum[10]), .\next_accum[11] (next_accum[11]), 
           .\next_accum[12] (next_accum[12]), .\next_accum[13] (next_accum[13]), 
           .\next_accum[14] (next_accum[14]), .\next_accum[15] (next_accum[15]), 
           .\next_accum[16] (next_accum[16]), .\next_accum[17] (next_accum[17]), 
           .\next_accum[18] (next_accum[18]), .\next_accum[19] (next_accum[19]), 
           .\next_accum[4] (next_accum[4])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(111[12] 150[6])
    FD1S3AX debug_rd_r_i2 (.D(debug_rd[2]), .CK(clk_c), .Q(debug_rd_r[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(241[12] 243[8])
    defparam debug_rd_r_i2.GSR = "DISABLED";
    FD1S3AX ui_in_sync0_i1 (.D(ui_in_c_0), .CK(clk_c), .Q(ui_in_sync0[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i1.GSR = "DISABLED";
    FD1S3AX debug_rd_r_i1 (.D(debug_rd[1]), .CK(clk_c), .Q(debug_rd_r[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(241[12] 243[8])
    defparam debug_rd_r_i1.GSR = "DISABLED";
    CCU2C _add_1_4402_add_4_24 (.A0(imm[23]), .B0(pc[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19942), .S0(early_branch_addr[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_24.INIT1 = 16'h0000;
    defparam _add_1_4402_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_24.INJECT1_1 = "NO";
    LUT4 i12604_3_lut_4_lut (.A(n27224), .B(n17432), .C(data_from_read[2]), 
         .D(gpio_out_sel[6]), .Z(data_from_read[6])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C+(D))) */ ;
    defparam i12604_3_lut_4_lut.init = 16'hfdf0;
    OB uo_out_pad_5 (.I(uo_out_c_5), .O(uo_out[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_6 (.I(uo_out_c_6), .O(uo_out[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    FD1S3IX time_count_3234__i0 (.D(n45), .CK(clk_c), .CD(n808), .Q(time_count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234__i0.GSR = "DISABLED";
    OB uo_out_pad_3 (.I(uo_out_c_3), .O(uo_out[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_7 (.I(GND_net), .O(uo_out[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    CCU2C _add_1_4402_add_4_22 (.A0(imm[21]), .B0(pc[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[22]), .B1(pc[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19941), .COUT(n19942), .S0(early_branch_addr[21]), .S1(early_branch_addr[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_4402_add_4_20 (.A0(imm[19]), .B0(pc[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[20]), .B1(pc[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19940), .COUT(n19941), .S0(early_branch_addr[19]), .S1(early_branch_addr[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_20 (.A0(d_3__N_1868[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_3__N_1868[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19980), .S0(next_accum[18]), .S1(next_accum[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_add_4_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_add_4_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_18 (.A0(d_3__N_1868[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_3__N_1868[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19979), .COUT(n19980), .S0(next_accum[16]), 
          .S1(next_accum[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_add_4_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_add_4_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_16 (.A0(accum[14]), .B0(d_3__N_1868[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[15]), .B1(d_3__N_1868[15]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19978), .COUT(n19979), .S0(next_accum[14]), 
          .S1(next_accum[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_4402_add_4_18 (.A0(imm[17]), .B0(pc[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[18]), .B1(pc[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19939), .COUT(n19940), .S0(early_branch_addr[17]), .S1(early_branch_addr[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_4402_add_4_16 (.A0(imm[15]), .B0(pc[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[16]), .B1(pc[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19938), .COUT(n19939), .S0(early_branch_addr[15]), .S1(early_branch_addr[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_14 (.A0(accum[12]), .B0(d_3__N_1868[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[13]), .B1(d_3__N_1868[13]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19977), .COUT(n19978), .S0(next_accum[12]), 
          .S1(next_accum[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_4402_add_4_14 (.A0(imm[13]), .B0(pc[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[14]), .B1(pc[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19937), .COUT(n19938), .S0(early_branch_addr[13]), .S1(early_branch_addr[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_4402_add_4_12 (.A0(imm[11]), .B0(pc[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[12]), .B1(pc[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19936), .COUT(n19937), .S0(early_branch_addr[11]), .S1(early_branch_addr[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_12 (.A0(accum[10]), .B0(d_3__N_1868[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[11]), .B1(d_3__N_1868[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19976), .COUT(n19977), .S0(next_accum[10]), 
          .S1(next_accum[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_12.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(addr_adj_2809[20]), .B(n22097), .C(n4309), .D(fsm_state_adj_2808[0]), 
         .Z(qspi_data_in_3__N_1[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(43[23:51])
    defparam i1_4_lut.init = 16'hc088;
    CCU2C _add_1_4402_add_4_10 (.A0(imm[9]), .B0(pc[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[10]), .B1(pc[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19935), .COUT(n19936), .S0(early_branch_addr[9]), .S1(early_branch_addr[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_10 (.A0(accum[8]), .B0(d_3__N_1868[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[9]), .B1(d_3__N_1868[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19975), .COUT(n19976), .S0(next_accum[8]), 
          .S1(next_accum[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_4402_add_4_8 (.A0(imm[7]), .B0(pc[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[8]), .B1(pc[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19934), .COUT(n19935), .S0(early_branch_addr[7]), .S1(early_branch_addr[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_8 (.A0(accum[6]), .B0(d_3__N_1868[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[7]), .B1(d_3__N_1868[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19974), .COUT(n19975), .S0(next_accum[6]), 
          .S1(next_accum[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_8.INJECT1_1 = "NO";
    LUT4 qspi_data_out_3__I_0_i2_3_lut (.A(n4319), .B(qspi_data_oe[3]), 
         .C(n27365), .Z(qspi_data_in_3__N_1[1])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(43[23:51])
    defparam qspi_data_out_3__I_0_i2_3_lut.init = 16'h8c8c;
    LUT4 i1_4_lut_adj_490 (.A(addr_adj_2809[22]), .B(n22097), .C(n4307), 
         .D(fsm_state_adj_2808[0]), .Z(qspi_data_in_3__N_1[2])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(43[23:51])
    defparam i1_4_lut_adj_490.init = 16'hc088;
    LUT4 qspi_data_out_3__I_0_i4_3_lut (.A(n26711), .B(qspi_data_oe[3]), 
         .C(n27365), .Z(qspi_data_in_3__N_1[3])) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(43[23:51])
    defparam qspi_data_out_3__I_0_i4_3_lut.init = 16'h8c8c;
    LUT4 i1_2_lut (.A(addr[4]), .B(addr[5]), .Z(n24140)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_adj_491 (.A(addr[2]), .B(addr[3]), .Z(n3)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_2_lut_adj_491.init = 16'h8888;
    CCU2C _add_1_add_4_add_4_6 (.A0(accum[4]), .B0(d_3__N_1868[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[5]), .B1(d_3__N_1868[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19973), .COUT(n19974), .S0(next_accum[4]), 
          .S1(next_accum[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_4 (.A0(accum[2]), .B0(d_3__N_1868[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[3]), .B1(d_3__N_1868[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19972), .COUT(n19973), .S0(mul_out[2]), 
          .S1(mul_out[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_4402_add_4_6 (.A0(imm[5]), .B0(pc[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[6]), .B1(pc[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19933), .COUT(n19934), .S0(early_branch_addr[5]), .S1(early_branch_addr[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_5 (.A0(early_branch_addr[5]), .B0(was_early_branch), 
          .C0(pc[5]), .D0(VCC_net), .A1(early_branch_addr[6]), .B1(was_early_branch), 
          .C1(pc[6]), .D1(VCC_net), .CIN(n19921), .COUT(n19922), .S0(instr_addr_23__N_318[4]), 
          .S1(instr_addr_23__N_318[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_5.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_5.INIT1 = 16'hb8b8;
    defparam _add_1_4407_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_4407_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(was_early_branch), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n19920));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_4407_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_4407_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_4402_add_4_4 (.A0(imm[3]), .B0(pc[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[4]), .B1(pc[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19932), .COUT(n19933), .S0(early_branch_addr[3]), .S1(early_branch_addr[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_4402_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_4402_add_4_2 (.A0(imm[1]), .B0(pc[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[2]), .B1(pc[2]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n19932), .S1(early_branch_addr[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4402_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_4402_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_4402_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_4402_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_2 (.A0(accum[0]), .B0(d_3__N_1868[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[1]), .B1(d_3__N_1868[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n19972), .S1(mul_out[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_add_4_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_2.INJECT1_1 = "NO";
    LUT4 i1340_4_lut (.A(pc[2]), .B(n2096), .C(debug_instr_valid), .D(pc[1]), 
         .Z(n2055)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i1340_4_lut.init = 16'hcac0;
    FD1P3IX gpio_out_sel_i6 (.D(data_to_write[6]), .SP(clk_c_enable_420), 
            .CD(n15210), .CK(clk_c), .Q(gpio_out_sel[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(204[12] 211[8])
    defparam gpio_out_sel_i6.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_492 (.A(n27237), .B(n22303), .C(n11), .D(n24260), 
         .Z(debug_uart_tx_start)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_4_lut_adj_492.init = 16'h1000;
    LUT4 i1_2_lut_adj_493 (.A(n17432), .B(addr[5]), .Z(n11)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_2_lut_adj_493.init = 16'hbbbb;
    FD1S3IX time_count_3234__i1 (.D(n44), .CK(clk_c), .CD(n808), .Q(time_count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234__i1.GSR = "DISABLED";
    FD1S3IX time_count_3234__i2 (.D(n43), .CK(clk_c), .CD(n808), .Q(time_count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234__i2.GSR = "DISABLED";
    FD1S3IX time_count_3234__i3 (.D(n42), .CK(clk_c), .CD(n808), .Q(time_count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234__i3.GSR = "DISABLED";
    FD1S3IX time_count_3234__i4 (.D(n41), .CK(clk_c), .CD(n808), .Q(time_count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234__i4.GSR = "DISABLED";
    FD1S3IX time_count_3234__i5 (.D(n40), .CK(clk_c), .CD(n808), .Q(time_count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234__i5.GSR = "DISABLED";
    FD1S3IX time_count_3234__i6 (.D(n39), .CK(clk_c), .CD(n808), .Q(time_count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234__i6.GSR = "DISABLED";
    FD1S3IX time_count_3234__i7 (.D(n38), .CK(clk_c), .CD(n808), .Q(time_count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234__i7.GSR = "DISABLED";
    CCU2C _add_1_4407_add_4_23 (.A0(early_branch_addr[23]), .B0(was_early_branch), 
          .C0(pc[23]), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19930), .S0(instr_addr_23__N_318[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4407_add_4_23.INIT0 = 16'hb8b8;
    defparam _add_1_4407_add_4_23.INIT1 = 16'h0000;
    defparam _add_1_4407_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_4407_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_4396_add_4_15 (.A0(addr_adj_2695[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_2695[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19964), .S0(addr_24__N_228[13]), .S1(addr_24__N_228[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_4396_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_4396_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_4396_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_4396_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_4396_add_4_13 (.A0(addr_adj_2695[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_2695[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19963), .COUT(n19964), .S0(addr_24__N_228[11]), 
          .S1(addr_24__N_228[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_4396_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_4396_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_4396_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_4396_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_4396_add_4_11 (.A0(addr_adj_2695[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_2695[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19962), .COUT(n19963), .S0(addr_24__N_228[9]), 
          .S1(addr_24__N_228[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_4396_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_4396_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_4396_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_4396_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_4396_add_4_9 (.A0(addr_adj_2695[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_2695[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19961), .COUT(n19962), .S0(addr_24__N_228[7]), 
          .S1(addr_24__N_228[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_4396_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_4396_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_4396_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_4396_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_4396_add_4_7 (.A0(addr_adj_2695[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_2695[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19960), .COUT(n19961), .S0(addr_24__N_228[5]), 
          .S1(addr_24__N_228[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_4396_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_4396_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_4396_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_4396_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_4396_add_4_5 (.A0(addr_adj_2695[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_2695[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19959), .COUT(n19960), .S0(addr_24__N_228[3]), 
          .S1(addr_24__N_228[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_4396_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_4396_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_4396_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_4396_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_4396_add_4_3 (.A0(addr_adj_2695[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_2695[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19958), .COUT(n19959), .S0(addr_24__N_228[1]), 
          .S1(addr_24__N_228[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_4396_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_4396_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_4396_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_4396_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_4396_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr_adj_2695[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n19958), .S1(addr_24__N_228[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_4396_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_4396_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_4396_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_4396_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_4399_add_4_21 (.A0(pc[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[23]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19956), .S0(next_pc_for_core[22]), .S1(next_pc_for_core[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_21.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync_i1 (.D(ui_in_sync0[0]), .CK(clk_c), .Q(next_fsm_state_3__N_2499[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i1.GSR = "DISABLED";
    VLO i1 (.Z(GND_net));
    LUT4 instr_addr_23__I_0_i1_3_lut_4_lut (.A(imm[1]), .B(pc[1]), .C(was_early_branch), 
         .D(instr_addr_23__N_318[0]), .Z(instr_addr[1])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam instr_addr_23__I_0_i1_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_2792_i1_3_lut_4_lut (.A(imm[1]), .B(pc[1]), .C(n27350), .D(addr_out[1]), 
         .Z(n4577)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_2792_i1_3_lut_4_lut.init = 16'h6f60;
    CCU2C _add_1_4399_add_4_19 (.A0(pc[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[21]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19955), .COUT(n19956), .S0(next_pc_for_core[20]), .S1(next_pc_for_core[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_19.INJECT1_1 = "NO";
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    CCU2C _add_1_4399_add_4_17 (.A0(pc[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[19]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19954), .COUT(n19955), .S0(next_pc_for_core[18]), .S1(next_pc_for_core[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_4399_add_4_15 (.A0(pc[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19953), .COUT(n19954), .S0(next_pc_for_core[16]), .S1(next_pc_for_core[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_4399_add_4_13 (.A0(pc[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[15]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19952), .COUT(n19953), .S0(next_pc_for_core[14]), .S1(next_pc_for_core[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_13.INJECT1_1 = "NO";
    LUT4 i12327_2_lut_rep_733 (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .Z(n27358)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12327_2_lut_rep_733.init = 16'h8888;
    LUT4 i1_2_lut_rep_595_3_lut_4_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(addr[2]), .D(is_timer_addr), .Z(n27220)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;
    defparam i1_2_lut_rep_595_3_lut_4_lut.init = 16'h0700;
    LUT4 i1_2_lut_rep_616_3_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(is_timer_addr), .Z(n27241)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_rep_616_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_3_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(data_ready_sync), .Z(n24126)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_598_3_lut_4_lut (.A(qv_data_write_n[0]), .B(qv_data_write_n[1]), 
         .C(addr[2]), .D(is_timer_addr), .Z(n27223)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam i1_2_lut_rep_598_3_lut_4_lut.init = 16'h7000;
    CCU2C _add_1_4399_add_4_11 (.A0(pc[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[13]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19951), .COUT(n19952), .S0(next_pc_for_core[12]), .S1(next_pc_for_core[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_4399_add_4_9 (.A0(pc[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[11]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19950), .COUT(n19951), .S0(next_pc_for_core[10]), .S1(next_pc_for_core[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_4399_add_4_7 (.A0(pc[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[9]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19949), .COUT(n19950), .S0(next_pc_for_core[8]), .S1(next_pc_for_core[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_4399_add_4_5 (.A0(pc[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[7]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19948), .COUT(n19949), .S0(next_pc_for_core[6]), .S1(next_pc_for_core[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_5.INJECT1_1 = "NO";
    LUT4 mux_34_i2_3_lut (.A(ui_in_c_0), .B(data_to_write[7]), .C(n805), 
         .Z(gpio_out_sel_7__N_13[1])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(209[13:93])
    defparam mux_34_i2_3_lut.init = 16'hc5c5;
    CCU2C _add_1_4399_add_4_3 (.A0(pc[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[5]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n19947), .COUT(n19948), .S0(next_pc_for_core[4]), .S1(next_pc_for_core[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_4399_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_4399_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_494 (.A(n27224), .B(n27269), .C(n24522), .D(addr[2]), 
         .Z(n805)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_494.init = 16'h0100;
    LUT4 i22245_3_lut (.A(n24118), .B(n17432), .C(addr[3]), .Z(n24522)) /* synthesis lut_function=(A (B)+!A (B+!(C))) */ ;
    defparam i22245_3_lut.init = 16'hcdcd;
    CCU2C _add_1_4399_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[3]), .B1(n27354), .C1(instr_len[2]), 
          .D1(pc[2]), .COUT(n19947), .S1(next_pc_for_core[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4399_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_4399_add_4_1.INIT1 = 16'h566a;
    defparam _add_1_4399_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_4399_add_4_1.INJECT1_1 = "NO";
    CCU2C time_count_3234_add_4_9 (.A0(time_count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19946), .S0(n38));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234_add_4_9.INIT0 = 16'haaa0;
    defparam time_count_3234_add_4_9.INIT1 = 16'h0000;
    defparam time_count_3234_add_4_9.INJECT1_0 = "NO";
    defparam time_count_3234_add_4_9.INJECT1_1 = "NO";
    LUT4 i12099_2_lut (.A(qspi_data_in[0]), .B(rst_reg_n), .Z(qspi_data_out_3__N_5[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(127[22:56])
    defparam i12099_2_lut.init = 16'h8888;
    CCU2C time_count_3234_add_4_7 (.A0(time_count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19945), .COUT(n19946), .S0(n40), .S1(n39));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3234_add_4_7.INIT0 = 16'haaa0;
    defparam time_count_3234_add_4_7.INIT1 = 16'haaa0;
    defparam time_count_3234_add_4_7.INJECT1_0 = "NO";
    defparam time_count_3234_add_4_7.INJECT1_1 = "NO";
    LUT4 i22459_4_lut (.A(is_writing), .B(is_writing_N_2331), .C(n27082), 
         .D(n6930), .Z(n24802)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i22459_4_lut.init = 16'hcaaa;
    LUT4 i12100_2_lut (.A(debug_rd_r[0]), .B(debug_register_data), .Z(uo_out_c_2)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(154[24:73])
    defparam i12100_2_lut.init = 16'h8888;
    LUT4 i3367_4_lut (.A(n23252), .B(n27083), .C(n5508), .D(n27080), 
         .Z(clk_c_enable_358)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C))) */ ;
    defparam i3367_4_lut.init = 16'hfcdc;
    LUT4 i23470_4_lut (.A(n27279), .B(rst_reg_n_adj_2691), .C(n27306), 
         .D(interrupt_core), .Z(clk_c_enable_367)) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))))) */ ;
    defparam i23470_4_lut.init = 16'h3f3b;
    LUT4 i3361_4_lut (.A(n23276), .B(n27083), .C(n5505), .D(n27080), 
         .Z(clk_c_enable_369)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C))) */ ;
    defparam i3361_4_lut.init = 16'hfcdc;
    LUT4 i1_2_lut_rep_612 (.A(n24118), .B(n17432), .Z(n27237)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_2_lut_rep_612.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_495 (.A(n24118), .B(n17432), .C(addr[4]), 
         .Z(n44_adj_2692)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_2_lut_3_lut_adj_495.init = 16'h1010;
    LUT4 i1_3_lut_rep_599_4_lut (.A(n24118), .B(n17432), .C(addr[5]), 
         .D(addr[4]), .Z(n27224)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_3_lut_rep_599_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_4_lut (.A(n24118), .B(n17432), .C(n3), .D(n24140), 
         .Z(data_from_read[2])) /* synthesis lut_function=(A (B)+!A (B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_4_lut_4_lut.init = 16'hddcd;
    LUT4 rst_reg_n_bdd_4_lut (.A(cycle[0]), .B(n27110), .C(n27342), .D(cycle[1]), 
         .Z(n26801)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C)))) */ ;
    defparam rst_reg_n_bdd_4_lut.init = 16'h3a1a;
    LUT4 i1345_4_lut (.A(pc[2]), .B(n2101), .C(debug_instr_valid), .D(pc[1]), 
         .Z(n2035)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i1345_4_lut.init = 16'hc5c0;
    LUT4 gnd_bdd_2_lut_24180 (.A(n26801), .B(rst_reg_n_adj_2691), .Z(n26802)) /* synthesis lut_function=(A (B)) */ ;
    defparam gnd_bdd_2_lut_24180.init = 16'h8888;
    LUT4 i3370_4_lut (.A(n22992), .B(n27083), .C(n27081), .D(n27299), 
         .Z(clk_c_enable_346)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;
    defparam i3370_4_lut.init = 16'heefc;
    LUT4 i22460_4_lut (.A(writing), .B(n22999), .C(n24428), .Z(n24803)) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam i22460_4_lut.init = 16'hbaba;
    sim_qspi_pmod i_qspi (.qspi_data_in({qspi_data_in}), .qspi_clk_N_56(qspi_clk_N_56), 
            .spi_clk_pos_derived_59(spi_clk_pos_derived_59), .GND_net(GND_net), 
            .VCC_net(VCC_net), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .\addr[14] (addr_adj_2695[14]), .\addr_24__N_228[14] (addr_24__N_228[14]), 
            .\addr[13] (addr_adj_2695[13]), .\addr[12] (addr_adj_2695[12]), 
            .\addr[11] (addr_adj_2695[11]), .\addr[10] (addr_adj_2695[10]), 
            .\addr[9] (addr_adj_2695[9]), .\addr[8] (addr_adj_2695[8]), 
            .writing(writing), .\addr[7] (addr_adj_2695[7]), .\addr[6] (addr_adj_2695[6]), 
            .\addr[5] (addr_adj_2695[5]), .\addr[4] (addr_adj_2695[4]), 
            .\addr[3] (addr_adj_2695[3]), .\addr[2] (addr_adj_2695[2]), 
            .\addr[1] (addr_adj_2695[1]), .n24803(n24803), .\addr[0] (addr_adj_2695[0]), 
            .qspi_ram_a_select(qspi_ram_a_select), .\addr_24__N_228[0] (addr_24__N_228[0]), 
            .n22999(n22999), .\writing_N_164[3] (writing_N_164[3]), .qspi_ram_b_select(qspi_ram_b_select), 
            .\addr_24__N_228[12] (addr_24__N_228[12]), .\addr_24__N_228[2] (addr_24__N_228[2]), 
            .\addr_24__N_228[1] (addr_24__N_228[1]), .\addr_24__N_228[3] (addr_24__N_228[3]), 
            .\addr_24__N_228[4] (addr_24__N_228[4]), .\addr_24__N_228[5] (addr_24__N_228[5]), 
            .\addr_24__N_228[6] (addr_24__N_228[6]), .\addr_24__N_228[7] (addr_24__N_228[7]), 
            .\addr_24__N_228[8] (addr_24__N_228[8]), .\addr_24__N_228[9] (addr_24__N_228[9]), 
            .\addr_24__N_228[10] (addr_24__N_228[10]), .\addr_24__N_228[13] (addr_24__N_228[13]), 
            .\addr_24__N_228[11] (addr_24__N_228[11]), .n27335(n27335), 
            .n24428(n24428)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(42[19] 50[6])
    LUT4 i1_2_lut_adj_496 (.A(addr[4]), .B(addr[3]), .Z(n24260)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_2_lut_adj_496.init = 16'h8888;
    LUT4 i1_4_lut_adj_497 (.A(addr[10]), .B(n24114), .C(n24110), .D(addr[8]), 
         .Z(n24118)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_4_lut_adj_497.init = 16'hfffe;
    LUT4 i1_3_lut (.A(addr[1]), .B(addr[7]), .C(addr[0]), .Z(n24114)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_498 (.A(addr[6]), .B(addr[9]), .Z(n24110)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_2_lut_adj_498.init = 16'heeee;
    LUT4 i1_2_lut_adj_499 (.A(addr[3]), .B(addr[5]), .Z(n24376)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_2_lut_adj_499.init = 16'h4444;
    LUT4 i4850_3_lut (.A(ui_in_c_1), .B(data_to_write[0]), .C(rst_reg_n), 
         .Z(n7164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(234[12] 239[8])
    defparam i4850_3_lut.init = 16'hcaca;
    LUT4 i12136_2_lut (.A(qspi_data_in[2]), .B(rst_reg_n), .Z(qspi_data_out_3__N_5[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(127[22:56])
    defparam i12136_2_lut.init = 16'h8888;
    LUT4 i22657_2_lut_rep_502_4_lut (.A(pc[2]), .B(n27297), .C(debug_instr_valid), 
         .D(n4057), .Z(n27127)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i22657_2_lut_rep_502_4_lut.init = 16'h0035;
    LUT4 i12102_2_lut (.A(debug_rd_r[2]), .B(debug_register_data), .Z(uo_out_c_4)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(156[24:73])
    defparam i12102_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_500 (.A(n24314), .B(n24561), .C(time_count[2]), 
         .D(n24312), .Z(n8869)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_500.init = 16'hffbf;
    LUT4 i1_3_lut_adj_501 (.A(time_count[4]), .B(time_count[1]), .C(time_count[7]), 
         .Z(n24314)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_501.init = 16'hfefe;
    LUT4 i22461_4_lut (.A(mem_op_increment_reg), .B(mem_op_increment_reg_de), 
         .C(n23908), .D(n27106), .Z(n24804)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i22461_4_lut.init = 16'hcaaa;
    LUT4 i22283_2_lut (.A(time_count[3]), .B(time_count[0]), .Z(n24561)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22283_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_502 (.A(time_count[5]), .B(time_count[6]), .Z(n24312)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_502.init = 16'heeee;
    LUT4 i12103_2_lut (.A(debug_rd_r[3]), .B(debug_register_data), .Z(uo_out_c_5)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(157[24:73])
    defparam i12103_2_lut.init = 16'h8888;
    LUT4 i12105_2_lut (.A(debug_uart_txd), .B(gpio_out_sel[6]), .Z(uo_out_c_6)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(158[24:70])
    defparam i12105_2_lut.init = 16'h2222;
    LUT4 i23487_2_lut (.A(n8869), .B(rst_reg_n), .Z(n808)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i23487_2_lut.init = 16'h7777;
    LUT4 i12101_2_lut (.A(debug_rd_r[1]), .B(debug_register_data), .Z(uo_out_c_3)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(155[24:73])
    defparam i12101_2_lut.init = 16'h8888;
    PFUMX i24345 (.BLUT(n27392), .ALUT(n27393), .C0(n1167), .Z(clk_c_enable_350));
    
endmodule
//
// Verilog Description of module \uart_tx(BIT_RATE=1000000,CLK_HZ=14000000) 
//

module \uart_tx(BIT_RATE=1000000,CLK_HZ=14000000)  (debug_uart_txd, clk_c, 
            clk_c_enable_341, clk_c_enable_426, n27294, debug_uart_tx_start, 
            \data_to_write[4] , \data_to_write[5] , \data_to_write[6] , 
            rst_reg_n, n27210, next_bit, uart_txd_N_2596, \data_to_write[2] , 
            \data_to_write[1] , \data_to_write[0] , \data_to_write[7] , 
            \data_to_write[3] ) /* synthesis syn_module_defined=1 */ ;
    output debug_uart_txd;
    input clk_c;
    input clk_c_enable_341;
    input clk_c_enable_426;
    output n27294;
    input debug_uart_tx_start;
    input \data_to_write[4] ;
    input \data_to_write[5] ;
    input \data_to_write[6] ;
    input rst_reg_n;
    output n27210;
    output next_bit;
    output uart_txd_N_2596;
    input \data_to_write[2] ;
    input \data_to_write[1] ;
    input \data_to_write[0] ;
    input \data_to_write[7] ;
    input \data_to_write[3] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire uart_txd_N_2594;
    wire [7:0]data_to_send;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(51[24:36])
    
    wire n23012;
    wire [7:0]data_to_send_7__N_2574;
    wire [3:0]fsm_state;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(59[11:20])
    
    wire n27406;
    wire [4:0]cycle_counter;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(55[25:38])
    wire [4:0]n50;
    
    wire n27261;
    wire [4:0]n18;
    
    wire n27030, n27036, n27363, n27194, n7228, clk_c_enable_362, 
        clk_c_enable_342, n27379;
    wire [3:0]n122;
    
    wire n24446;
    
    FD1S3JX txd_reg_46 (.D(uart_txd_N_2594), .CK(clk_c), .PD(clk_c_enable_341), 
            .Q(debug_uart_txd)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(135[8] 145[4])
    defparam txd_reg_46.GSR = "DISABLED";
    FD1P3AX data_to_send__i7 (.D(n23012), .SP(clk_c_enable_426), .CK(clk_c), 
            .Q(data_to_send[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i7.GSR = "DISABLED";
    LUT4 mux_13_i5_3_lut_4_lut (.A(n27294), .B(debug_uart_tx_start), .C(\data_to_write[4] ), 
         .D(data_to_send[5]), .Z(data_to_send_7__N_2574[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i6_3_lut_4_lut (.A(n27294), .B(debug_uart_tx_start), .C(\data_to_write[5] ), 
         .D(data_to_send[6]), .Z(data_to_send_7__N_2574[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 fsm_state_0__bdd_4_lut (.A(fsm_state[0]), .B(fsm_state[2]), .C(fsm_state[1]), 
         .D(fsm_state[3]), .Z(n27406)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;
    defparam fsm_state_0__bdd_4_lut.init = 16'h4555;
    LUT4 i3627_2_lut (.A(cycle_counter[1]), .B(cycle_counter[0]), .Z(n50[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3627_2_lut.init = 16'h6666;
    LUT4 mux_13_i7_3_lut_4_lut (.A(n27294), .B(debug_uart_tx_start), .C(\data_to_write[6] ), 
         .D(data_to_send[7]), .Z(data_to_send_7__N_2574[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i7_3_lut_4_lut.init = 16'hfb40;
    FD1S3IX cycle_counter__i0 (.D(n18[0]), .CK(clk_c), .CD(n27261), .Q(cycle_counter[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i0.GSR = "DISABLED";
    LUT4 fsm_state_3__bdd_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(fsm_state[0]), .Z(n27030)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B (C (D))))) */ ;
    defparam fsm_state_3__bdd_4_lut.init = 16'h6aa2;
    LUT4 fsm_state_2__bdd_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(fsm_state[0]), 
         .Z(n27036)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam fsm_state_2__bdd_3_lut.init = 16'h6a6a;
    LUT4 i23566_3_lut_rep_569_4_lut (.A(fsm_state[0]), .B(n27363), .C(debug_uart_tx_start), 
         .D(rst_reg_n), .Z(n27194)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(79[9:30])
    defparam i23566_3_lut_rep_569_4_lut.init = 16'h01ff;
    LUT4 i232_2_lut_rep_585_3_lut (.A(fsm_state[0]), .B(n27363), .C(debug_uart_tx_start), 
         .Z(n27210)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(79[9:30])
    defparam i232_2_lut_rep_585_3_lut.init = 16'h1010;
    LUT4 i4913_2_lut_4_lut_2_lut_3_lut (.A(fsm_state[0]), .B(n27363), .C(rst_reg_n), 
         .Z(n7228)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(79[9:30])
    defparam i4913_2_lut_4_lut_2_lut_3_lut.init = 16'h1f1f;
    LUT4 i3274_2_lut_rep_615_3_lut_4_lut (.A(fsm_state[0]), .B(n27363), 
         .C(rst_reg_n), .D(next_bit), .Z(clk_c_enable_362)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(79[9:30])
    defparam i3274_2_lut_rep_615_3_lut_4_lut.init = 16'hffef;
    FD1P3IX fsm_state__i0 (.D(n27406), .SP(clk_c_enable_342), .CD(n27194), 
            .CK(clk_c), .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam fsm_state__i0.GSR = "DISABLED";
    FD1P3IX data_to_send__i1 (.D(data_to_send_7__N_2574[1]), .SP(clk_c_enable_426), 
            .CD(clk_c_enable_341), .CK(clk_c), .Q(data_to_send[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i1.GSR = "DISABLED";
    FD1P3IX data_to_send__i0 (.D(data_to_send_7__N_2574[0]), .SP(clk_c_enable_426), 
            .CD(clk_c_enable_341), .CK(clk_c), .Q(data_to_send[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i0.GSR = "DISABLED";
    LUT4 i12135_4_lut (.A(data_to_send[0]), .B(fsm_state[0]), .C(uart_txd_N_2596), 
         .D(n27363), .Z(uart_txd_N_2594)) /* synthesis lut_function=(A ((D)+!B)+!A !(B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(140[14] 144[8])
    defparam i12135_4_lut.init = 16'haf23;
    LUT4 i3648_3_lut_4_lut (.A(cycle_counter[2]), .B(n27379), .C(cycle_counter[3]), 
         .D(cycle_counter[4]), .Z(n50[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3648_3_lut_4_lut.init = 16'h7f80;
    FD1P3IX data_to_send__i2 (.D(data_to_send_7__N_2574[2]), .SP(clk_c_enable_426), 
            .CD(clk_c_enable_341), .CK(clk_c), .Q(data_to_send[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i2.GSR = "DISABLED";
    FD1P3IX data_to_send__i3 (.D(data_to_send_7__N_2574[3]), .SP(clk_c_enable_426), 
            .CD(clk_c_enable_341), .CK(clk_c), .Q(data_to_send[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i3.GSR = "DISABLED";
    FD1P3IX data_to_send__i4 (.D(data_to_send_7__N_2574[4]), .SP(clk_c_enable_426), 
            .CD(clk_c_enable_341), .CK(clk_c), .Q(data_to_send[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i4.GSR = "DISABLED";
    FD1P3IX fsm_state__i1 (.D(n122[1]), .SP(next_bit), .CD(n7228), .CK(clk_c), 
            .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam fsm_state__i1.GSR = "DISABLED";
    FD1P3IX fsm_state__i2 (.D(n27036), .SP(next_bit), .CD(n7228), .CK(clk_c), 
            .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1P3IX fsm_state__i3 (.D(n27030), .SP(next_bit), .CD(n7228), .CK(clk_c), 
            .Q(fsm_state[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam fsm_state__i3.GSR = "DISABLED";
    FD1P3IX cycle_counter__i1 (.D(n50[1]), .SP(clk_c_enable_362), .CD(n27261), 
            .CK(clk_c), .Q(cycle_counter[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i1.GSR = "DISABLED";
    FD1P3IX cycle_counter__i2 (.D(n50[2]), .SP(clk_c_enable_362), .CD(n27261), 
            .CK(clk_c), .Q(cycle_counter[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i2.GSR = "DISABLED";
    FD1P3IX cycle_counter__i3 (.D(n50[3]), .SP(clk_c_enable_362), .CD(n27261), 
            .CK(clk_c), .Q(cycle_counter[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i3.GSR = "DISABLED";
    FD1P3IX cycle_counter__i4 (.D(n50[4]), .SP(clk_c_enable_362), .CD(n27261), 
            .CK(clk_c), .Q(cycle_counter[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i4.GSR = "DISABLED";
    LUT4 i12175_3_lut_3_lut_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(fsm_state[0]), .Z(n122[1])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(D)))) */ ;
    defparam i12175_3_lut_3_lut_4_lut.init = 16'h33c4;
    LUT4 i23444_4_lut (.A(cycle_counter[0]), .B(cycle_counter[2]), .C(cycle_counter[3]), 
         .D(n24446), .Z(next_bit)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(74[21:71])
    defparam i23444_4_lut.init = 16'h0080;
    LUT4 i1_2_lut (.A(cycle_counter[1]), .B(cycle_counter[4]), .Z(n24446)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3IX data_to_send__i5 (.D(data_to_send_7__N_2574[5]), .SP(clk_c_enable_426), 
            .CD(clk_c_enable_341), .CK(clk_c), .Q(data_to_send[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i5.GSR = "DISABLED";
    FD1P3IX data_to_send__i6 (.D(data_to_send_7__N_2574[6]), .SP(clk_c_enable_426), 
            .CD(clk_c_enable_341), .CK(clk_c), .Q(data_to_send[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i6.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_738 (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[3]), 
         .Z(n27363)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(84[17:37])
    defparam i1_3_lut_rep_738.init = 16'hfefe;
    LUT4 i1_2_lut_rep_669_4_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[3]), 
         .D(fsm_state[0]), .Z(n27294)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(84[17:37])
    defparam i1_2_lut_rep_669_4_lut.init = 16'hfffe;
    LUT4 uart_txd_I_227_4_lut_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(fsm_state[3]), .Z(uart_txd_N_2596)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(84[17:37])
    defparam uart_txd_I_227_4_lut_3_lut.init = 16'h1e1e;
    LUT4 i3629_2_lut_rep_754 (.A(cycle_counter[1]), .B(cycle_counter[0]), 
         .Z(n27379)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3629_2_lut_rep_754.init = 16'h8888;
    LUT4 i3634_2_lut_3_lut (.A(cycle_counter[1]), .B(cycle_counter[0]), 
         .C(cycle_counter[2]), .Z(n50[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3634_2_lut_3_lut.init = 16'h7878;
    LUT4 i3641_2_lut_3_lut_4_lut (.A(cycle_counter[1]), .B(cycle_counter[0]), 
         .C(cycle_counter[3]), .D(cycle_counter[2]), .Z(n50[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3641_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_3_lut_4_lut (.A(n27294), .B(debug_uart_tx_start), .C(next_bit), 
         .D(n27194), .Z(clk_c_enable_342)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam i1_3_lut_4_lut.init = 16'hfff4;
    LUT4 mux_13_i3_3_lut_4_lut (.A(n27294), .B(debug_uart_tx_start), .C(\data_to_write[2] ), 
         .D(data_to_send[3]), .Z(data_to_send_7__N_2574[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i2_3_lut_4_lut (.A(n27294), .B(debug_uart_tx_start), .C(\data_to_write[1] ), 
         .D(data_to_send[2]), .Z(data_to_send_7__N_2574[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i1_3_lut_4_lut (.A(n27294), .B(debug_uart_tx_start), .C(\data_to_write[0] ), 
         .D(data_to_send[1]), .Z(data_to_send_7__N_2574[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut_adj_489 (.A(n27294), .B(debug_uart_tx_start), .C(\data_to_write[7] ), 
         .D(rst_reg_n), .Z(n23012)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam i1_3_lut_4_lut_adj_489.init = 16'h4000;
    LUT4 mux_13_i4_3_lut_4_lut (.A(n27294), .B(debug_uart_tx_start), .C(\data_to_write[3] ), 
         .D(data_to_send[4]), .Z(data_to_send_7__N_2574[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 i23568_2_lut_rep_636 (.A(next_bit), .B(rst_reg_n), .Z(n27261)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i23568_2_lut_rep_636.init = 16'hbbbb;
    LUT4 i4478_2_lut_3_lut_4_lut (.A(next_bit), .B(rst_reg_n), .C(cycle_counter[0]), 
         .D(n27294), .Z(n18[0])) /* synthesis lut_function=(!(A (C)+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam i4478_2_lut_3_lut_4_lut.init = 16'h0f4b;
    
endmodule
//
// Verilog Description of module \peripherals_min(CLOCK_MHZ=14) 
//

module \peripherals_min(CLOCK_MHZ=14)  (peri_data_ready, clk_c, clk_c_enable_341, 
            read_en) /* synthesis syn_module_defined=1 */ ;
    output peri_data_ready;
    input clk_c;
    input clk_c_enable_341;
    input read_en;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    FD1S3DX data_ready_51 (.D(read_en), .CK(clk_c), .CD(clk_c_enable_341), 
            .Q(peri_data_ready)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(139[13:35])
    defparam data_ready_51.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module tinyQV
//

module tinyQV (rst_reg_n_adj_15, clk_c, rst_reg_n, \data_from_read[2] , 
            n27358, \addr[2] , n22303, read_en, n17432, \addr[5] , 
            n24260, n24118, n27269, counter_hi, peri_data_ready, clk_c_enable_341, 
            \instr_addr_23__N_318[0] , \instr_addr_23__N_318[18] , \instr_addr_23__N_318[14] , 
            \instr_addr_23__N_318[15] , \instr_addr_23__N_318[16] , \instr_addr_23__N_318[17] , 
            \instr_addr_23__N_318[6] , \addr[7] , \instr_addr_23__N_318[5] , 
            \addr[6] , \instr_addr_23__N_318[7] , \addr[8] , \instr_addr_23__N_318[3] , 
            \addr[4] , \instr_addr_23__N_318[10] , data_stall, \instr_addr_23__N_318[9] , 
            \addr[10] , \instr_addr_23__N_318[11] , \instr_addr_23__N_318[8] , 
            \addr[9] , \instr_addr[1] , \addr[1] , \instr_addr_23__N_318[12] , 
            \instr_addr_23__N_318[22] , \instr_addr_23__N_318[13] , \instr_addr_23__N_318[4] , 
            \instr_addr_23__N_318[19] , \instr_addr_23__N_318[20] , \instr_addr_23__N_318[21] , 
            n27081, is_writing_N_2331, n27299, \data_to_write[7] , \data_to_write[6] , 
            continue_txn_N_2131, data_stall_N_2158, \data_to_write[5] , 
            \pc[1] , \pc[2] , n24806, \data_to_write[4] , qv_data_write_n, 
            \data_to_write[0] , \data_to_write[3] , \data_to_write[2] , 
            \data_to_write[1] , n27082, \addr[0] , is_writing, \instr_addr_23__N_318[2] , 
            \addr[3] , n6930, \writing_N_164[3] , n27083, qspi_ram_b_select, 
            \qspi_data_out_3__N_5[0] , qspi_ram_a_select, n24802, qspi_data_in, 
            \fsm_state[0] , n23276, clk_c_enable_358, clk_c_enable_369, 
            n23252, clk_N_45, \qspi_data_out_3__N_5[2] , n4319, n4307, 
            \qspi_data_oe[3] , clk_c_enable_346, n27080, \qspi_data_out_3__N_5[3] , 
            \addr[20] , \addr[22] , spi_clk_pos_derived_59, qspi_clk_N_56, 
            next_bit, n27210, uart_txd_N_2596, clk_c_enable_426, n24376, 
            n44, clk_c_enable_273, n805, clk_c_enable_420, n27365, 
            n22097, n4309, n26711, n5508, n5505, n22992, \instr_len[2] , 
            VCC_net, interrupt_core, n2055, debug_instr_valid, was_early_branch, 
            n2035, \pc[10] , n27106, data_ready_sync, n2096, n2101, 
            \imm[23] , n4057, n26793, \imm[22] , \imm[1] , \imm[10] , 
            \imm[21] , \imm[20] , \imm[6] , \imm[19] , \imm[18] , 
            \imm[17] , \imm[16] , \imm[15] , \imm[14] , \imm[13] , 
            \imm[12] , \imm[11] , \imm[9] , \imm[8] , \imm[7] , \imm[5] , 
            \imm[4] , \imm[3] , \imm[2] , is_timer_addr, n27354, n27342, 
            \addr_out[1] , \instr_write_offset[3] , n27297, mem_op_increment_reg, 
            n24804, \pc[23] , \next_pc_for_core[6] , \next_pc_for_core[4] , 
            \next_pc_for_core[9] , \next_pc_for_core[13] , \pc[8] , \pc[12] , 
            \next_pc_for_core[3] , \next_pc_for_core[5] , \pc[4] , \next_pc_for_core[7] , 
            \next_pc_for_core[8] , \next_pc_for_core[10] , \next_pc_for_core[12] , 
            \next_pc_for_core[11] , \next_pc_for_core[14] , \next_pc_for_core[15] , 
            \next_pc_for_core[16] , \next_pc_for_core[17] , \next_pc_for_core[18] , 
            \next_pc_for_core[19] , \next_pc_for_core[20] , \next_pc_for_core[21] , 
            \next_pc_for_core[22] , \next_pc_for_core[23] , \pc[22] , 
            \pc[21] , \pc[20] , \pc[19] , \pc[18] , \pc[17] , \pc[16] , 
            \pc[15] , \pc[14] , \pc[13] , \pc[11] , \pc[9] , \pc[7] , 
            \pc[6] , \pc[5] , \pc[3] , n27127, n27110, cycle, n27350, 
            \early_branch_addr[3] , \early_branch_addr[6] , \early_branch_addr[2] , 
            \early_branch_addr[5] , \early_branch_addr[4] , \early_branch_addr[7] , 
            \early_branch_addr[8] , \early_branch_addr[9] , \early_branch_addr[10] , 
            \early_branch_addr[11] , \early_branch_addr[12] , \early_branch_addr[13] , 
            \early_branch_addr[14] , \early_branch_addr[15] , \early_branch_addr[16] , 
            \early_branch_addr[17] , \early_branch_addr[18] , \early_branch_addr[19] , 
            \early_branch_addr[20] , \early_branch_addr[21] , \early_branch_addr[22] , 
            \early_branch_addr[23] , n27294, n27306, \data_from_read[6] , 
            n24126, n27241, n8869, n27279, n23908, n27220, mem_op_increment_reg_de, 
            n27218, \next_fsm_state_3__N_2499[3] , clk_c_enable_350, clk_c_enable_367, 
            \mul_out[2] , \mul_out[3] , \mul_out[1] , \ui_in_sync[1] , 
            n1167, debug_rd, accum, d_3__N_1868, n4577, n26802, 
            n27223, \next_accum[5] , \next_accum[6] , \next_accum[7] , 
            GND_net, \next_accum[8] , \next_accum[9] , \next_accum[10] , 
            \next_accum[11] , \next_accum[12] , \next_accum[13] , \next_accum[14] , 
            \next_accum[15] , \next_accum[16] , \next_accum[17] , \next_accum[18] , 
            \next_accum[19] , \next_accum[4] ) /* synthesis syn_module_defined=1 */ ;
    output rst_reg_n_adj_15;
    input clk_c;
    input rst_reg_n;
    input \data_from_read[2] ;
    input n27358;
    output \addr[2] ;
    output n22303;
    output read_en;
    output n17432;
    output \addr[5] ;
    input n24260;
    input n24118;
    output n27269;
    output [4:2]counter_hi;
    input peri_data_ready;
    output clk_c_enable_341;
    output \instr_addr_23__N_318[0] ;
    input \instr_addr_23__N_318[18] ;
    input \instr_addr_23__N_318[14] ;
    input \instr_addr_23__N_318[15] ;
    input \instr_addr_23__N_318[16] ;
    input \instr_addr_23__N_318[17] ;
    input \instr_addr_23__N_318[6] ;
    output \addr[7] ;
    input \instr_addr_23__N_318[5] ;
    output \addr[6] ;
    input \instr_addr_23__N_318[7] ;
    output \addr[8] ;
    input \instr_addr_23__N_318[3] ;
    output \addr[4] ;
    input \instr_addr_23__N_318[10] ;
    output data_stall;
    input \instr_addr_23__N_318[9] ;
    output \addr[10] ;
    input \instr_addr_23__N_318[11] ;
    input \instr_addr_23__N_318[8] ;
    output \addr[9] ;
    input \instr_addr[1] ;
    output \addr[1] ;
    input \instr_addr_23__N_318[12] ;
    input \instr_addr_23__N_318[22] ;
    input \instr_addr_23__N_318[13] ;
    input \instr_addr_23__N_318[4] ;
    input \instr_addr_23__N_318[19] ;
    input \instr_addr_23__N_318[20] ;
    input \instr_addr_23__N_318[21] ;
    output n27081;
    output is_writing_N_2331;
    output n27299;
    output \data_to_write[7] ;
    output \data_to_write[6] ;
    output continue_txn_N_2131;
    output data_stall_N_2158;
    output \data_to_write[5] ;
    output \pc[1] ;
    output \pc[2] ;
    input n24806;
    output \data_to_write[4] ;
    output [1:0]qv_data_write_n;
    output \data_to_write[0] ;
    output \data_to_write[3] ;
    output \data_to_write[2] ;
    output \data_to_write[1] ;
    output n27082;
    output \addr[0] ;
    output is_writing;
    input \instr_addr_23__N_318[2] ;
    output \addr[3] ;
    output n6930;
    output \writing_N_164[3] ;
    output n27083;
    output qspi_ram_b_select;
    input \qspi_data_out_3__N_5[0] ;
    output qspi_ram_a_select;
    input n24802;
    input [3:0]qspi_data_in;
    output \fsm_state[0] ;
    output n23276;
    input clk_c_enable_358;
    input clk_c_enable_369;
    output n23252;
    input clk_N_45;
    input \qspi_data_out_3__N_5[2] ;
    output n4319;
    output n4307;
    output \qspi_data_oe[3] ;
    input clk_c_enable_346;
    output n27080;
    input \qspi_data_out_3__N_5[3] ;
    output \addr[20] ;
    output \addr[22] ;
    output spi_clk_pos_derived_59;
    output qspi_clk_N_56;
    input next_bit;
    input n27210;
    input uart_txd_N_2596;
    output clk_c_enable_426;
    input n24376;
    input n44;
    output clk_c_enable_273;
    input n805;
    output clk_c_enable_420;
    output n27365;
    output n22097;
    output n4309;
    output n26711;
    output n5508;
    output n5505;
    output n22992;
    output \instr_len[2] ;
    input VCC_net;
    output interrupt_core;
    input n2055;
    output debug_instr_valid;
    output was_early_branch;
    input n2035;
    output \pc[10] ;
    output n27106;
    output data_ready_sync;
    output n2096;
    output n2101;
    output \imm[23] ;
    output n4057;
    input n26793;
    output \imm[22] ;
    output \imm[1] ;
    output \imm[10] ;
    output \imm[21] ;
    output \imm[20] ;
    output \imm[6] ;
    output \imm[19] ;
    output \imm[18] ;
    output \imm[17] ;
    output \imm[16] ;
    output \imm[15] ;
    output \imm[14] ;
    output \imm[13] ;
    output \imm[12] ;
    output \imm[11] ;
    output \imm[9] ;
    output \imm[8] ;
    output \imm[7] ;
    output \imm[5] ;
    output \imm[4] ;
    output \imm[3] ;
    output \imm[2] ;
    output is_timer_addr;
    output n27354;
    output n27342;
    output \addr_out[1] ;
    output \instr_write_offset[3] ;
    output n27297;
    output mem_op_increment_reg;
    input n24804;
    output \pc[23] ;
    input \next_pc_for_core[6] ;
    input \next_pc_for_core[4] ;
    input \next_pc_for_core[9] ;
    input \next_pc_for_core[13] ;
    output \pc[8] ;
    output \pc[12] ;
    input \next_pc_for_core[3] ;
    input \next_pc_for_core[5] ;
    output \pc[4] ;
    input \next_pc_for_core[7] ;
    input \next_pc_for_core[8] ;
    input \next_pc_for_core[10] ;
    input \next_pc_for_core[12] ;
    input \next_pc_for_core[11] ;
    input \next_pc_for_core[14] ;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[16] ;
    input \next_pc_for_core[17] ;
    input \next_pc_for_core[18] ;
    input \next_pc_for_core[19] ;
    input \next_pc_for_core[20] ;
    input \next_pc_for_core[21] ;
    input \next_pc_for_core[22] ;
    input \next_pc_for_core[23] ;
    output \pc[22] ;
    output \pc[21] ;
    output \pc[20] ;
    output \pc[19] ;
    output \pc[18] ;
    output \pc[17] ;
    output \pc[16] ;
    output \pc[15] ;
    output \pc[14] ;
    output \pc[13] ;
    output \pc[11] ;
    output \pc[9] ;
    output \pc[7] ;
    output \pc[6] ;
    output \pc[5] ;
    output \pc[3] ;
    input n27127;
    output n27110;
    output [1:0]cycle;
    output n27350;
    input \early_branch_addr[3] ;
    input \early_branch_addr[6] ;
    input \early_branch_addr[2] ;
    input \early_branch_addr[5] ;
    input \early_branch_addr[4] ;
    input \early_branch_addr[7] ;
    input \early_branch_addr[8] ;
    input \early_branch_addr[9] ;
    input \early_branch_addr[10] ;
    input \early_branch_addr[11] ;
    input \early_branch_addr[12] ;
    input \early_branch_addr[13] ;
    input \early_branch_addr[14] ;
    input \early_branch_addr[15] ;
    input \early_branch_addr[16] ;
    input \early_branch_addr[17] ;
    input \early_branch_addr[18] ;
    input \early_branch_addr[19] ;
    input \early_branch_addr[20] ;
    input \early_branch_addr[21] ;
    input \early_branch_addr[22] ;
    input \early_branch_addr[23] ;
    input n27294;
    output n27306;
    input \data_from_read[6] ;
    input n24126;
    input n27241;
    input n8869;
    output n27279;
    output n23908;
    input n27220;
    output mem_op_increment_reg_de;
    output n27218;
    input \next_fsm_state_3__N_2499[3] ;
    input clk_c_enable_350;
    input clk_c_enable_367;
    input \mul_out[2] ;
    input \mul_out[3] ;
    input \mul_out[1] ;
    input \ui_in_sync[1] ;
    output n1167;
    output [3:0]debug_rd;
    output [15:0]accum;
    output [19:0]d_3__N_1868;
    input n4577;
    input n26802;
    input n27223;
    input \next_accum[5] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input GND_net;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[4] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    wire [27:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    
    wire n27357, n24751, n24753, n24745, n24747, n27356, n22344;
    wire [31:0]mem_data_from_read;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(74[15:33])
    
    wire n24778, n24757, n24759, n24744, n9091, n25239;
    wire [59:0]debug_branch_N_840;
    wire [1:0]qv_data_read_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(65[15:29])
    
    wire n26088, n26089, n27271, n27298, n27268, n28575, mem_data_ready, 
        n10, n24100, n24102, n24092, n24088, n24098, n24080, debug_data_continue;
    wire [1:0]data_txn_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(49[15:27])
    wire [15:0]instr_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(61[15:25])
    
    wire start_instr, instr_fetch_running, n27334, n23526, n27333, 
        n23532, n27255, n27327, n23536;
    wire [31:0]qspi_data_buf;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(58[16:29])
    wire [23:1]instr_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(56[15:25])
    wire [31:0]data_to_write;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(56[17:30])
    
    wire instr_fetch_stopped;
    wire [3:1]next_instr_write_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[16:39])
    
    wire instr_fetch_running_N_945, n27093, n27150, debug_stop_txn_N_2148, 
        n27341, n23432, n27277, n27233, debug_stop_txn_N_2147, n22591, 
        n24743, n24742, n26794, n26730, n26714, n27227;
    
    FD1S3AX rst_reg_n_16 (.D(rst_reg_n), .CK(clk_c), .Q(rst_reg_n_adj_15)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=111, LSE_RLINE=150 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(92[10:43])
    defparam rst_reg_n_16.GSR = "DISABLED";
    LUT4 i22410_3_lut_4_lut (.A(addr[27]), .B(n27357), .C(\data_from_read[2] ), 
         .D(n24751), .Z(n24753)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i22410_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i22404_3_lut_4_lut (.A(addr[27]), .B(n27357), .C(\data_from_read[2] ), 
         .D(n24745), .Z(n24747)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i22404_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i20124_3_lut_4_lut (.A(addr[27]), .B(n27357), .C(n27358), .D(n27356), 
         .Z(n22344)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i20124_3_lut_4_lut.init = 16'hfeee;
    LUT4 i20084_2_lut_3_lut_4_lut (.A(addr[27]), .B(n27357), .C(\addr[2] ), 
         .D(n27358), .Z(n22303)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i20084_2_lut_3_lut_4_lut.init = 16'hfff1;
    LUT4 i22435_3_lut_4_lut (.A(addr[27]), .B(n27357), .C(\data_from_read[2] ), 
         .D(mem_data_from_read[3]), .Z(n24778)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i22435_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i22416_3_lut_4_lut (.A(addr[27]), .B(n27357), .C(\data_from_read[2] ), 
         .D(n24757), .Z(n24759)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i22416_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6751_3_lut_4_lut (.A(addr[27]), .B(n27357), .C(\data_from_read[2] ), 
         .D(n24744), .Z(n9091)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i6751_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6779_3_lut_4_lut (.A(addr[27]), .B(n27357), .C(\data_from_read[2] ), 
         .D(n25239), .Z(debug_branch_N_840[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i6779_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23527_3_lut_4_lut (.A(addr[27]), .B(n27357), .C(qv_data_read_n[0]), 
         .D(qv_data_read_n[1]), .Z(read_en)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i23527_3_lut_4_lut.init = 16'h0e00;
    LUT4 n26088_bdd_2_lut (.A(n26088), .B(n17432), .Z(n26089)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n26088_bdd_2_lut.init = 16'h2222;
    LUT4 addr_2__bdd_4_lut_24096 (.A(\addr[2] ), .B(\addr[5] ), .C(n24260), 
         .D(n24118), .Z(n26088)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam addr_2__bdd_4_lut_24096.init = 16'hff80;
    LUT4 i1_2_lut_rep_732 (.A(addr[26]), .B(addr[25]), .Z(n27357)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_rep_732.init = 16'heeee;
    LUT4 i12800_2_lut_rep_646_3_lut_4_lut (.A(addr[26]), .B(addr[25]), .C(n27358), 
         .D(addr[27]), .Z(n27271)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i12800_2_lut_rep_646_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_673_3_lut (.A(addr[26]), .B(addr[25]), .C(addr[27]), 
         .Z(n27298)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_rep_673_3_lut.init = 16'hfefe;
    LUT4 i12827_2_lut_rep_644_3_lut_4_lut (.A(addr[26]), .B(addr[25]), .C(n27358), 
         .D(addr[27]), .Z(n27269)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i12827_2_lut_rep_644_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i23680_2_lut_rep_643_3_lut_4_lut (.A(addr[26]), .B(addr[25]), .C(counter_hi[3]), 
         .D(addr[27]), .Z(n27268)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i23680_2_lut_rep_643_3_lut_4_lut.init = 16'hffef;
    FD1S3AX rst_reg_n_16_rep_766 (.D(rst_reg_n), .CK(clk_c), .Q(n28575)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=111, LSE_RLINE=150 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(92[10:43])
    defparam rst_reg_n_16_rep_766.GSR = "DISABLED";
    LUT4 i25_4_lut (.A(mem_data_ready), .B(peri_data_ready), .C(n27298), 
         .D(n26089), .Z(n10)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C)+!B !((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(77[26:62])
    defparam i25_4_lut.init = 16'h3505;
    LUT4 i1_4_lut (.A(n24100), .B(addr[27]), .C(n24102), .D(n27357), 
         .Z(n17432)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i1_4_lut_adj_484 (.A(addr[12]), .B(n24092), .C(n24088), .D(addr[11]), 
         .Z(n24100)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_4_lut_adj_484.init = 16'hfffe;
    LUT4 i1_4_lut_adj_485 (.A(addr[15]), .B(n24098), .C(n24080), .D(addr[21]), 
         .Z(n24102)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_4_lut_adj_485.init = 16'hfffe;
    LUT4 i1_2_lut (.A(addr[24]), .B(addr[18]), .Z(n24092)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_486 (.A(addr[20]), .B(addr[23]), .Z(n24088)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_adj_486.init = 16'heeee;
    LUT4 i1_4_lut_adj_487 (.A(addr[17]), .B(addr[14]), .C(addr[19]), .D(addr[22]), 
         .Z(n24098)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_4_lut_adj_487.init = 16'hfffe;
    LUT4 i1_2_lut_adj_488 (.A(addr[16]), .B(addr[13]), .Z(n24080)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_adj_488.init = 16'heeee;
    tinyqv_mem_ctrl mem (.clk_c(clk_c), .clk_c_enable_341(clk_c_enable_341), 
            .debug_data_continue(debug_data_continue), .data_txn_len({Open_0, 
            data_txn_len[0]}), .instr_data({instr_data}), .start_instr(start_instr), 
            .instr_fetch_running(instr_fetch_running), .n27334(n27334), 
            .n23526(n23526), .n27333(n27333), .n23532(n23532), .\instr_addr_23__N_318[0] (\instr_addr_23__N_318[0] ), 
            .n27255(n27255), .n27327(n27327), .n23536(n23536), .\instr_addr_23__N_318[18] (\instr_addr_23__N_318[18] ), 
            .\addr[19] (addr[19]), .\instr_addr_23__N_318[14] (\instr_addr_23__N_318[14] ), 
            .\addr[15] (addr[15]), .\qspi_data_buf[29] (qspi_data_buf[29]), 
            .\qspi_data_buf[25] (qspi_data_buf[25]), .\mem_data_from_read[23] (mem_data_from_read[23]), 
            .\mem_data_from_read[22] (mem_data_from_read[22]), .\mem_data_from_read[21] (mem_data_from_read[21]), 
            .\mem_data_from_read[20] (mem_data_from_read[20]), .\mem_data_from_read[19] (mem_data_from_read[19]), 
            .\mem_data_from_read[18] (mem_data_from_read[18]), .\mem_data_from_read[17] (mem_data_from_read[17]), 
            .\mem_data_from_read[16] (mem_data_from_read[16]), .\qspi_data_buf[14] (qspi_data_buf[14]), 
            .\qspi_data_buf[12] (qspi_data_buf[12]), .\qspi_data_buf[10] (qspi_data_buf[10]), 
            .\qspi_data_buf[8] (qspi_data_buf[8]), .\instr_addr_23__N_318[15] (\instr_addr_23__N_318[15] ), 
            .\addr[16] (addr[16]), .\instr_addr_23__N_318[16] (\instr_addr_23__N_318[16] ), 
            .\addr[17] (addr[17]), .\instr_addr_23__N_318[17] (\instr_addr_23__N_318[17] ), 
            .\addr[18] (addr[18]), .\instr_addr_23__N_318[6] (\instr_addr_23__N_318[6] ), 
            .\addr[7] (\addr[7] ), .\instr_addr_23__N_318[5] (\instr_addr_23__N_318[5] ), 
            .\addr[6] (\addr[6] ), .\instr_addr[2] (instr_addr[2]), .\addr[2] (\addr[2] ), 
            .\instr_addr_23__N_318[7] (\instr_addr_23__N_318[7] ), .\addr[8] (\addr[8] ), 
            .\instr_addr_23__N_318[3] (\instr_addr_23__N_318[3] ), .\addr[4] (\addr[4] ), 
            .\instr_addr_23__N_318[10] (\instr_addr_23__N_318[10] ), .\addr[11] (addr[11]), 
            .data_stall(data_stall), .data_to_write({data_to_write[31:8], 
            \data_to_write[7] , \data_to_write[6] , \data_to_write[5] , 
            \data_to_write[4] , \data_to_write[3] , \data_to_write[2] , 
            \data_to_write[1] , \data_to_write[0] }), .\instr_addr_23__N_318[9] (\instr_addr_23__N_318[9] ), 
            .\addr[10] (\addr[10] ), .instr_fetch_stopped(instr_fetch_stopped), 
            .\instr_addr_23__N_318[11] (\instr_addr_23__N_318[11] ), .\addr[12] (addr[12]), 
            .\instr_addr_23__N_318[8] (\instr_addr_23__N_318[8] ), .\addr[9] (\addr[9] ), 
            .rst_reg_n(rst_reg_n), .\instr_addr[1] (\instr_addr[1] ), .\addr[1] (\addr[1] ), 
            .\instr_addr_23__N_318[12] (\instr_addr_23__N_318[12] ), .\addr[13] (addr[13]), 
            .\instr_addr_23__N_318[22] (\instr_addr_23__N_318[22] ), .\addr[23] (addr[23]), 
            .\instr_addr_23__N_318[13] (\instr_addr_23__N_318[13] ), .\addr[14] (addr[14]), 
            .\instr_addr_23__N_318[4] (\instr_addr_23__N_318[4] ), .\addr[5] (\addr[5] ), 
            .\next_instr_write_offset[3] (next_instr_write_offset[3]), .\instr_addr_23__N_318[19] (\instr_addr_23__N_318[19] ), 
            .\addr[20] (addr[20]), .instr_fetch_running_N_945(instr_fetch_running_N_945), 
            .n27093(n27093), .\instr_addr_23__N_318[20] (\instr_addr_23__N_318[20] ), 
            .\addr[21] (addr[21]), .\instr_addr_23__N_318[21] (\instr_addr_23__N_318[21] ), 
            .\addr[22] (addr[22]), .mem_data_ready(mem_data_ready), .n27150(n27150), 
            .n27081(n27081), .is_writing_N_2331(is_writing_N_2331), .\mem_data_from_read[31] (mem_data_from_read[31]), 
            .\mem_data_from_read[27] (mem_data_from_read[27]), .\mem_data_from_read[30] (mem_data_from_read[30]), 
            .\mem_data_from_read[26] (mem_data_from_read[26]), .\mem_data_from_read[28] (mem_data_from_read[28]), 
            .\mem_data_from_read[24] (mem_data_from_read[24]), .n27299(n27299), 
            .debug_stop_txn_N_2148(debug_stop_txn_N_2148), .n27341(n27341), 
            .n23432(n23432), .continue_txn_N_2131(continue_txn_N_2131), 
            .data_stall_N_2158(data_stall_N_2158), .n27271(n27271), .n27277(n27277), 
            .n27233(n27233), .\pc[1] (\pc[1] ), .\pc[2] (\pc[2] ), .n24806(n24806), 
            .n27298(n27298), .debug_stop_txn_N_2147(debug_stop_txn_N_2147), 
            .\addr[24] (addr[24]), .qv_data_write_n({qv_data_write_n}), 
            .qv_data_read_n({qv_data_read_n}), .n22591(n22591), .n22344(n22344), 
            .n27356(n27356), .n27357(n27357), .\addr[27] (addr[27]), .\mem_data_from_read[13] (mem_data_from_read[13]), 
            .\mem_data_from_read[9] (mem_data_from_read[9]), .n24743(n24743), 
            .n24742(n24742), .n26794(n26794), .n26730(n26730), .n26714(n26714), 
            .\mem_data_from_read[4] (mem_data_from_read[4]), .\mem_data_from_read[3] (mem_data_from_read[3]), 
            .\mem_data_from_read[5] (mem_data_from_read[5]), .\mem_data_from_read[1] (mem_data_from_read[1]), 
            .\mem_data_from_read[6] (mem_data_from_read[6]), .n27082(n27082), 
            .\addr[0] (\addr[0] ), .n27358(n27358), .n27227(n27227), .is_writing(is_writing), 
            .\instr_addr_23__N_318[2] (\instr_addr_23__N_318[2] ), .\addr[3] (\addr[3] ), 
            .n6930(n6930), .\writing_N_164[3] (\writing_N_164[3] ), .n27083(n27083), 
            .qspi_ram_b_select(qspi_ram_b_select), .\qspi_data_out_3__N_5[0] (\qspi_data_out_3__N_5[0] ), 
            .qspi_ram_a_select(qspi_ram_a_select), .n24802(n24802), .qspi_data_in({qspi_data_in}), 
            .\fsm_state[0] (\fsm_state[0] ), .n23276(n23276), .clk_c_enable_358(clk_c_enable_358), 
            .clk_c_enable_369(clk_c_enable_369), .n23252(n23252), .clk_N_45(clk_N_45), 
            .\qspi_data_out_3__N_5[2] (\qspi_data_out_3__N_5[2] ), .n4319(n4319), 
            .n4307(n4307), .\qspi_data_oe[3] (\qspi_data_oe[3] ), .clk_c_enable_346(clk_c_enable_346), 
            .n27080(n27080), .\qspi_data_out_3__N_5[3] (\qspi_data_out_3__N_5[3] ), 
            .\addr[20]_adj_13 (\addr[20] ), .\addr[22]_adj_14 (\addr[22] ), 
            .spi_clk_pos_derived_59(spi_clk_pos_derived_59), .qspi_clk_N_56(qspi_clk_N_56), 
            .next_bit(next_bit), .n27210(n27210), .uart_txd_N_2596(uart_txd_N_2596), 
            .clk_c_enable_426(clk_c_enable_426), .n24376(n24376), .n22303(n22303), 
            .n44(n44), .clk_c_enable_273(clk_c_enable_273), .n805(n805), 
            .clk_c_enable_420(clk_c_enable_420), .n27365(n27365), .n22097(n22097), 
            .n4309(n4309), .n26711(n26711), .n5508(n5508), .n5505(n5505), 
            .n22992(n22992)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(132[19] 164[6])
    tinyqv_cpu cpu (.clk_c(clk_c), .instr_len({\instr_len[2] , Open_1}), 
            .VCC_net(VCC_net), .interrupt_core(interrupt_core), .data_to_write({data_to_write[31:8], 
            \data_to_write[7] , \data_to_write[6] , \data_to_write[5] , 
            \data_to_write[4] , \data_to_write[3] , \data_to_write[2] , 
            \data_to_write[1] , \data_to_write[0] }), .n2055(n2055), .qv_data_read_n({qv_data_read_n}), 
            .\instr_addr_23__N_318[0] (\instr_addr_23__N_318[0] ), .addr({addr[27:11], 
            \addr[10] , \addr[9] , \addr[8] , \addr[7] , \addr[6] , 
            \addr[5] , \addr[4] , \addr[3] , \addr[2] , \addr[1] , 
            \addr[0] }), .debug_data_continue(debug_data_continue), .counter_hi({counter_hi}), 
            .debug_instr_valid(debug_instr_valid), .was_early_branch(was_early_branch), 
            .n2035(n2035), .\pc[2] (\pc[2] ), .\pc[10] (\pc[10] ), .mem_data_ready(mem_data_ready), 
            .n27106(n27106), .data_ready_sync(data_ready_sync), .\pc[1] (\pc[1] ), 
            .n2096(n2096), .n2101(n2101), .n28575(n28575), .rst_reg_n(rst_reg_n_adj_15), 
            .instr_data({instr_data}), .\data_txn_len[0] (data_txn_len[0]), 
            .\qspi_data_buf[12] (qspi_data_buf[12]), .n27150(n27150), .\qspi_data_buf[8] (qspi_data_buf[8]), 
            .\qspi_data_buf[14] (qspi_data_buf[14]), .\qspi_data_buf[10] (qspi_data_buf[10]), 
            .\imm[23] (\imm[23] ), .n4057(n4057), .n26794(n26794), .n26793(n26793), 
            .n27298(n27298), .\imm[22] (\imm[22] ), .\imm[1] (\imm[1] ), 
            .\imm[10] (\imm[10] ), .instr_fetch_running(instr_fetch_running), 
            .\imm[21] (\imm[21] ), .\imm[20] (\imm[20] ), .\imm[6] (\imm[6] ), 
            .\imm[19] (\imm[19] ), .\imm[18] (\imm[18] ), .\imm[17] (\imm[17] ), 
            .qv_data_write_n({qv_data_write_n}), .\imm[16] (\imm[16] ), 
            .\imm[15] (\imm[15] ), .\imm[14] (\imm[14] ), .\imm[13] (\imm[13] ), 
            .\imm[12] (\imm[12] ), .\imm[11] (\imm[11] ), .\imm[9] (\imm[9] ), 
            .\imm[8] (\imm[8] ), .\imm[7] (\imm[7] ), .\imm[5] (\imm[5] ), 
            .\imm[4] (\imm[4] ), .\imm[3] (\imm[3] ), .\imm[2] (\imm[2] ), 
            .is_timer_addr(is_timer_addr), .n27354(n27354), .n27342(n27342), 
            .\addr_out[1] (\addr_out[1] ), .\instr_write_offset[3] (\instr_write_offset[3] ), 
            .\next_instr_write_offset[3] (next_instr_write_offset[3]), .n27297(n27297), 
            .n26730(n26730), .\mem_data_from_read[4] (mem_data_from_read[4]), 
            .mem_op_increment_reg(mem_op_increment_reg), .n24804(n24804), 
            .n26714(n26714), .\mem_data_from_read[6] (mem_data_from_read[6]), 
            .\mem_data_from_read[27] (mem_data_from_read[27]), .\mem_data_from_read[31] (mem_data_from_read[31]), 
            .\pc[23] (\pc[23] ), .debug_stop_txn_N_2148(debug_stop_txn_N_2148), 
            .debug_stop_txn_N_2147(debug_stop_txn_N_2147), .\next_pc_for_core[6] (\next_pc_for_core[6] ), 
            .n24747(n24747), .n24753(n24753), .\next_pc_for_core[4] (\next_pc_for_core[4] ), 
            .\next_pc_for_core[9] (\next_pc_for_core[9] ), .\next_pc_for_core[13] (\next_pc_for_core[13] ), 
            .n24778(n24778), .n25239(n25239), .\pc[8] (\pc[8] ), .\pc[12] (\pc[12] ), 
            .\next_pc_for_core[3] (\next_pc_for_core[3] ), .\next_pc_for_core[5] (\next_pc_for_core[5] ), 
            .\pc[4] (\pc[4] ), .\next_pc_for_core[7] (\next_pc_for_core[7] ), 
            .\next_pc_for_core[8] (\next_pc_for_core[8] ), .\next_pc_for_core[10] (\next_pc_for_core[10] ), 
            .\next_pc_for_core[12] (\next_pc_for_core[12] ), .\next_pc_for_core[11] (\next_pc_for_core[11] ), 
            .\next_pc_for_core[14] (\next_pc_for_core[14] ), .\next_pc_for_core[15] (\next_pc_for_core[15] ), 
            .\next_pc_for_core[16] (\next_pc_for_core[16] ), .\next_pc_for_core[17] (\next_pc_for_core[17] ), 
            .\next_pc_for_core[18] (\next_pc_for_core[18] ), .\next_pc_for_core[19] (\next_pc_for_core[19] ), 
            .\next_pc_for_core[20] (\next_pc_for_core[20] ), .\next_pc_for_core[21] (\next_pc_for_core[21] ), 
            .\next_pc_for_core[22] (\next_pc_for_core[22] ), .\next_pc_for_core[23] (\next_pc_for_core[23] ), 
            .\pc[22] (\pc[22] ), .\pc[21] (\pc[21] ), .\pc[20] (\pc[20] ), 
            .\pc[19] (\pc[19] ), .\pc[18] (\pc[18] ), .\pc[17] (\pc[17] ), 
            .\pc[16] (\pc[16] ), .\pc[15] (\pc[15] ), .\pc[14] (\pc[14] ), 
            .\pc[13] (\pc[13] ), .\pc[11] (\pc[11] ), .\pc[9] (\pc[9] ), 
            .\pc[7] (\pc[7] ), .\pc[6] (\pc[6] ), .\pc[5] (\pc[5] ), .\pc[3] (\pc[3] ), 
            .\mem_data_from_read[19] (mem_data_from_read[19]), .\mem_data_from_read[23] (mem_data_from_read[23]), 
            .n24757(n24757), .n27327(n27327), .\mem_data_from_read[16] (mem_data_from_read[16]), 
            .\mem_data_from_read[20] (mem_data_from_read[20]), .n24745(n24745), 
            .\mem_data_from_read[18] (mem_data_from_read[18]), .\mem_data_from_read[22] (mem_data_from_read[22]), 
            .n24751(n24751), .n27127(n27127), .n27333(n27333), .n27334(n27334), 
            .n27110(n27110), .n27341(n27341), .cycle({cycle}), .n27227(n27227), 
            .start_instr(start_instr), .n23432(n23432), .n27350(n27350), 
            .\early_branch_addr[3] (\early_branch_addr[3] ), .\early_branch_addr[6] (\early_branch_addr[6] ), 
            .\early_branch_addr[2] (\early_branch_addr[2] ), .\early_branch_addr[5] (\early_branch_addr[5] ), 
            .\early_branch_addr[4] (\early_branch_addr[4] ), .\early_branch_addr[7] (\early_branch_addr[7] ), 
            .\early_branch_addr[8] (\early_branch_addr[8] ), .\early_branch_addr[9] (\early_branch_addr[9] ), 
            .\early_branch_addr[10] (\early_branch_addr[10] ), .\early_branch_addr[11] (\early_branch_addr[11] ), 
            .\early_branch_addr[12] (\early_branch_addr[12] ), .\early_branch_addr[13] (\early_branch_addr[13] ), 
            .\early_branch_addr[14] (\early_branch_addr[14] ), .\early_branch_addr[15] (\early_branch_addr[15] ), 
            .\early_branch_addr[16] (\early_branch_addr[16] ), .\early_branch_addr[17] (\early_branch_addr[17] ), 
            .\early_branch_addr[18] (\early_branch_addr[18] ), .\early_branch_addr[19] (\early_branch_addr[19] ), 
            .\early_branch_addr[20] (\early_branch_addr[20] ), .\early_branch_addr[21] (\early_branch_addr[21] ), 
            .\early_branch_addr[22] (\early_branch_addr[22] ), .\early_branch_addr[23] (\early_branch_addr[23] ), 
            .n44(n44), .\data_from_read[2] (\data_from_read[2] ), .n27294(n27294), 
            .n10(n10), .n27093(n27093), .n27277(n27277), .n23526(n23526), 
            .n22591(n22591), .n9091(n9091), .n23532(n23532), .n27306(n27306), 
            .n24742(n24742), .n24743(n24743), .n24744(n24744), .n23536(n23536), 
            .\mem_data_from_read[1] (mem_data_from_read[1]), .\mem_data_from_read[5] (mem_data_from_read[5]), 
            .\mem_data_from_read[9] (mem_data_from_read[9]), .\mem_data_from_read[13] (mem_data_from_read[13]), 
            .\data_from_read[6] (\data_from_read[6] ), .instr_fetch_running_N_945(instr_fetch_running_N_945), 
            .instr_fetch_stopped(instr_fetch_stopped), .\instr_addr[2] (instr_addr[2]), 
            .n24759(n24759), .n27268(n27268), .\mem_data_from_read[24] (mem_data_from_read[24]), 
            .\mem_data_from_read[28] (mem_data_from_read[28]), .\mem_data_from_read[26] (mem_data_from_read[26]), 
            .\mem_data_from_read[30] (mem_data_from_read[30]), .n24126(n24126), 
            .n27241(n27241), .n27255(n27255), .\qspi_data_buf[25] (qspi_data_buf[25]), 
            .\qspi_data_buf[29] (qspi_data_buf[29]), .\mem_data_from_read[17] (mem_data_from_read[17]), 
            .\mem_data_from_read[21] (mem_data_from_read[21]), .n27233(n27233), 
            .n8869(n8869), .n27279(n27279), .n23908(n23908), .n27358(n27358), 
            .n27220(n27220), .mem_op_increment_reg_de(mem_op_increment_reg_de), 
            .n27218(n27218), .\next_fsm_state_3__N_2499[3] (\next_fsm_state_3__N_2499[3] ), 
            .clk_c_enable_350(clk_c_enable_350), .clk_c_enable_367(clk_c_enable_367), 
            .\debug_branch_N_840[29] (debug_branch_N_840[29]), .\mul_out[2] (\mul_out[2] ), 
            .\mul_out[3] (\mul_out[3] ), .\mul_out[1] (\mul_out[1] ), .\ui_in_sync[1] (\ui_in_sync[1] ), 
            .n1167(n1167), .debug_rd({debug_rd}), .accum({accum}), .d_3__N_1868({d_3__N_1868}), 
            .n4577(n4577), .n26802(n26802), .n27223(n27223), .\next_accum[5] (\next_accum[5] ), 
            .\next_accum[6] (\next_accum[6] ), .\next_accum[7] (\next_accum[7] ), 
            .GND_net(GND_net), .\next_accum[8] (\next_accum[8] ), .\next_accum[9] (\next_accum[9] ), 
            .\next_accum[10] (\next_accum[10] ), .\next_accum[11] (\next_accum[11] ), 
            .\next_accum[12] (\next_accum[12] ), .\next_accum[13] (\next_accum[13] ), 
            .\next_accum[14] (\next_accum[14] ), .\next_accum[15] (\next_accum[15] ), 
            .\next_accum[16] (\next_accum[16] ), .\next_accum[17] (\next_accum[17] ), 
            .\next_accum[18] (\next_accum[18] ), .\next_accum[19] (\next_accum[19] ), 
            .\next_accum[4] (\next_accum[4] )) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(94[14] 130[6])
    
endmodule
//
// Verilog Description of module tinyqv_mem_ctrl
//

module tinyqv_mem_ctrl (clk_c, clk_c_enable_341, debug_data_continue, 
            data_txn_len, instr_data, start_instr, instr_fetch_running, 
            n27334, n23526, n27333, n23532, \instr_addr_23__N_318[0] , 
            n27255, n27327, n23536, \instr_addr_23__N_318[18] , \addr[19] , 
            \instr_addr_23__N_318[14] , \addr[15] , \qspi_data_buf[29] , 
            \qspi_data_buf[25] , \mem_data_from_read[23] , \mem_data_from_read[22] , 
            \mem_data_from_read[21] , \mem_data_from_read[20] , \mem_data_from_read[19] , 
            \mem_data_from_read[18] , \mem_data_from_read[17] , \mem_data_from_read[16] , 
            \qspi_data_buf[14] , \qspi_data_buf[12] , \qspi_data_buf[10] , 
            \qspi_data_buf[8] , \instr_addr_23__N_318[15] , \addr[16] , 
            \instr_addr_23__N_318[16] , \addr[17] , \instr_addr_23__N_318[17] , 
            \addr[18] , \instr_addr_23__N_318[6] , \addr[7] , \instr_addr_23__N_318[5] , 
            \addr[6] , \instr_addr[2] , \addr[2] , \instr_addr_23__N_318[7] , 
            \addr[8] , \instr_addr_23__N_318[3] , \addr[4] , \instr_addr_23__N_318[10] , 
            \addr[11] , data_stall, data_to_write, \instr_addr_23__N_318[9] , 
            \addr[10] , instr_fetch_stopped, \instr_addr_23__N_318[11] , 
            \addr[12] , \instr_addr_23__N_318[8] , \addr[9] , rst_reg_n, 
            \instr_addr[1] , \addr[1] , \instr_addr_23__N_318[12] , \addr[13] , 
            \instr_addr_23__N_318[22] , \addr[23] , \instr_addr_23__N_318[13] , 
            \addr[14] , \instr_addr_23__N_318[4] , \addr[5] , \next_instr_write_offset[3] , 
            \instr_addr_23__N_318[19] , \addr[20] , instr_fetch_running_N_945, 
            n27093, \instr_addr_23__N_318[20] , \addr[21] , \instr_addr_23__N_318[21] , 
            \addr[22] , mem_data_ready, n27150, n27081, is_writing_N_2331, 
            \mem_data_from_read[31] , \mem_data_from_read[27] , \mem_data_from_read[30] , 
            \mem_data_from_read[26] , \mem_data_from_read[28] , \mem_data_from_read[24] , 
            n27299, debug_stop_txn_N_2148, n27341, n23432, continue_txn_N_2131, 
            data_stall_N_2158, n27271, n27277, n27233, \pc[1] , \pc[2] , 
            n24806, n27298, debug_stop_txn_N_2147, \addr[24] , qv_data_write_n, 
            qv_data_read_n, n22591, n22344, n27356, n27357, \addr[27] , 
            \mem_data_from_read[13] , \mem_data_from_read[9] , n24743, 
            n24742, n26794, n26730, n26714, \mem_data_from_read[4] , 
            \mem_data_from_read[3] , \mem_data_from_read[5] , \mem_data_from_read[1] , 
            \mem_data_from_read[6] , n27082, \addr[0] , n27358, n27227, 
            is_writing, \instr_addr_23__N_318[2] , \addr[3] , n6930, 
            \writing_N_164[3] , n27083, qspi_ram_b_select, \qspi_data_out_3__N_5[0] , 
            qspi_ram_a_select, n24802, qspi_data_in, \fsm_state[0] , 
            n23276, clk_c_enable_358, clk_c_enable_369, n23252, clk_N_45, 
            \qspi_data_out_3__N_5[2] , n4319, n4307, \qspi_data_oe[3] , 
            clk_c_enable_346, n27080, \qspi_data_out_3__N_5[3] , \addr[20]_adj_13 , 
            \addr[22]_adj_14 , spi_clk_pos_derived_59, qspi_clk_N_56, 
            next_bit, n27210, uart_txd_N_2596, clk_c_enable_426, n24376, 
            n22303, n44, clk_c_enable_273, n805, clk_c_enable_420, 
            n27365, n22097, n4309, n26711, n5508, n5505, n22992) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output clk_c_enable_341;
    input debug_data_continue;
    output [1:0]data_txn_len;
    output [15:0]instr_data;
    input start_instr;
    input instr_fetch_running;
    input n27334;
    output n23526;
    input n27333;
    output n23532;
    input \instr_addr_23__N_318[0] ;
    output n27255;
    input n27327;
    output n23536;
    input \instr_addr_23__N_318[18] ;
    input \addr[19] ;
    input \instr_addr_23__N_318[14] ;
    input \addr[15] ;
    output \qspi_data_buf[29] ;
    output \qspi_data_buf[25] ;
    output \mem_data_from_read[23] ;
    output \mem_data_from_read[22] ;
    output \mem_data_from_read[21] ;
    output \mem_data_from_read[20] ;
    output \mem_data_from_read[19] ;
    output \mem_data_from_read[18] ;
    output \mem_data_from_read[17] ;
    output \mem_data_from_read[16] ;
    output \qspi_data_buf[14] ;
    output \qspi_data_buf[12] ;
    output \qspi_data_buf[10] ;
    output \qspi_data_buf[8] ;
    input \instr_addr_23__N_318[15] ;
    input \addr[16] ;
    input \instr_addr_23__N_318[16] ;
    input \addr[17] ;
    input \instr_addr_23__N_318[17] ;
    input \addr[18] ;
    input \instr_addr_23__N_318[6] ;
    input \addr[7] ;
    input \instr_addr_23__N_318[5] ;
    input \addr[6] ;
    input \instr_addr[2] ;
    input \addr[2] ;
    input \instr_addr_23__N_318[7] ;
    input \addr[8] ;
    input \instr_addr_23__N_318[3] ;
    input \addr[4] ;
    input \instr_addr_23__N_318[10] ;
    input \addr[11] ;
    output data_stall;
    input [31:0]data_to_write;
    input \instr_addr_23__N_318[9] ;
    input \addr[10] ;
    output instr_fetch_stopped;
    input \instr_addr_23__N_318[11] ;
    input \addr[12] ;
    input \instr_addr_23__N_318[8] ;
    input \addr[9] ;
    input rst_reg_n;
    input \instr_addr[1] ;
    input \addr[1] ;
    input \instr_addr_23__N_318[12] ;
    input \addr[13] ;
    input \instr_addr_23__N_318[22] ;
    input \addr[23] ;
    input \instr_addr_23__N_318[13] ;
    input \addr[14] ;
    input \instr_addr_23__N_318[4] ;
    input \addr[5] ;
    input \next_instr_write_offset[3] ;
    input \instr_addr_23__N_318[19] ;
    input \addr[20] ;
    output instr_fetch_running_N_945;
    input n27093;
    input \instr_addr_23__N_318[20] ;
    input \addr[21] ;
    input \instr_addr_23__N_318[21] ;
    input \addr[22] ;
    output mem_data_ready;
    output n27150;
    output n27081;
    output is_writing_N_2331;
    output \mem_data_from_read[31] ;
    output \mem_data_from_read[27] ;
    output \mem_data_from_read[30] ;
    output \mem_data_from_read[26] ;
    output \mem_data_from_read[28] ;
    output \mem_data_from_read[24] ;
    output n27299;
    output debug_stop_txn_N_2148;
    input n27341;
    output n23432;
    output continue_txn_N_2131;
    output data_stall_N_2158;
    input n27271;
    output n27277;
    input n27233;
    input \pc[1] ;
    input \pc[2] ;
    input n24806;
    input n27298;
    input debug_stop_txn_N_2147;
    input \addr[24] ;
    input [1:0]qv_data_write_n;
    input [1:0]qv_data_read_n;
    input n22591;
    input n22344;
    output n27356;
    input n27357;
    input \addr[27] ;
    output \mem_data_from_read[13] ;
    output \mem_data_from_read[9] ;
    output n24743;
    output n24742;
    output n26794;
    output n26730;
    output n26714;
    output \mem_data_from_read[4] ;
    output \mem_data_from_read[3] ;
    output \mem_data_from_read[5] ;
    output \mem_data_from_read[1] ;
    output \mem_data_from_read[6] ;
    output n27082;
    input \addr[0] ;
    input n27358;
    output n27227;
    output is_writing;
    input \instr_addr_23__N_318[2] ;
    input \addr[3] ;
    output n6930;
    output \writing_N_164[3] ;
    output n27083;
    output qspi_ram_b_select;
    input \qspi_data_out_3__N_5[0] ;
    output qspi_ram_a_select;
    input n24802;
    input [3:0]qspi_data_in;
    output \fsm_state[0] ;
    output n23276;
    input clk_c_enable_358;
    input clk_c_enable_369;
    output n23252;
    input clk_N_45;
    input \qspi_data_out_3__N_5[2] ;
    output n4319;
    output n4307;
    output \qspi_data_oe[3] ;
    input clk_c_enable_346;
    output n27080;
    input \qspi_data_out_3__N_5[3] ;
    output \addr[20]_adj_13 ;
    output \addr[22]_adj_14 ;
    output spi_clk_pos_derived_59;
    output qspi_clk_N_56;
    input next_bit;
    input n27210;
    input uart_txd_N_2596;
    output clk_c_enable_426;
    input n24376;
    input n22303;
    input n44;
    output clk_c_enable_273;
    input n805;
    output clk_c_enable_420;
    output n27365;
    output n22097;
    output n4309;
    output n26711;
    output n5508;
    output n5505;
    output n22992;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    
    wire continue_txn, clk_c_enable_5, qspi_write_done, n9653, n27301, 
        clk_c_enable_279, n22180, clk_c_enable_206;
    wire [31:0]instr_data_7__N_1969;
    wire [1:0]qspi_data_byte_idx;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(59[15:33])
    
    wire clk_c_enable_291, qspi_data_byte_idx_1__N_2025, n9, instr_active, 
        clk_c_enable_79, instr_active_N_2106, qspi_data_ready, n27307;
    wire [24:0]addr_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(57[17:24])
    wire [31:0]qspi_data_buf;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(58[16:29])
    
    wire clk_c_enable_183, clk_c_enable_191, clk_c_enable_199, debug_stall_txn, 
        n27105, n27310, n1055, n9624, n27375;
    wire [1:0]read_cycles_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(105[15:32])
    
    wire n27100, n6942, debug_stop_txn_N_2119, n5423, n27087, n22307, 
        n8804;
    wire [1:0]data_txn_len_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(49[15:27])
    
    wire n27265, n27217, ram_b_block_N_2303, ram_a_block_N_2299, n27251, 
        n23418, n482, n9702, clk_c_enable_392;
    wire [1:0]n174;
    
    wire debug_stop_txn_N_2145, n27360, data_ready_N_2108, n27254, data_ready_N_2113, 
        n27273, n24390, n27361;
    wire [1:0]write_qspi_data_byte_idx_1__N_2021;
    
    wire data_ready_N_2112, n22387, debug_stop_txn_N_2142, n27324, n9276, 
        n27325, debug_stop_txn_N_2120, n23438, n28559, n24701, n24704, 
        n24707, n24710, n24697, n24694, n24691, n26951, n26945, 
        n26939, n26130, n24688, n24700, n24703, n24706, n24709, 
        n27344, n27345, n23258, last_ram_b_sel, n27352, n27272;
    wire [1:0]txn_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(56[16:23])
    
    wire n45, spi_ram_a_select_N_2309, spi_ram_b_select_N_2313, n27090, 
        n23424;
    wire [23:0]addr_23__N_2188;
    
    wire n27232, n27250, n5909, spi_clk_pos, stop_txn_now_N_2363;
    
    FD1P3IX continue_txn_187 (.D(debug_data_continue), .SP(clk_c_enable_5), 
            .CD(clk_c_enable_341), .CK(clk_c), .Q(continue_txn)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam continue_txn_187.GSR = "DISABLED";
    FD1S3IX qspi_write_done_185 (.D(n27301), .CK(clk_c), .CD(n9653), .Q(qspi_write_done)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(173[12] 175[8])
    defparam qspi_write_done_185.GSR = "DISABLED";
    FD1P3AX data_txn_len_i0_i0 (.D(n22180), .SP(clk_c_enable_279), .CK(clk_c), 
            .Q(data_txn_len[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(177[12] 183[8])
    defparam data_txn_len_i0_i0.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i1 (.D(instr_data_7__N_1969[0]), .SP(clk_c_enable_206), 
            .CK(clk_c), .Q(instr_data[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i1.GSR = "DISABLED";
    FD1P3IX qspi_data_byte_idx__i0 (.D(n9), .SP(clk_c_enable_291), .CD(qspi_data_byte_idx_1__N_2025), 
            .CK(clk_c), .Q(qspi_data_byte_idx[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam qspi_data_byte_idx__i0.GSR = "DISABLED";
    FD1P3IX instr_active_180 (.D(start_instr), .SP(clk_c_enable_79), .CD(instr_active_N_2106), 
            .CK(clk_c), .Q(instr_active)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(103[12] 109[8])
    defparam instr_active_180.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(qspi_data_ready), .B(n27307), .C(instr_fetch_running), 
         .D(n27334), .Z(n23526)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(65[22:102])
    defparam i1_2_lut_4_lut.init = 16'hff7f;
    LUT4 i1_2_lut_4_lut_adj_471 (.A(qspi_data_ready), .B(n27307), .C(instr_fetch_running), 
         .D(n27333), .Z(n23532)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(65[22:102])
    defparam i1_2_lut_4_lut_adj_471.init = 16'hff7f;
    LUT4 i4134_2_lut_rep_630_4_lut (.A(qspi_data_ready), .B(n27307), .C(instr_fetch_running), 
         .D(\instr_addr_23__N_318[0] ), .Z(n27255)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(65[22:102])
    defparam i4134_2_lut_rep_630_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_472 (.A(qspi_data_ready), .B(n27307), .C(instr_fetch_running), 
         .D(n27327), .Z(n23536)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(65[22:102])
    defparam i1_2_lut_4_lut_adj_472.init = 16'hff7f;
    LUT4 data_addr_24__I_0_i20_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[18] ), .D(\addr[19] ), .Z(addr_in[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i20_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX qspi_data_buf_i32 (.D(instr_data_7__N_1969[31]), .SP(clk_c_enable_183), 
            .CK(clk_c), .Q(qspi_data_buf[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i32.GSR = "DISABLED";
    LUT4 data_addr_24__I_0_i16_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[14] ), .D(\addr[15] ), .Z(addr_in[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i16_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX qspi_data_buf_i31 (.D(instr_data_7__N_1969[30]), .SP(clk_c_enable_183), 
            .CK(clk_c), .Q(qspi_data_buf[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i31.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i30 (.D(instr_data_7__N_1969[29]), .SP(clk_c_enable_183), 
            .CK(clk_c), .Q(\qspi_data_buf[29] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i30.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i29 (.D(instr_data_7__N_1969[28]), .SP(clk_c_enable_183), 
            .CK(clk_c), .Q(qspi_data_buf[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i29.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i28 (.D(instr_data_7__N_1969[27]), .SP(clk_c_enable_183), 
            .CK(clk_c), .Q(qspi_data_buf[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i28.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i27 (.D(instr_data_7__N_1969[26]), .SP(clk_c_enable_183), 
            .CK(clk_c), .Q(qspi_data_buf[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i27.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i26 (.D(instr_data_7__N_1969[25]), .SP(clk_c_enable_183), 
            .CK(clk_c), .Q(\qspi_data_buf[25] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i26.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i25 (.D(instr_data_7__N_1969[24]), .SP(clk_c_enable_183), 
            .CK(clk_c), .Q(qspi_data_buf[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i25.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i24 (.D(instr_data_7__N_1969[23]), .SP(clk_c_enable_191), 
            .CK(clk_c), .Q(\mem_data_from_read[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i24.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i23 (.D(instr_data_7__N_1969[22]), .SP(clk_c_enable_191), 
            .CK(clk_c), .Q(\mem_data_from_read[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i23.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i22 (.D(instr_data_7__N_1969[21]), .SP(clk_c_enable_191), 
            .CK(clk_c), .Q(\mem_data_from_read[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i22.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i21 (.D(instr_data_7__N_1969[20]), .SP(clk_c_enable_191), 
            .CK(clk_c), .Q(\mem_data_from_read[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i21.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i20 (.D(instr_data_7__N_1969[19]), .SP(clk_c_enable_191), 
            .CK(clk_c), .Q(\mem_data_from_read[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i20.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i19 (.D(instr_data_7__N_1969[18]), .SP(clk_c_enable_191), 
            .CK(clk_c), .Q(\mem_data_from_read[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i19.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i18 (.D(instr_data_7__N_1969[17]), .SP(clk_c_enable_191), 
            .CK(clk_c), .Q(\mem_data_from_read[17] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i18.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i17 (.D(instr_data_7__N_1969[16]), .SP(clk_c_enable_191), 
            .CK(clk_c), .Q(\mem_data_from_read[16] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i17.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i16 (.D(instr_data_7__N_1969[15]), .SP(clk_c_enable_199), 
            .CK(clk_c), .Q(qspi_data_buf[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i16.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i15 (.D(instr_data_7__N_1969[14]), .SP(clk_c_enable_199), 
            .CK(clk_c), .Q(\qspi_data_buf[14] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i15.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i14 (.D(instr_data_7__N_1969[13]), .SP(clk_c_enable_199), 
            .CK(clk_c), .Q(qspi_data_buf[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i14.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i13 (.D(instr_data_7__N_1969[12]), .SP(clk_c_enable_199), 
            .CK(clk_c), .Q(\qspi_data_buf[12] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i13.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i12 (.D(instr_data_7__N_1969[11]), .SP(clk_c_enable_199), 
            .CK(clk_c), .Q(qspi_data_buf[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i12.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i11 (.D(instr_data_7__N_1969[10]), .SP(clk_c_enable_199), 
            .CK(clk_c), .Q(\qspi_data_buf[10] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i11.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i10 (.D(instr_data_7__N_1969[9]), .SP(clk_c_enable_199), 
            .CK(clk_c), .Q(qspi_data_buf[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i10.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i9 (.D(instr_data_7__N_1969[8]), .SP(clk_c_enable_199), 
            .CK(clk_c), .Q(\qspi_data_buf[8] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i9.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i8 (.D(instr_data_7__N_1969[7]), .SP(clk_c_enable_206), 
            .CK(clk_c), .Q(instr_data[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i8.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i7 (.D(instr_data_7__N_1969[6]), .SP(clk_c_enable_206), 
            .CK(clk_c), .Q(instr_data[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i7.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i6 (.D(instr_data_7__N_1969[5]), .SP(clk_c_enable_206), 
            .CK(clk_c), .Q(instr_data[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i6.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i5 (.D(instr_data_7__N_1969[4]), .SP(clk_c_enable_206), 
            .CK(clk_c), .Q(instr_data[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i5.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i4 (.D(instr_data_7__N_1969[3]), .SP(clk_c_enable_206), 
            .CK(clk_c), .Q(instr_data[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i4.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i3 (.D(instr_data_7__N_1969[2]), .SP(clk_c_enable_206), 
            .CK(clk_c), .Q(instr_data[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i3.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i2 (.D(instr_data_7__N_1969[1]), .SP(clk_c_enable_206), 
            .CK(clk_c), .Q(instr_data[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i2.GSR = "DISABLED";
    LUT4 data_addr_24__I_0_i17_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[15] ), .D(\addr[16] ), .Z(addr_in[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i18_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[16] ), .D(\addr[17] ), .Z(addr_in[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i19_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[17] ), .D(\addr[18] ), .Z(addr_in[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i8_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[6] ), .D(\addr[7] ), .Z(addr_in[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i7_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[5] ), .D(\addr[6] ), .Z(addr_in[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i3_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr[2] ), .D(\addr[2] ), .Z(addr_in[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i9_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[7] ), .D(\addr[8] ), .Z(addr_in[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr_23__N_318[3] ), 
         .D(\addr[4] ), .Z(addr_in[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i12_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[10] ), .D(\addr[11] ), .Z(addr_in[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 debug_stall_txn_I_0_2_lut_rep_480 (.A(debug_stall_txn), .B(data_stall), 
         .Z(n27105)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(129[20:43])
    defparam debug_stall_txn_I_0_2_lut_rep_480.init = 16'heeee;
    LUT4 i7217_3_lut_4_lut (.A(debug_stall_txn), .B(data_stall), .C(n27310), 
         .D(n1055), .Z(n9624)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(129[20:43])
    defparam i7217_3_lut_4_lut.init = 16'hefe0;
    LUT4 instr_data_7__I_173_i10_4_lut (.A(data_to_write[9]), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n27375), .Z(instr_data_7__N_1969[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i10_4_lut.init = 16'h0aca;
    LUT4 i12362_2_lut_rep_475_3_lut (.A(debug_stall_txn), .B(data_stall), 
         .C(read_cycles_count[1]), .Z(n27100)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(129[20:43])
    defparam i12362_2_lut_rep_475_3_lut.init = 16'hfefe;
    LUT4 data_addr_24__I_0_i11_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[9] ), .D(\addr[10] ), .Z(addr_in[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i11_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX instr_fetch_stopped_182 (.D(debug_stop_txn_N_2119), .CK(clk_c), 
            .CD(n6942), .Q(instr_fetch_stopped)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam instr_fetch_stopped_182.GSR = "DISABLED";
    LUT4 data_addr_24__I_0_i13_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[11] ), .D(\addr[12] ), .Z(addr_in[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr_23__N_318[8] ), 
         .D(\addr[9] ), .Z(addr_in[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3412_2_lut (.A(continue_txn), .B(rst_reg_n), .Z(n5423)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i3412_2_lut.init = 16'h4444;
    LUT4 data_addr_24__I_0_i2_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr[1] ), .D(\addr[1] ), .Z(addr_in[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i14_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[12] ), .D(\addr[13] ), .Z(addr_in[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i24_3_lut_rep_462_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[22] ), .D(\addr[23] ), .Z(n27087)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i24_3_lut_rep_462_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i15_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[13] ), .D(\addr[14] ), .Z(addr_in[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i18_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr_23__N_318[4] ), 
         .D(\addr[5] ), .Z(addr_in[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut (.A(n22307), .B(\next_instr_write_offset[3] ), .C(n27307), 
         .D(qspi_data_ready), .Z(debug_stall_txn)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut.init = 16'h0040;
    LUT4 data_addr_24__I_0_i21_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[19] ), .D(\addr[20] ), .Z(addr_in[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i21_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX instr_fetch_started_181 (.D(n27093), .CK(clk_c), .CD(n8804), 
            .Q(instr_fetch_running_N_945)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam instr_fetch_started_181.GSR = "DISABLED";
    LUT4 data_addr_24__I_0_i22_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[20] ), .D(\addr[21] ), .Z(addr_in[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 instr_data_7__I_173_i9_4_lut (.A(data_to_write[8]), .B(instr_data[8]), 
         .C(qspi_data_ready), .D(n27375), .Z(instr_data_7__N_1969[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i9_4_lut.init = 16'h0aca;
    LUT4 data_addr_24__I_0_i23_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[21] ), .D(\addr[22] ), .Z(addr_in[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_525 (.A(mem_data_ready), .B(data_txn_len_c[1]), .Z(n27150)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_525.init = 16'h2222;
    FD1P3AX data_txn_len_i0_i1 (.D(n27265), .SP(clk_c_enable_279), .CK(clk_c), 
            .Q(data_txn_len_c[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(177[12] 183[8])
    defparam data_txn_len_i0_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_456_3_lut_4_lut (.A(n27217), .B(start_instr), .C(ram_b_block_N_2303), 
         .D(ram_a_block_N_2299), .Z(n27081)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i1_2_lut_rep_456_3_lut_4_lut.init = 16'hd000;
    LUT4 i1_4_lut_3_lut (.A(start_instr), .B(n27251), .C(n23418), .Z(is_writing_N_2331)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_4_lut_3_lut.init = 16'h4040;
    LUT4 qspi_data_buf_31__I_0_189_3_lut (.A(qspi_data_buf[31]), .B(instr_data[15]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[31] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_31__I_0_189_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_27__I_0_3_lut (.A(qspi_data_buf[27]), .B(instr_data[11]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[27] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_27__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_30__I_0_3_lut (.A(qspi_data_buf[30]), .B(instr_data[14]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[30] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_30__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_26__I_0_3_lut (.A(qspi_data_buf[26]), .B(instr_data[10]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[26] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_26__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_28__I_0_3_lut (.A(qspi_data_buf[28]), .B(instr_data[12]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[28] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_28__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_24__I_0_3_lut (.A(qspi_data_buf[24]), .B(instr_data[8]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_24__I_0_3_lut.init = 16'hcaca;
    LUT4 i7355_2_lut_3_lut_4_lut (.A(n27217), .B(start_instr), .C(n482), 
         .D(n27299), .Z(n9702)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i7355_2_lut_3_lut_4_lut.init = 16'hf020;
    LUT4 debug_stop_txn_I_194_2_lut (.A(instr_fetch_running_N_945), .B(debug_stall_txn), 
         .Z(debug_stop_txn_N_2148)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(78[44:79])
    defparam debug_stop_txn_I_194_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n27217), .B(start_instr), .C(n482), 
         .D(n27299), .Z(clk_c_enable_392)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf0fd;
    FD1P3IX qspi_data_byte_idx__i1 (.D(n174[1]), .SP(clk_c_enable_291), 
            .CD(qspi_data_byte_idx_1__N_2025), .CK(clk_c), .Q(qspi_data_byte_idx[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam qspi_data_byte_idx__i1.GSR = "DISABLED";
    LUT4 debug_stop_txn_I_193_4_lut (.A(qspi_data_ready), .B(n22307), .C(n27375), 
         .D(\next_instr_write_offset[3] ), .Z(debug_stop_txn_N_2145)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[30:99])
    defparam debug_stop_txn_I_193_4_lut.init = 16'h3b0a;
    LUT4 i1_2_lut_4_lut_adj_473 (.A(qspi_data_ready), .B(n27307), .C(instr_fetch_running), 
         .D(n27341), .Z(n23432)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(65[22:102])
    defparam i1_2_lut_4_lut_adj_473.init = 16'h8000;
    LUT4 instr_data_7__I_173_i8_3_lut (.A(data_to_write[7]), .B(instr_data[15]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i8_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i7_3_lut (.A(data_to_write[6]), .B(instr_data[14]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i7_3_lut.init = 16'hcaca;
    LUT4 qspi_data_ready_I_0_202_2_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(n27360), 
         .C(data_txn_len[0]), .D(qspi_data_ready), .Z(data_ready_N_2108)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[64:98])
    defparam qspi_data_ready_I_0_202_2_lut_4_lut.init = 16'h2100;
    LUT4 i4132_2_lut_rep_629_4_lut (.A(qspi_data_ready), .B(n27307), .C(instr_fetch_running), 
         .D(\instr_addr_23__N_318[0] ), .Z(n27254)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(65[22:102])
    defparam i4132_2_lut_rep_629_4_lut.init = 16'h7f80;
    LUT4 i4676_4_lut (.A(n27217), .B(continue_txn_N_2131), .C(continue_txn), 
         .D(data_stall_N_2158), .Z(clk_c_enable_5)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(198[22] 203[16])
    defparam i4676_4_lut.init = 16'h05c5;
    LUT4 data_ready_N_2113_I_0_4_lut (.A(data_ready_N_2113), .B(n27273), 
         .C(n27271), .D(mem_data_ready), .Z(continue_txn_N_2131)) /* synthesis lut_function=(!((B (C)+!B (C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(194[30:139])
    defparam data_ready_N_2113_I_0_4_lut.init = 16'h0a2a;
    LUT4 continue_txn_I_189_4_lut (.A(n24390), .B(data_ready_N_2108), .C(n27361), 
         .D(data_txn_len_c[1]), .Z(data_stall_N_2158)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(190[21] 191[76])
    defparam continue_txn_I_189_4_lut.init = 16'hecce;
    LUT4 i1_3_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(data_txn_len[0]), .Z(n24390)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4848;
    LUT4 instr_data_7__I_173_i6_3_lut (.A(data_to_write[5]), .B(instr_data[13]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i6_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_652_4_lut (.A(n27375), .B(instr_active), .C(instr_fetch_running), 
         .D(qspi_data_ready), .Z(n27277)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(65[22:102])
    defparam i1_3_lut_rep_652_4_lut.init = 16'h4000;
    LUT4 i20088_4_lut (.A(n27254), .B(n27233), .C(\pc[1] ), .D(\pc[2] ), 
         .Z(n22307)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i20088_4_lut.init = 16'h7bde;
    LUT4 data_ready_I_0_206_4_lut (.A(instr_active), .B(data_ready_N_2108), 
         .C(n27271), .D(data_ready_N_2112), .Z(mem_data_ready)) /* synthesis lut_function=(!(A+!(B+!(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[25:190])
    defparam data_ready_I_0_206_4_lut.init = 16'h4544;
    FD1P3IX data_stall_188 (.D(n24806), .SP(rst_reg_n), .CD(n5423), .CK(clk_c), 
            .Q(data_stall)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam data_stall_188.GSR = "DISABLED";
    LUT4 instr_data_7__I_173_i5_3_lut (.A(data_to_write[4]), .B(instr_data[12]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i5_3_lut.init = 16'hcaca;
    LUT4 i12177_4_lut (.A(n27298), .B(debug_stop_txn_N_2147), .C(debug_stop_txn_N_2145), 
         .D(n22387), .Z(debug_stop_txn_N_2142)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[26] 86[20])
    defparam i12177_4_lut.init = 16'hccdc;
    LUT4 i105_2_lut_rep_699 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n27324)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i105_2_lut_rep_699.init = 16'hbbbb;
    LUT4 i23677_2_lut_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n9276), .D(qspi_data_ready), .Z(clk_c_enable_191)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C)+!B !((D)+!C)))) */ ;
    defparam i23677_2_lut_3_lut_4_lut.init = 16'h40f0;
    LUT4 i12772_2_lut_rep_700 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n27325)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12772_2_lut_rep_700.init = 16'h8888;
    LUT4 i23675_2_lut_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n9276), .D(qspi_data_ready), .Z(clk_c_enable_183)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i23675_2_lut_3_lut_4_lut.init = 16'h80f0;
    PFUMX debug_stop_txn_I_182 (.BLUT(debug_stop_txn_N_2120), .ALUT(debug_stop_txn_N_2142), 
          .C0(instr_active), .Z(debug_stop_txn_N_2119)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;
    LUT4 i1_2_lut_3_lut (.A(qspi_data_ready), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(rst_reg_n), .Z(n23438)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[26:60])
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut (.A(instr_active), .B(\addr[24] ), .Z(n23418)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 instr_active_I_0_2_lut_rep_755 (.A(instr_active), .B(start_instr), 
         .Z(n28559)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam instr_active_I_0_2_lut_rep_755.init = 16'heeee;
    LUT4 i22358_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[28]), .D(\mem_data_from_read[20] ), .Z(n24701)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22358_3_lut_4_lut.init = 16'hf960;
    LUT4 i22361_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[29] ), .D(\mem_data_from_read[21] ), .Z(n24704)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22361_3_lut_4_lut.init = 16'hf960;
    LUT4 i22364_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[30]), .D(\mem_data_from_read[22] ), .Z(n24707)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22364_3_lut_4_lut.init = 16'hf960;
    LUT4 i22367_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[31]), .D(\mem_data_from_read[23] ), .Z(n24710)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22367_3_lut_4_lut.init = 16'hf960;
    LUT4 i22354_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[11]), .D(instr_data[3]), .Z(n24697)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22354_3_lut_4_lut.init = 16'hf960;
    LUT4 i22351_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[10] ), .D(instr_data[2]), .Z(n24694)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22351_3_lut_4_lut.init = 16'hf960;
    LUT4 i22348_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[9]), .D(instr_data[1]), .Z(n24691)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22348_3_lut_4_lut.init = 16'hf960;
    LUT4 n5072_bdd_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[25] ), .D(\mem_data_from_read[17] ), .Z(n26951)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n5072_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 n15156_bdd_3_lut_24318_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[26]), .D(\mem_data_from_read[18] ), .Z(n26945)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n15156_bdd_3_lut_24318_4_lut.init = 16'hf960;
    LUT4 n15156_bdd_3_lut_24255_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[27]), .D(\mem_data_from_read[19] ), .Z(n26939)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n15156_bdd_3_lut_24255_4_lut.init = 16'hf960;
    LUT4 n15156_bdd_3_lut_23902_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[24]), .D(\mem_data_from_read[16] ), .Z(n26130)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n15156_bdd_3_lut_23902_4_lut.init = 16'hf960;
    LUT4 i22345_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[8] ), .D(instr_data[0]), .Z(n24688)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22345_3_lut_4_lut.init = 16'hf960;
    LUT4 i22357_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[12] ), .D(instr_data[4]), .Z(n24700)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22357_3_lut_4_lut.init = 16'hf960;
    LUT4 i22360_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[13]), .D(instr_data[5]), .Z(n24703)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22360_3_lut_4_lut.init = 16'hf960;
    LUT4 i22363_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[14] ), .D(instr_data[6]), .Z(n24706)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22363_3_lut_4_lut.init = 16'hf960;
    LUT4 i22366_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[15]), .D(instr_data[7]), .Z(n24709)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i22366_3_lut_4_lut.init = 16'hf960;
    LUT4 i4873_2_lut_rep_719 (.A(qv_data_write_n[1]), .B(qv_data_read_n[1]), 
         .Z(n27344)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(73[22:48])
    defparam i4873_2_lut_rep_719.init = 16'h8888;
    LUT4 i4665_2_lut_rep_720 (.A(qv_data_write_n[0]), .B(qv_data_read_n[0]), 
         .Z(n27345)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(73[22:48])
    defparam i4665_2_lut_rep_720.init = 16'h8888;
    LUT4 i20167_2_lut_3_lut_4_lut (.A(qv_data_write_n[0]), .B(qv_data_read_n[0]), 
         .C(qv_data_read_n[1]), .D(qv_data_write_n[1]), .Z(n22387)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(73[22:48])
    defparam i20167_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_474 (.A(start_instr), .B(n27087), .C(\addr[24] ), 
         .D(n23258), .Z(ram_b_block_N_2303)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_4_lut_adj_474.init = 16'hffbf;
    LUT4 i1_2_lut_adj_475 (.A(instr_active), .B(last_ram_b_sel), .Z(n23258)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_2_lut_adj_475.init = 16'heeee;
    LUT4 instr_data_7__I_173_i1_3_lut (.A(data_to_write[0]), .B(instr_data[8]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i1_3_lut.init = 16'hcaca;
    LUT4 qspi_data_byte_idx_1__I_0_i3_2_lut_rep_727 (.A(qspi_data_byte_idx[0]), 
         .B(qspi_data_byte_idx[1]), .Z(n27352)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[144:171])
    defparam qspi_data_byte_idx_1__I_0_i3_2_lut_rep_727.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_476 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n9276), .D(qspi_data_ready), .Z(clk_c_enable_206)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[144:171])
    defparam i1_2_lut_3_lut_4_lut_adj_476.init = 16'h10f0;
    LUT4 data_stall_I_0_213_2_lut_3_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(data_stall), .Z(data_ready_N_2113)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[144:171])
    defparam data_stall_I_0_213_2_lut_3_lut.init = 16'h1010;
    LUT4 i23660_4_lut (.A(n23438), .B(n27272), .C(n22591), .D(n22344), 
         .Z(clk_c_enable_291)) /* synthesis lut_function=(!(A (B+(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(149[13:62])
    defparam i23660_4_lut.init = 16'h5777;
    LUT4 i12183_2_lut_rep_731 (.A(qv_data_read_n[0]), .B(qv_data_read_n[1]), 
         .Z(n27356)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12183_2_lut_rep_731.init = 16'h8888;
    LUT4 i12803_2_lut_rep_648_3_lut_4_lut (.A(qv_data_read_n[0]), .B(qv_data_read_n[1]), 
         .C(n27357), .D(\addr[27] ), .Z(n27273)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i12803_2_lut_rep_648_3_lut_4_lut.init = 16'hfff8;
    LUT4 i3791_2_lut_rep_736 (.A(qspi_data_byte_idx[1]), .B(qspi_data_byte_idx[0]), 
         .Z(n27361)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(153[39:65])
    defparam i3791_2_lut_rep_736.init = 16'h6666;
    LUT4 i1_4_lut_4_lut (.A(qspi_data_byte_idx[1]), .B(qspi_data_byte_idx[0]), 
         .C(txn_len[0]), .D(n45), .Z(n174[1])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(153[39:65])
    defparam i1_4_lut_4_lut.init = 16'h6624;
    LUT4 i1_4_lut_adj_477 (.A(start_instr), .B(n27087), .C(\addr[24] ), 
         .D(instr_active), .Z(spi_ram_a_select_N_2309)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_4_lut_adj_477.init = 16'hffef;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\addr[24] ), .D(\addr[23] ), .Z(spi_ram_b_select_N_2313)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hefff;
    LUT4 i1_4_lut_adj_478 (.A(n27090), .B(start_instr), .C(n27299), .D(n23424), 
         .Z(addr_23__N_2188[0])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_478.init = 16'h0200;
    LUT4 i1_3_lut_4_lut_4_lut (.A(continue_txn), .B(n27301), .C(write_qspi_data_byte_idx_1__N_2021[0]), 
         .D(qspi_data_ready), .Z(debug_stop_txn_N_2120)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[102:115])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 qspi_data_byte_idx_1__I_0_197_i3_2_lut_rep_750 (.A(qspi_data_byte_idx[0]), 
         .B(qspi_data_byte_idx[1]), .Z(n27375)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam qspi_data_byte_idx_1__I_0_197_i3_2_lut_rep_750.init = 16'hdddd;
    LUT4 i1_2_lut_rep_682_3_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(instr_active), .Z(n27307)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam i1_2_lut_rep_682_3_lut.init = 16'h2020;
    LUT4 i23639_2_lut_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n9276), .D(qspi_data_ready), .Z(clk_c_enable_199)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam i23639_2_lut_3_lut_4_lut.init = 16'h20f0;
    LUT4 instr_data_7__I_173_i32_3_lut (.A(data_to_write[31]), .B(instr_data[15]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i32_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i31_3_lut (.A(data_to_write[30]), .B(instr_data[14]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i31_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i30_3_lut (.A(data_to_write[29]), .B(instr_data[13]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i30_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i29_3_lut (.A(data_to_write[28]), .B(instr_data[12]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i29_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i28_3_lut (.A(data_to_write[27]), .B(instr_data[11]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i28_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i25_4_lut (.A(data_to_write[24]), .B(instr_data[8]), 
         .C(qspi_data_ready), .D(n27325), .Z(instr_data_7__N_1969[24])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i25_4_lut.init = 16'hca0a;
    LUT4 instr_data_7__I_173_i24_3_lut (.A(data_to_write[23]), .B(instr_data[15]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i24_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i23_3_lut (.A(data_to_write[22]), .B(instr_data[14]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i23_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i22_3_lut (.A(data_to_write[21]), .B(instr_data[13]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i22_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i21_3_lut (.A(data_to_write[20]), .B(instr_data[12]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i21_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i20_3_lut (.A(data_to_write[19]), .B(instr_data[11]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i20_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i19_4_lut (.A(data_to_write[18]), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n27324), .Z(instr_data_7__N_1969[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i19_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i18_4_lut (.A(data_to_write[17]), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n27324), .Z(instr_data_7__N_1969[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i18_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i17_4_lut (.A(data_to_write[16]), .B(instr_data[8]), 
         .C(qspi_data_ready), .D(n27324), .Z(instr_data_7__N_1969[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i17_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i16_3_lut (.A(data_to_write[15]), .B(instr_data[15]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i16_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i15_3_lut (.A(data_to_write[14]), .B(instr_data[14]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i15_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i11_4_lut (.A(data_to_write[10]), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n27375), .Z(instr_data_7__N_1969[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i11_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i12_3_lut (.A(data_to_write[11]), .B(instr_data[11]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i12_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i14_3_lut (.A(data_to_write[13]), .B(instr_data[13]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i14_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i13_3_lut (.A(data_to_write[12]), .B(instr_data[12]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i13_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i4_4_lut (.A(data_to_write[3]), .B(instr_data[11]), 
         .C(qspi_data_ready), .D(n27352), .Z(instr_data_7__N_1969[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i4_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i3_4_lut (.A(data_to_write[2]), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n27352), .Z(instr_data_7__N_1969[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i3_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i2_4_lut (.A(data_to_write[1]), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n27352), .Z(instr_data_7__N_1969[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i2_4_lut.init = 16'h0aca;
    LUT4 qspi_data_buf_15__I_0_i6_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), 
         .C(instr_data[13]), .D(qspi_data_buf[13]), .Z(\mem_data_from_read[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam qspi_data_buf_15__I_0_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 qspi_data_buf_15__I_0_i2_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), 
         .C(instr_data[9]), .D(qspi_data_buf[9]), .Z(\mem_data_from_read[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam qspi_data_buf_15__I_0_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i22400_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), .C(instr_data[15]), 
         .D(qspi_data_buf[15]), .Z(n24743)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i22400_3_lut_4_lut.init = 16'hf780;
    LUT4 i22399_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), .C(instr_data[11]), 
         .D(qspi_data_buf[11]), .Z(n24742)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i22399_3_lut_4_lut.init = 16'hf780;
    LUT4 n5057_bdd_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), .C(instr_data[15]), 
         .D(instr_data[7]), .Z(n26794)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n5057_bdd_3_lut_4_lut.init = 16'hfb40;
    LUT4 mem_data_from_read_4__bdd_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), 
         .C(instr_data[8]), .D(instr_data[0]), .Z(n26730)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mem_data_from_read_4__bdd_3_lut_4_lut.init = 16'hfb40;
    LUT4 mem_data_from_read_6__bdd_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), 
         .C(instr_data[10]), .D(instr_data[2]), .Z(n26714)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mem_data_from_read_6__bdd_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i5_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), 
         .C(instr_data[12]), .D(instr_data[4]), .Z(\mem_data_from_read[4] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_adj_479 (.A(instr_active), .B(start_instr), .C(data_txn_len[0]), 
         .Z(txn_len[0])) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_3_lut_adj_479.init = 16'hfefe;
    LUT4 instr_data_7__I_0_i4_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), 
         .C(instr_data[11]), .D(instr_data[3]), .Z(\mem_data_from_read[3] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i6_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), 
         .C(instr_data[13]), .D(instr_data[5]), .Z(\mem_data_from_read[5] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i2_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), 
         .C(instr_data[9]), .D(instr_data[1]), .Z(\mem_data_from_read[1] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i7_3_lut_4_lut (.A(data_txn_len[0]), .B(n27150), 
         .C(instr_data[14]), .D(instr_data[6]), .Z(\mem_data_from_read[6] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_457_3_lut_4_lut (.A(n27251), .B(n27232), .C(ram_a_block_N_2299), 
         .D(start_instr), .Z(n27082)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_rep_457_3_lut_4_lut.init = 16'hf070;
    LUT4 i12383_2_lut_rep_626_3_lut_4_lut (.A(n27298), .B(n27356), .C(qspi_write_done), 
         .D(n27299), .Z(n27251)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12383_2_lut_rep_626_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_480 (.A(n27271), .B(n27250), .C(n23418), 
         .D(n27093), .Z(addr_in[24])) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(95[18] 98[33])
    defparam i1_2_lut_3_lut_4_lut_adj_480.init = 16'hd0f0;
    LUT4 i1_2_lut_adj_481 (.A(instr_active), .B(\addr[0] ), .Z(n23424)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_481.init = 16'h4444;
    LUT4 i3770_2_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .Z(n5909)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i3770_2_lut.init = 16'h8888;
    LUT4 i23447_2_lut_3_lut_4_lut (.A(n27271), .B(n27250), .C(rst_reg_n), 
         .D(n27251), .Z(clk_c_enable_279)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam i23447_2_lut_3_lut_4_lut.init = 16'h1fff;
    LUT4 i1_2_lut_rep_465_3_lut_4_lut (.A(n27271), .B(n27250), .C(start_instr), 
         .D(n27251), .Z(n27090)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam i1_2_lut_rep_465_3_lut_4_lut.init = 16'hf1ff;
    LUT4 i1_4_lut_4_lut_adj_482 (.A(n27271), .B(n27250), .C(data_stall), 
         .D(qspi_data_ready), .Z(n9276)) /* synthesis lut_function=(A (D)+!A ((C+(D))+!B)) */ ;
    defparam i1_4_lut_4_lut_adj_482.init = 16'hff51;
    LUT4 i1_2_lut_rep_625_3_lut_4_lut (.A(n27298), .B(n27356), .C(qspi_write_done), 
         .D(n27299), .Z(n27250)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;
    defparam i1_2_lut_rep_625_3_lut_4_lut.init = 16'hfff1;
    LUT4 i1_2_lut_rep_602_3_lut_4_lut_4_lut (.A(n27298), .B(n27356), .C(n27272), 
         .D(n27358), .Z(n27227)) /* synthesis lut_function=(A (C)+!A ((C+!(D))+!B)) */ ;
    defparam i1_2_lut_rep_602_3_lut_4_lut_4_lut.init = 16'hf1f5;
    LUT4 i1_2_lut_rep_607_3_lut_4_lut_4_lut (.A(n27298), .B(n27356), .C(n27272), 
         .D(n27358), .Z(n27232)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_2_lut_rep_607_3_lut_4_lut_4_lut.init = 16'hfffb;
    LUT4 i12806_2_lut_rep_592_3_lut_4_lut_3_lut_4_lut_4_lut (.A(n27298), .B(n27356), 
         .C(n27272), .D(n27358), .Z(n27217)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i12806_2_lut_rep_592_3_lut_4_lut_3_lut_4_lut_4_lut.init = 16'hfefa;
    LUT4 data_ready_I_178_2_lut_3_lut_4_lut (.A(n27272), .B(n27273), .C(data_ready_N_2113), 
         .D(n27271), .Z(data_ready_N_2112)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(95[18] 98[33])
    defparam data_ready_I_178_2_lut_3_lut_4_lut.init = 16'hf0f4;
    LUT4 i1_4_lut_adj_483 (.A(n27272), .B(debug_stop_txn_N_2119), .C(is_writing), 
         .D(spi_clk_pos), .Z(stop_txn_now_N_2363)) /* synthesis lut_function=(A (B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(91[18] 99[12])
    defparam i1_4_lut_adj_483.init = 16'h8808;
    LUT4 data_addr_24__I_0_i4_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[2] ), .D(\addr[3] ), .Z(addr_in[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i4_3_lut_4_lut.init = 16'hf1e0;
    qspi_controller q_ctrl (.\write_qspi_data_byte_idx_1__N_2021[0] (write_qspi_data_byte_idx_1__N_2021[0]), 
            .clk_c(clk_c), .qspi_data_ready(qspi_data_ready), .n6930(n6930), 
            .\writing_N_164[3] (\writing_N_164[3] ), .n27083(n27083), .\addr_in[24] (addr_in[24]), 
            .qspi_ram_b_select(qspi_ram_b_select), .spi_ram_b_select_N_2313(spi_ram_b_select_N_2313), 
            .clk_c_enable_341(clk_c_enable_341), .qspi_data_out_3__N_5({Open_2, 
            Open_3, Open_4, \qspi_data_out_3__N_5[0] }), .qspi_ram_a_select(qspi_ram_a_select), 
            .spi_ram_a_select_N_2309(spi_ram_a_select_N_2309), .is_writing(is_writing), 
            .ram_b_block_N_2303(ram_b_block_N_2303), .n24802(n24802), .qspi_data_in({qspi_data_in}), 
            .rst_reg_n(rst_reg_n), .\fsm_state[0] (\fsm_state[0] ), .n27082(n27082), 
            .n27299(n27299), .n23276(n23276), .spi_clk_pos(spi_clk_pos), 
            .clk_c_enable_358(clk_c_enable_358), .n27090(n27090), .\addr_in[14] (addr_in[14]), 
            .clk_c_enable_369(clk_c_enable_369), .n23252(n23252), .n9624(n9624), 
            .n27100(n27100), .\instr_data[8] (instr_data[8]), .last_ram_b_sel(last_ram_b_sel), 
            .clk_N_45(clk_N_45), .\addr_in[13] (addr_in[13]), .\addr_in[12] (addr_in[12]), 
            .\addr_in[11] (addr_in[11]), .\addr_in[15] (addr_in[15]), .\addr_in[9] (addr_in[9]), 
            .\addr_in[8] (addr_in[8]), .\addr_in[7] (addr_in[7]), .\addr_in[6] (addr_in[6]), 
            .\addr_in[10] (addr_in[10]), .\qspi_data_out_3__N_5[2] (\qspi_data_out_3__N_5[2] ), 
            .\addr_in[4] (addr_in[4]), .\instr_data[15] (instr_data[15]), 
            .\addr_in[5] (addr_in[5]), .clk_c_enable_392(clk_c_enable_392), 
            .\addr_23__N_2188[0] (addr_23__N_2188[0]), .n27081(n27081), 
            .n9702(n9702), .\addr_in[3] (addr_in[3]), .\addr_in[2] (addr_in[2]), 
            .\addr_in[1] (addr_in[1]), .\addr_in[16] (addr_in[16]), .\addr_in[17] (addr_in[17]), 
            .\addr_in[18] (addr_in[18]), .\addr_in[19] (addr_in[19]), .\addr_in[20] (addr_in[20]), 
            .\addr_in[21] (addr_in[21]), .n27105(n27105), .n27310(n27310), 
            .n1055(n1055), .clk_c_enable_79(clk_c_enable_79), .\addr_in[22] (addr_in[22]), 
            .n4319(n4319), .\instr_data[13] (instr_data[13]), .debug_stop_txn_N_2119(debug_stop_txn_N_2119), 
            .qspi_write_done(qspi_write_done), .n6942(n6942), .n27087(n27087), 
            .\instr_data[14] (instr_data[14]), .n4307(n4307), .\qspi_data_oe[3] (\qspi_data_oe[3] ), 
            .clk_c_enable_346(clk_c_enable_346), .ram_a_block_N_2299(ram_a_block_N_2299), 
            .n27080(n27080), .debug_stall_txn(debug_stall_txn), .data_stall(data_stall), 
            .\read_cycles_count[1] (read_cycles_count[1]), .n26130(n26130), 
            .n24688(n24688), .\qspi_data_out_3__N_5[3] (\qspi_data_out_3__N_5[3] ), 
            .\addr[20] (\addr[20]_adj_13 ), .\addr[22] (\addr[22]_adj_14 ), 
            .\instr_data[9] (instr_data[9]), .\instr_data[10] (instr_data[10]), 
            .\instr_data[11] (instr_data[11]), .\instr_data[12] (instr_data[12]), 
            .n482(n482), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .qspi_clk_N_56(qspi_clk_N_56), .start_instr(start_instr), .\addr[24] (\addr[24] ), 
            .instr_active(instr_active), .qspi_data_byte_idx({qspi_data_byte_idx}), 
            .n9(n9), .data_txn_len({data_txn_len_c[1], data_txn_len[0]}), 
            .n27272(n27272), .n27360(n27360), .n45(n45), .n27301(n27301), 
            .n27344(n27344), .n27357(n27357), .\addr[27] (\addr[27] ), 
            .n27265(n27265), .stop_txn_now_N_2363(stop_txn_now_N_2363), 
            .next_bit(next_bit), .n27210(n27210), .uart_txd_N_2596(uart_txd_N_2596), 
            .clk_c_enable_426(clk_c_enable_426), .n27271(n27271), .n27273(n27273), 
            .n8804(n8804), .n24376(n24376), .n22303(n22303), .n44(n44), 
            .clk_c_enable_273(clk_c_enable_273), .instr_active_N_2106(instr_active_N_2106), 
            .n805(n805), .clk_c_enable_420(clk_c_enable_420), .n27093(n27093), 
            .n22344(n22344), .qspi_data_byte_idx_1__N_2025(qspi_data_byte_idx_1__N_2025), 
            .n27345(n27345), .n27298(n27298), .n22180(n22180), .n27365(n27365), 
            .n22097(n22097), .n4309(n4309), .n24709(n24709), .n24700(n24700), 
            .n24703(n24703), .n24706(n24706), .n28559(n28559), .\data_to_write[26] (data_to_write[26]), 
            .n27325(n27325), .\instr_data_7__N_1969[26] (instr_data_7__N_1969[26]), 
            .\data_to_write[25] (data_to_write[25]), .\instr_data_7__N_1969[25] (instr_data_7__N_1969[25]), 
            .n9653(n9653), .n26711(n26711), .n5508(n5508), .n24704(n24704), 
            .n24707(n24707), .n5505(n5505), .n5909(n5909), .n22992(n22992), 
            .n24701(n24701), .n24710(n24710), .n26951(n26951), .n24691(n24691), 
            .n26945(n26945), .n24694(n24694), .n26939(n26939), .n24697(n24697)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(112[21] 136[6])
    
endmodule
//
// Verilog Description of module qspi_controller
//

module qspi_controller (\write_qspi_data_byte_idx_1__N_2021[0] , clk_c, 
            qspi_data_ready, n6930, \writing_N_164[3] , n27083, \addr_in[24] , 
            qspi_ram_b_select, spi_ram_b_select_N_2313, clk_c_enable_341, 
            qspi_data_out_3__N_5, qspi_ram_a_select, spi_ram_a_select_N_2309, 
            is_writing, ram_b_block_N_2303, n24802, qspi_data_in, rst_reg_n, 
            \fsm_state[0] , n27082, n27299, n23276, spi_clk_pos, clk_c_enable_358, 
            n27090, \addr_in[14] , clk_c_enable_369, n23252, n9624, 
            n27100, \instr_data[8] , last_ram_b_sel, clk_N_45, \addr_in[13] , 
            \addr_in[12] , \addr_in[11] , \addr_in[15] , \addr_in[9] , 
            \addr_in[8] , \addr_in[7] , \addr_in[6] , \addr_in[10] , 
            \qspi_data_out_3__N_5[2] , \addr_in[4] , \instr_data[15] , 
            \addr_in[5] , clk_c_enable_392, \addr_23__N_2188[0] , n27081, 
            n9702, \addr_in[3] , \addr_in[2] , \addr_in[1] , \addr_in[16] , 
            \addr_in[17] , \addr_in[18] , \addr_in[19] , \addr_in[20] , 
            \addr_in[21] , n27105, n27310, n1055, clk_c_enable_79, 
            \addr_in[22] , n4319, \instr_data[13] , debug_stop_txn_N_2119, 
            qspi_write_done, n6942, n27087, \instr_data[14] , n4307, 
            \qspi_data_oe[3] , clk_c_enable_346, ram_a_block_N_2299, n27080, 
            debug_stall_txn, data_stall, \read_cycles_count[1] , n26130, 
            n24688, \qspi_data_out_3__N_5[3] , \addr[20] , \addr[22] , 
            \instr_data[9] , \instr_data[10] , \instr_data[11] , \instr_data[12] , 
            n482, spi_clk_pos_derived_59, qspi_clk_N_56, start_instr, 
            \addr[24] , instr_active, qspi_data_byte_idx, n9, data_txn_len, 
            n27272, n27360, n45, n27301, n27344, n27357, \addr[27] , 
            n27265, stop_txn_now_N_2363, next_bit, n27210, uart_txd_N_2596, 
            clk_c_enable_426, n27271, n27273, n8804, n24376, n22303, 
            n44, clk_c_enable_273, instr_active_N_2106, n805, clk_c_enable_420, 
            n27093, n22344, qspi_data_byte_idx_1__N_2025, n27345, n27298, 
            n22180, n27365, n22097, n4309, n24709, n24700, n24703, 
            n24706, n28559, \data_to_write[26] , n27325, \instr_data_7__N_1969[26] , 
            \data_to_write[25] , \instr_data_7__N_1969[25] , n9653, n26711, 
            n5508, n24704, n24707, n5505, n5909, n22992, n24701, 
            n24710, n26951, n24691, n26945, n24694, n26939, n24697) /* synthesis syn_module_defined=1 */ ;
    output \write_qspi_data_byte_idx_1__N_2021[0] ;
    input clk_c;
    output qspi_data_ready;
    output n6930;
    output \writing_N_164[3] ;
    output n27083;
    input \addr_in[24] ;
    output qspi_ram_b_select;
    input spi_ram_b_select_N_2313;
    output clk_c_enable_341;
    input [3:0]qspi_data_out_3__N_5;
    output qspi_ram_a_select;
    input spi_ram_a_select_N_2309;
    output is_writing;
    input ram_b_block_N_2303;
    input n24802;
    input [3:0]qspi_data_in;
    input rst_reg_n;
    output \fsm_state[0] ;
    input n27082;
    output n27299;
    output n23276;
    output spi_clk_pos;
    input clk_c_enable_358;
    input n27090;
    input \addr_in[14] ;
    input clk_c_enable_369;
    output n23252;
    input n9624;
    input n27100;
    output \instr_data[8] ;
    output last_ram_b_sel;
    input clk_N_45;
    input \addr_in[13] ;
    input \addr_in[12] ;
    input \addr_in[11] ;
    input \addr_in[15] ;
    input \addr_in[9] ;
    input \addr_in[8] ;
    input \addr_in[7] ;
    input \addr_in[6] ;
    input \addr_in[10] ;
    input \qspi_data_out_3__N_5[2] ;
    input \addr_in[4] ;
    output \instr_data[15] ;
    input \addr_in[5] ;
    input clk_c_enable_392;
    input \addr_23__N_2188[0] ;
    input n27081;
    input n9702;
    input \addr_in[3] ;
    input \addr_in[2] ;
    input \addr_in[1] ;
    input \addr_in[16] ;
    input \addr_in[17] ;
    input \addr_in[18] ;
    input \addr_in[19] ;
    input \addr_in[20] ;
    input \addr_in[21] ;
    input n27105;
    output n27310;
    output n1055;
    output clk_c_enable_79;
    input \addr_in[22] ;
    output n4319;
    output \instr_data[13] ;
    input debug_stop_txn_N_2119;
    input qspi_write_done;
    output n6942;
    input n27087;
    output \instr_data[14] ;
    output n4307;
    output \qspi_data_oe[3] ;
    input clk_c_enable_346;
    output ram_a_block_N_2299;
    output n27080;
    input debug_stall_txn;
    input data_stall;
    output \read_cycles_count[1] ;
    input n26130;
    input n24688;
    input \qspi_data_out_3__N_5[3] ;
    output \addr[20] ;
    output \addr[22] ;
    output \instr_data[9] ;
    output \instr_data[10] ;
    output \instr_data[11] ;
    output \instr_data[12] ;
    output n482;
    output spi_clk_pos_derived_59;
    output qspi_clk_N_56;
    input start_instr;
    input \addr[24] ;
    input instr_active;
    input [1:0]qspi_data_byte_idx;
    output n9;
    input [1:0]data_txn_len;
    output n27272;
    output n27360;
    output n45;
    output n27301;
    input n27344;
    input n27357;
    input \addr[27] ;
    output n27265;
    input stop_txn_now_N_2363;
    input next_bit;
    input n27210;
    input uart_txd_N_2596;
    output clk_c_enable_426;
    input n27271;
    input n27273;
    output n8804;
    input n24376;
    input n22303;
    input n44;
    output clk_c_enable_273;
    output instr_active_N_2106;
    input n805;
    output clk_c_enable_420;
    input n27093;
    input n22344;
    output qspi_data_byte_idx_1__N_2025;
    input n27345;
    input n27298;
    output n22180;
    output n27365;
    output n22097;
    output n4309;
    input n24709;
    input n24700;
    input n24703;
    input n24706;
    input n28559;
    input \data_to_write[26] ;
    input n27325;
    output \instr_data_7__N_1969[26] ;
    input \data_to_write[25] ;
    output \instr_data_7__N_1969[25] ;
    output n9653;
    output n26711;
    output n5508;
    input n24704;
    input n24707;
    output n5505;
    input n5909;
    output n22992;
    input n24701;
    input n24710;
    input n26951;
    input n24691;
    input n26945;
    input n24694;
    input n26939;
    input n24697;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    
    wire n23033, data_req_N_2318, data_ready_N_2338, clk_c_enable_97;
    wire [1:0]delay_cycles_cfg;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(87[15:31])
    
    wire n27262;
    wire [3:0]spi_in_buffer;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(91[15:28])
    
    wire n26936, n26942;
    wire [1:0]read_cycles_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(105[15:32])
    
    wire clk_c_enable_349;
    wire [1:0]n396;
    wire [1:0]n4772;
    wire [2:0]nibbles_remaining;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(86[15:32])
    
    wire n27284, n8989;
    wire [2:0]n4136;
    
    wire stop_txn_reg, stop_txn_reg_N_2360;
    wire [2:0]fsm_state;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(82[15:24])
    
    wire n27411, n1102, n4, n9128, n27410, clk_c_enable_348, n27285, 
        n27221, n27239, clk_c_enable_419, n27312, n14701, n27283, 
        n14670, n27314, n6, clk_c_enable_355, n27225, n1094;
    wire [3:0]qspi_data_out_3__N_5_c;
    
    wire n26950;
    wire [23:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(84[31:35])
    wire [23:0]addr_23__N_2188;
    
    wire n1085, n27311, n27264, n27253, n1183, n5501, clk_c_enable_415;
    wire [7:0]data_out_7__N_2177;
    
    wire last_ram_a_sel, spi_clk_neg, n27313, spi_clk_use_neg, n26710, 
        n27412, n1087, n5;
    wire [1:0]n333;
    
    wire n27359, debug_stop_txn, n23358;
    wire [3:0]n4305;
    
    wire n23078, n27282;
    wire [2:0]n329;
    
    wire n26131, n26128, n25112, n15202, n25016, n26129, n27286, 
        n26127, n27370, n1086, n27323, n27378;
    wire [2:0]n312;
    
    wire n27281, n27373;
    wire [1:0]n381;
    wire [1:0]n181;
    wire [2:0]n356;
    wire [0:0]n4760;
    
    wire n1072, n23284, n23394, n24382, n23376;
    wire [7:0]data_out_7__N_2273;
    
    wire n24484;
    wire [55:0]instr_data_15__N_1959;
    
    wire n22112, n26948, n26944, n26938, n10, n26952, n26949, 
        n26946, n26943, n26940, n26937;
    
    FD1S3IX data_req_230 (.D(data_req_N_2318), .CK(clk_c), .CD(n23033), 
            .Q(\write_qspi_data_byte_idx_1__N_2021[0] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam data_req_230.GSR = "DISABLED";
    FD1S3IX data_ready_224 (.D(data_ready_N_2338), .CK(clk_c), .CD(n6930), 
            .Q(qspi_data_ready)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam data_ready_224.GSR = "DISABLED";
    FD1P3JX spi_flash_select_227 (.D(\addr_in[24] ), .SP(clk_c_enable_97), 
            .PD(n27083), .CK(clk_c), .Q(\writing_N_164[3] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_flash_select_227.GSR = "DISABLED";
    FD1P3JX spi_ram_b_select_229 (.D(spi_ram_b_select_N_2313), .SP(clk_c_enable_97), 
            .PD(n27083), .CK(clk_c), .Q(qspi_ram_b_select)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_ram_b_select_229.GSR = "DISABLED";
    FD1P3AX delay_cycles_cfg_i0_i0 (.D(qspi_data_out_3__N_5[0]), .SP(clk_c_enable_341), 
            .CK(clk_c), .Q(delay_cycles_cfg[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(112[12] 117[8])
    defparam delay_cycles_cfg_i0_i0.GSR = "DISABLED";
    FD1P3JX spi_ram_a_select_228 (.D(spi_ram_a_select_N_2309), .SP(clk_c_enable_97), 
            .PD(n27083), .CK(clk_c), .Q(qspi_ram_a_select)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_ram_a_select_228.GSR = "DISABLED";
    FD1P3IX is_writing_222 (.D(n24802), .SP(ram_b_block_N_2303), .CD(n27083), 
            .CK(clk_c), .Q(is_writing)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam is_writing_222.GSR = "DISABLED";
    LUT4 n9_bdd_4_lut_24252 (.A(n27262), .B(qspi_data_in[3]), .C(spi_in_buffer[3]), 
         .D(rst_reg_n), .Z(n26936)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam n9_bdd_4_lut_24252.init = 16'he4a0;
    LUT4 n9_bdd_4_lut_24327 (.A(n27262), .B(qspi_data_in[2]), .C(spi_in_buffer[2]), 
         .D(rst_reg_n), .Z(n26942)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam n9_bdd_4_lut_24327.init = 16'he4a0;
    FD1P3IX read_cycles_count__i0 (.D(n396[0]), .SP(clk_c_enable_349), .CD(n27083), 
            .CK(clk_c), .Q(read_cycles_count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam read_cycles_count__i0.GSR = "DISABLED";
    LUT4 mux_2616_i2_4_lut (.A(n4772[1]), .B(nibbles_remaining[1]), .C(n27284), 
         .D(n8989), .Z(n4136[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_2616_i2_4_lut.init = 16'hcac0;
    FD1S3IX stop_txn_reg_218 (.D(stop_txn_reg_N_2360), .CK(clk_c), .CD(clk_c_enable_341), 
            .Q(stop_txn_reg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(98[12] 103[8])
    defparam stop_txn_reg_218.GSR = "DISABLED";
    LUT4 mux_113_i3_4_lut_then_4_lut (.A(n27284), .B(fsm_state[2]), .C(fsm_state[1]), 
         .D(\fsm_state[0] ), .Z(n27411)) /* synthesis lut_function=(A (B (C (D)))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_113_i3_4_lut_then_4_lut.init = 16'hd454;
    LUT4 mux_681_i3_4_lut (.A(n4136[2]), .B(\addr_in[24] ), .C(n1102), 
         .D(n4), .Z(n9128)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam mux_681_i3_4_lut.init = 16'h3a35;
    LUT4 mux_113_i3_4_lut_else_4_lut (.A(n27284), .B(fsm_state[2]), .C(fsm_state[1]), 
         .D(\fsm_state[0] ), .Z(n27410)) /* synthesis lut_function=(A (B (C (D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_113_i3_4_lut_else_4_lut.init = 16'hd444;
    LUT4 i1_3_lut_4_lut (.A(n27082), .B(ram_b_block_N_2303), .C(n27299), 
         .D(n27083), .Z(clk_c_enable_348)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i1_3_lut_4_lut.init = 16'hfff8;
    LUT4 i23642_2_lut_4_lut_4_lut (.A(n27285), .B(is_writing), .C(n27221), 
         .D(n27239), .Z(clk_c_enable_419)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (C (D))))) */ ;
    defparam i23642_2_lut_4_lut_4_lut.init = 16'h1ddd;
    LUT4 i1_3_lut_4_lut_adj_450 (.A(\fsm_state[0] ), .B(n27312), .C(n27284), 
         .D(n14701), .Z(n23276)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_adj_450.init = 16'h0070;
    LUT4 i12368_3_lut_4_lut (.A(\fsm_state[0] ), .B(n27312), .C(is_writing), 
         .D(n27283), .Z(n14670)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;
    defparam i12368_3_lut_4_lut.init = 16'h7770;
    LUT4 i789_2_lut_rep_614_3_lut_4_lut (.A(fsm_state[2]), .B(n27314), .C(spi_clk_pos), 
         .D(n27284), .Z(n27239)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A ((D)+!C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i789_2_lut_rep_614_3_lut_4_lut.init = 16'hdf0f;
    LUT4 i1_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n27314), .C(spi_clk_pos), 
         .D(n27284), .Z(n6)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h20f0;
    FD1P3AX spi_in_buffer_i0_i0 (.D(qspi_data_out_3__N_5[0]), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(spi_in_buffer[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_451 (.A(fsm_state[2]), .B(n27314), .C(is_writing), 
         .D(n27284), .Z(data_req_N_2318)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_3_lut_4_lut_adj_451.init = 16'h0020;
    LUT4 i1_2_lut_rep_600_3_lut_4_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n27314), 
         .C(spi_clk_pos), .D(n27284), .Z(n27225)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_600_3_lut_4_lut_3_lut_4_lut.init = 16'h2000;
    FD1P3IX nibbles_remaining__i0 (.D(n1094), .SP(clk_c_enable_358), .CD(n27083), 
            .CK(clk_c), .Q(nibbles_remaining[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i0.GSR = "DISABLED";
    LUT4 n5072_bdd_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n27314), .C(qspi_data_out_3__N_5_c[1]), 
         .D(n27284), .Z(n26950)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam n5072_bdd_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 addr_23__I_0_i15_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[14] ), 
         .D(addr[10]), .Z(addr_23__N_2188[14])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i15_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX fsm_state__i0 (.D(n1085), .SP(clk_c_enable_369), .CD(n27083), 
            .CK(clk_c), .Q(\fsm_state[0] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i0.GSR = "DISABLED";
    LUT4 i3149_2_lut_rep_639_3_lut_4_lut (.A(nibbles_remaining[0]), .B(n27311), 
         .C(n27314), .D(fsm_state[2]), .Z(n27264)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i3149_2_lut_rep_639_3_lut_4_lut.init = 16'h0e00;
    LUT4 i1_4_lut_4_lut (.A(n27284), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(\fsm_state[0] ), .Z(n23252)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(209[30] 211[24])
    defparam i1_4_lut_4_lut.init = 16'h0041;
    LUT4 i1_3_lut_4_lut_adj_452 (.A(nibbles_remaining[0]), .B(n27311), .C(n9624), 
         .D(n27253), .Z(n1183)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_3_lut_4_lut_adj_452.init = 16'hefff;
    LUT4 i2892_3_lut_4_lut (.A(n27082), .B(ram_b_block_N_2303), .C(n27299), 
         .D(n27100), .Z(n5501)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i2892_3_lut_4_lut.init = 16'h08f8;
    FD1P3AX data_i1 (.D(data_out_7__N_2177[0]), .SP(clk_c_enable_415), .CK(clk_c), 
            .Q(\instr_data[8] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i1.GSR = "DISABLED";
    FD1S3JX last_ram_a_sel_235 (.D(qspi_ram_a_select), .CK(clk_c), .PD(clk_c_enable_341), 
            .Q(last_ram_a_sel)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(272[12] 280[8])
    defparam last_ram_a_sel_235.GSR = "DISABLED";
    FD1S3JX last_ram_b_sel_236 (.D(qspi_ram_b_select), .CK(clk_c), .PD(clk_c_enable_341), 
            .Q(last_ram_b_sel)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(272[12] 280[8])
    defparam last_ram_b_sel_236.GSR = "DISABLED";
    FD1S3AX spi_clk_neg_237 (.D(spi_clk_pos), .CK(clk_N_45), .Q(spi_clk_neg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(286[12:54])
    defparam spi_clk_neg_237.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_637_4_lut (.A(fsm_state[2]), .B(\fsm_state[0] ), .C(n27313), 
         .D(fsm_state[1]), .Z(n27262)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_637_4_lut.init = 16'hfff7;
    LUT4 addr_23__I_0_i14_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[13] ), 
         .D(addr[9]), .Z(addr_23__N_2188[13])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i13_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[12] ), 
         .D(addr[8]), .Z(addr_23__N_2188[12])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i12_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[11] ), 
         .D(addr[7]), .Z(addr_23__N_2188[11])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i16_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[15] ), 
         .D(addr[11]), .Z(addr_23__N_2188[15])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i16_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i10_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[9] ), 
         .D(addr[5]), .Z(addr_23__N_2188[9])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i9_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[8] ), 
         .D(addr[4]), .Z(addr_23__N_2188[8])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i9_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i8_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[7] ), 
         .D(addr[3]), .Z(addr_23__N_2188[7])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i7_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[6] ), 
         .D(addr[2]), .Z(addr_23__N_2188[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i11_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[10] ), 
         .D(addr[6]), .Z(addr_23__N_2188[10])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i11_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX spi_clk_use_neg_220 (.D(\qspi_data_out_3__N_5[2] ), .SP(clk_c_enable_341), 
            .CK(clk_c), .Q(spi_clk_use_neg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(112[12] 117[8])
    defparam spi_clk_use_neg_220.GSR = "DISABLED";
    LUT4 addr_23__I_0_i5_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[4] ), 
         .D(addr[0]), .Z(addr_23__N_2188[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__bdd_4_lut (.A(\instr_data[15] ), .B(fsm_state[2]), .C(is_writing), 
         .D(nibbles_remaining[0]), .Z(n26710)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B (C)+!B (C+(D)))) */ ;
    defparam addr_23__bdd_4_lut.init = 16'h8c8f;
    LUT4 addr_23__I_0_i6_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[5] ), 
         .D(addr[1]), .Z(addr_23__N_2188[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i6_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX addr_i0 (.D(\addr_23__N_2188[0] ), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i0.GSR = "DISABLED";
    LUT4 i12683_3_lut_4_lut (.A(n27299), .B(n27081), .C(n14701), .D(n27412), 
         .Z(n1087)) /* synthesis lut_function=(A (C+(D))+!A !(B+!(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i12683_3_lut_4_lut.init = 16'hbbb0;
    FD1P3IX addr_i3 (.D(\addr_in[3] ), .SP(clk_c_enable_392), .CD(n9702), 
            .CK(clk_c), .Q(addr[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i3.GSR = "DISABLED";
    FD1P3IX addr_i2 (.D(\addr_in[2] ), .SP(clk_c_enable_392), .CD(n9702), 
            .CK(clk_c), .Q(addr[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i2.GSR = "DISABLED";
    FD1P3IX addr_i1 (.D(\addr_in[1] ), .SP(clk_c_enable_392), .CD(n9702), 
            .CK(clk_c), .Q(addr[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i1.GSR = "DISABLED";
    LUT4 addr_23__I_0_i17_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[16] ), 
         .D(addr[12]), .Z(addr_23__N_2188[16])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i18_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[17] ), 
         .D(addr[13]), .Z(addr_23__N_2188[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i19_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[18] ), 
         .D(addr[14]), .Z(addr_23__N_2188[18])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i20_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[19] ), 
         .D(addr[15]), .Z(addr_23__N_2188[19])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i21_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[20] ), 
         .D(addr[16]), .Z(addr_23__N_2188[20])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(\fsm_state[0] ), 
         .Z(n5)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(169[58:88])
    defparam i1_3_lut.init = 16'hf7f7;
    LUT4 addr_23__I_0_i22_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[21] ), 
         .D(addr[17]), .Z(addr_23__N_2188[21])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i22_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_106_i1_4_lut (.A(delay_cycles_cfg[0]), .B(n27105), .C(n27310), 
         .D(n1055), .Z(n333[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(178[38] 204[32])
    defparam mux_106_i1_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut_4_lut_adj_453 (.A(fsm_state[2]), .B(n27359), .C(debug_stop_txn), 
         .D(rst_reg_n), .Z(clk_c_enable_79)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_3_lut_4_lut_adj_453.init = 16'hf1ff;
    LUT4 addr_23__I_0_i23_3_lut_4_lut (.A(n27299), .B(n27090), .C(\addr_in[22] ), 
         .D(addr[18]), .Z(addr_23__N_2188[22])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i23_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut_adj_454 (.A(fsm_state[2]), .B(n27359), .C(stop_txn_reg), 
         .D(spi_clk_pos), .Z(n23358)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_3_lut_4_lut_adj_454.init = 16'hfff1;
    FD1P3AX delay_cycles_cfg_i0_i1 (.D(qspi_data_out_3__N_5_c[1]), .SP(clk_c_enable_341), 
            .CK(clk_c), .Q(delay_cycles_cfg[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(112[12] 117[8])
    defparam delay_cycles_cfg_i0_i1.GSR = "DISABLED";
    LUT4 mux_2648_i2_3_lut (.A(addr[21]), .B(n4305[1]), .C(\fsm_state[0] ), 
         .Z(n4319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_2648_i2_3_lut.init = 16'hcaca;
    LUT4 mux_2641_i2_4_lut (.A(nibbles_remaining[0]), .B(\instr_data[13] ), 
         .C(fsm_state[2]), .D(is_writing), .Z(n4305[1])) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B+!(C (D)))) */ ;
    defparam mux_2641_i2_4_lut.init = 16'hc5f5;
    LUT4 i12178_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n27359), .C(debug_stop_txn_N_2119), 
         .D(qspi_write_done), .Z(debug_stop_txn)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i12178_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i23571_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n27359), .C(rst_reg_n), 
         .D(qspi_write_done), .Z(n6942)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i23571_2_lut_3_lut_4_lut.init = 16'h0f1f;
    LUT4 addr_23__I_0_i24_3_lut_4_lut (.A(n27299), .B(n27090), .C(n27087), 
         .D(addr[19]), .Z(addr_23__N_2188[23])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i24_3_lut_4_lut.init = 16'hfb40;
    LUT4 i12589_3_lut (.A(\instr_data[14] ), .B(fsm_state[2]), .C(is_writing), 
         .Z(n4307)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i12589_3_lut.init = 16'h8c8c;
    FD1P3IX spi_data_oe__i3 (.D(n1102), .SP(clk_c_enable_346), .CD(n27083), 
            .CK(clk_c), .Q(\qspi_data_oe[3] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_data_oe__i3.GSR = "DISABLED";
    FD1P3AX spi_clk_pos_225 (.D(n23078), .SP(clk_c_enable_348), .CK(clk_c), 
            .Q(spi_clk_pos)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_clk_pos_225.GSR = "DISABLED";
    LUT4 i674_rep_455_3_lut_4_lut (.A(ram_a_block_N_2299), .B(n27090), .C(n27299), 
         .D(ram_b_block_N_2303), .Z(n27080)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i674_rep_455_3_lut_4_lut.init = 16'h0800;
    LUT4 mux_105_i1_4_lut (.A(debug_stall_txn), .B(n27282), .C(n27284), 
         .D(data_stall), .Z(n329[0])) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(178[38] 204[32])
    defparam mux_105_i1_4_lut.init = 16'hc0c5;
    L6MUX21 i23776 (.D0(n26131), .D1(n26128), .SD(n25112), .Z(data_out_7__N_2177[0]));
    FD1P3IX read_cycles_count__i1 (.D(n396[1]), .SP(clk_c_enable_349), .CD(n27083), 
            .CK(clk_c), .Q(\read_cycles_count[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam read_cycles_count__i1.GSR = "DISABLED";
    LUT4 i23616_3_lut_4_lut (.A(nibbles_remaining[0]), .B(n27311), .C(n1102), 
         .D(n4136[1]), .Z(n15202)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+(D))+!B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam i23616_3_lut_4_lut.init = 16'h0b04;
    LUT4 i1_2_lut_rep_685 (.A(fsm_state[2]), .B(\fsm_state[0] ), .Z(n27310)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_685.init = 16'h8888;
    LUT4 i23684_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(\fsm_state[0] ), 
         .C(n27311), .D(nibbles_remaining[0]), .Z(n25016)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i23684_2_lut_3_lut_4_lut.init = 16'hfff8;
    LUT4 equal_117_i4_2_lut_rep_686 (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .Z(n27311)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam equal_117_i4_2_lut_rep_686.init = 16'heeee;
    LUT4 equal_117_i5_2_lut_rep_659_3_lut (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .C(nibbles_remaining[0]), .Z(n27284)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam equal_117_i5_2_lut_rep_659_3_lut.init = 16'hfefe;
    LUT4 i3811_2_lut_3_lut_4_lut (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .C(n4136[1]), .D(nibbles_remaining[0]), .Z(n4)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i3811_2_lut_3_lut_4_lut.init = 16'hfff1;
    PFUMX i23774 (.BLUT(n26130), .ALUT(n26129), .C0(n27221), .Z(n26131));
    LUT4 mux_2616_i3_3_lut_4_lut_4_lut (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .C(n27286), .D(nibbles_remaining[0]), .Z(n4136[2])) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam mux_2616_i3_3_lut_4_lut_4_lut.init = 16'hcccd;
    LUT4 i1_2_lut_rep_687 (.A(fsm_state[2]), .B(fsm_state[1]), .Z(n27312)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_687.init = 16'h8888;
    LUT4 i1_2_lut_rep_657_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(\fsm_state[0] ), 
         .Z(n27282)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_657_3_lut.init = 16'h8080;
    LUT4 i12195_2_lut_rep_688 (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .Z(n27313)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12195_2_lut_rep_688.init = 16'heeee;
    LUT4 i1_3_lut_rep_660_4_lut (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .C(\fsm_state[0] ), .D(fsm_state[2]), .Z(n27285)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_3_lut_rep_660_4_lut.init = 16'hefff;
    LUT4 i27_3_lut_4_lut (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .C(n14670), .D(spi_clk_pos), .Z(n27253)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam i27_3_lut_4_lut.init = 16'hf101;
    PFUMX i23771 (.BLUT(n24688), .ALUT(n26127), .C0(n27370), .Z(n26128));
    LUT4 i1_2_lut_rep_689 (.A(fsm_state[1]), .B(\fsm_state[0] ), .Z(n27314)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_689.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_658_3_lut (.A(fsm_state[1]), .B(\fsm_state[0] ), .C(fsm_state[2]), 
         .Z(n27283)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_658_3_lut.init = 16'hbfbf;
    FD1P3AX spi_in_buffer_i0_i1 (.D(qspi_data_out_3__N_5_c[1]), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(spi_in_buffer[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i1.GSR = "DISABLED";
    FD1P3AX spi_in_buffer_i0_i2 (.D(\qspi_data_out_3__N_5[2] ), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(spi_in_buffer[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX spi_in_buffer_i0_i3 (.D(\qspi_data_out_3__N_5[3] ), .SP(clk_c_enable_355), 
            .CK(clk_c), .Q(spi_in_buffer[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i3.GSR = "DISABLED";
    FD1P3IX nibbles_remaining__i1 (.D(n15202), .SP(clk_c_enable_358), .CD(n27083), 
            .CK(clk_c), .Q(nibbles_remaining[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_661_3_lut (.A(fsm_state[1]), .B(\fsm_state[0] ), .C(fsm_state[2]), 
         .Z(n27286)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_661_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_3_lut_3_lut (.A(fsm_state[1]), .B(\fsm_state[0] ), 
         .C(fsm_state[2]), .Z(n8989)) /* synthesis lut_function=(!(A (B (C))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_3_lut_3_lut_3_lut.init = 16'h3b3b;
    FD1P3IX nibbles_remaining__i2 (.D(n9128), .SP(clk_c_enable_358), .CD(n27083), 
            .CK(clk_c), .Q(nibbles_remaining[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i2.GSR = "DISABLED";
    FD1P3IX fsm_state__i1 (.D(n1086), .SP(clk_c_enable_369), .CD(n27083), 
            .CK(clk_c), .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i1.GSR = "DISABLED";
    FD1P3IX fsm_state__i2 (.D(n1087), .SP(clk_c_enable_369), .CD(n27083), 
            .CK(clk_c), .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1P3AX addr_i4 (.D(addr_23__N_2188[4]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i4.GSR = "DISABLED";
    FD1P3AX addr_i5 (.D(addr_23__N_2188[5]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i5.GSR = "DISABLED";
    FD1P3AX addr_i6 (.D(addr_23__N_2188[6]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i6.GSR = "DISABLED";
    FD1P3AX addr_i7 (.D(addr_23__N_2188[7]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i7.GSR = "DISABLED";
    FD1P3AX addr_i8 (.D(addr_23__N_2188[8]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i8.GSR = "DISABLED";
    FD1P3AX addr_i9 (.D(addr_23__N_2188[9]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i9.GSR = "DISABLED";
    FD1P3AX addr_i10 (.D(addr_23__N_2188[10]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i10.GSR = "DISABLED";
    FD1P3AX addr_i11 (.D(addr_23__N_2188[11]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i11.GSR = "DISABLED";
    FD1P3AX addr_i12 (.D(addr_23__N_2188[12]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i12.GSR = "DISABLED";
    FD1P3AX addr_i13 (.D(addr_23__N_2188[13]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i13.GSR = "DISABLED";
    FD1P3AX addr_i14 (.D(addr_23__N_2188[14]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i14.GSR = "DISABLED";
    FD1P3AX addr_i15 (.D(addr_23__N_2188[15]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i15.GSR = "DISABLED";
    FD1P3AX addr_i16 (.D(addr_23__N_2188[16]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i16.GSR = "DISABLED";
    FD1P3AX addr_i17 (.D(addr_23__N_2188[17]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i17.GSR = "DISABLED";
    FD1P3AX addr_i18 (.D(addr_23__N_2188[18]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i18.GSR = "DISABLED";
    FD1P3AX addr_i19 (.D(addr_23__N_2188[19]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i19.GSR = "DISABLED";
    FD1P3AX addr_i20 (.D(addr_23__N_2188[20]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\addr[20] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i20.GSR = "DISABLED";
    FD1P3AX addr_i21 (.D(addr_23__N_2188[21]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i21.GSR = "DISABLED";
    FD1P3AX addr_i22 (.D(addr_23__N_2188[22]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\addr[22] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i22.GSR = "DISABLED";
    FD1P3AX addr_i23 (.D(addr_23__N_2188[23]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(addr[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i23.GSR = "DISABLED";
    FD1P3AX data_i2 (.D(data_out_7__N_2177[1]), .SP(clk_c_enable_415), .CK(clk_c), 
            .Q(\instr_data[9] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i2.GSR = "DISABLED";
    FD1P3AX data_i3 (.D(data_out_7__N_2177[2]), .SP(clk_c_enable_415), .CK(clk_c), 
            .Q(\instr_data[10] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i3.GSR = "DISABLED";
    FD1P3AX data_i4 (.D(data_out_7__N_2177[3]), .SP(clk_c_enable_415), .CK(clk_c), 
            .Q(\instr_data[11] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i4.GSR = "DISABLED";
    FD1P3AX data_i5 (.D(data_out_7__N_2177[4]), .SP(clk_c_enable_419), .CK(clk_c), 
            .Q(\instr_data[12] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i5.GSR = "DISABLED";
    FD1P3AX data_i6 (.D(data_out_7__N_2177[5]), .SP(clk_c_enable_419), .CK(clk_c), 
            .Q(\instr_data[13] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i6.GSR = "DISABLED";
    FD1P3AX data_i7 (.D(data_out_7__N_2177[6]), .SP(clk_c_enable_419), .CK(clk_c), 
            .Q(\instr_data[14] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i7.GSR = "DISABLED";
    FD1P3AX data_i8 (.D(data_out_7__N_2177[7]), .SP(clk_c_enable_419), .CK(clk_c), 
            .Q(\instr_data[15] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i8.GSR = "DISABLED";
    LUT4 mux_2864_i2_3_lut_4_lut_3_lut_4_lut (.A(\writing_N_164[3] ), .B(is_writing), 
         .C(n27323), .D(\fsm_state[0] ), .Z(n4772[1])) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(187[46] 194[40])
    defparam mux_2864_i2_3_lut_4_lut_3_lut_4_lut.init = 16'h0f02;
    LUT4 fsm_state_2__I_0_240_i4_2_lut_rep_698 (.A(fsm_state[1]), .B(fsm_state[2]), 
         .Z(n27323)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(265[13:23])
    defparam fsm_state_2__I_0_240_i4_2_lut_rep_698.init = 16'hdddd;
    LUT4 i12669_3_lut_4_lut_4_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(n27378), .D(\fsm_state[0] ), .Z(n312[1])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(265[13:23])
    defparam i12669_3_lut_4_lut_4_lut_4_lut.init = 16'h558a;
    LUT4 fsm_state_2__I_0_239_i5_2_lut_rep_656_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(\fsm_state[0] ), .Z(n27281)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(265[13:23])
    defparam fsm_state_2__I_0_239_i5_2_lut_rep_656_3_lut.init = 16'hfdfd;
    LUT4 mux_114_i2_4_lut (.A(delay_cycles_cfg[1]), .B(n27373), .C(n1183), 
         .D(n9624), .Z(n381[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_114_i2_4_lut.init = 16'hcac0;
    LUT4 i171_2_lut_3_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(spi_clk_pos), 
         .D(\fsm_state[0] ), .Z(n482)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(265[13:23])
    defparam i171_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 spi_clk_pos_I_0_256_3_lut_rep_703 (.A(spi_clk_pos), .B(spi_clk_neg), 
         .C(spi_clk_use_neg), .Z(spi_clk_pos_derived_59)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(287[26:69])
    defparam spi_clk_pos_I_0_256_3_lut_rep_703.init = 16'hcaca;
    LUT4 qspi_clk_I_0_1_lut_3_lut (.A(spi_clk_pos), .B(spi_clk_neg), .C(spi_clk_use_neg), 
         .Z(qspi_clk_N_56)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(287[26:69])
    defparam qspi_clk_I_0_1_lut_3_lut.init = 16'h3535;
    PFUMX mux_129_i2 (.BLUT(n181[1]), .ALUT(n381[1]), .C0(n5), .Z(n396[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 n9_bdd_4_lut_23901 (.A(n27262), .B(qspi_data_in[0]), .C(spi_in_buffer[0]), 
         .D(rst_reg_n), .Z(n26127)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam n9_bdd_4_lut_23901.init = 16'he4a0;
    PFUMX mux_129_i1 (.BLUT(n181[0]), .ALUT(n381[0]), .C0(n5), .Z(n396[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX mux_662_i2 (.BLUT(n356[1]), .ALUT(n4760[0]), .C0(n14701), .Z(n1072));
    LUT4 i1_4_lut (.A(ram_a_block_N_2299), .B(ram_b_block_N_2303), .C(n27090), 
         .D(n27299), .Z(n1102)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i1_4_lut.init = 16'h0080;
    LUT4 i1_4_lut_adj_455 (.A(start_instr), .B(n27087), .C(\addr[24] ), 
         .D(n23284), .Z(ram_a_block_N_2299)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(109[49:72])
    defparam i1_4_lut_adj_455.init = 16'hffef;
    LUT4 i1_2_lut (.A(instr_active), .B(last_ram_a_sel), .Z(n23284)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(109[49:72])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i23657_4_lut (.A(qspi_data_byte_idx[0]), .B(n23394), .C(start_instr), 
         .D(instr_active), .Z(n9)) /* synthesis lut_function=(!(A+!((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[10:18])
    defparam i23657_4_lut.init = 16'h5551;
    LUT4 i1_3_lut_adj_456 (.A(data_txn_len[0]), .B(data_txn_len[1]), .C(qspi_data_byte_idx[1]), 
         .Z(n23394)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C)))) */ ;
    defparam i1_3_lut_adj_456.init = 16'h4141;
    LUT4 i1_2_lut_rep_734 (.A(\fsm_state[0] ), .B(fsm_state[1]), .Z(n27359)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_734.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(\fsm_state[0] ), .B(fsm_state[1]), 
         .C(n27311), .D(fsm_state[2]), .Z(n24382)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h0e03;
    LUT4 i1_2_lut_rep_674_3_lut (.A(\fsm_state[0] ), .B(fsm_state[1]), .C(fsm_state[2]), 
         .Z(n27299)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_674_3_lut.init = 16'hfefe;
    LUT4 qspi_busy_I_0_2_lut_rep_647_3_lut_4_lut (.A(\fsm_state[0] ), .B(fsm_state[1]), 
         .C(qspi_write_done), .D(fsm_state[2]), .Z(n27272)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam qspi_busy_I_0_2_lut_rep_647_3_lut_4_lut.init = 16'hfffe;
    PFUMX mux_113_i1 (.BLUT(n312[0]), .ALUT(n329[0]), .C0(n25016), .Z(n356[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_2_lut_3_lut (.A(\fsm_state[0] ), .B(fsm_state[1]), 
         .C(fsm_state[2]), .Z(n1055)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_3_lut_4_lut_2_lut_3_lut.init = 16'h1010;
    LUT4 i39_2_lut_rep_735 (.A(data_txn_len[1]), .B(qspi_data_byte_idx[1]), 
         .Z(n27360)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(59[15:33])
    defparam i39_2_lut_rep_735.init = 16'h6666;
    LUT4 i11080_3_lut_4_lut_4_lut (.A(data_txn_len[1]), .B(qspi_data_byte_idx[1]), 
         .C(start_instr), .D(instr_active), .Z(n45)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(59[15:33])
    defparam i11080_3_lut_4_lut_4_lut.init = 16'hccc6;
    LUT4 i23439_3_lut_rep_676_4_lut (.A(data_txn_len[1]), .B(qspi_data_byte_idx[1]), 
         .C(data_txn_len[0]), .D(qspi_data_byte_idx[0]), .Z(n27301)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(59[15:33])
    defparam i23439_3_lut_rep_676_4_lut.init = 16'h9009;
    LUT4 i12673_4_lut_4_lut (.A(n27284), .B(n27310), .C(n27105), .D(n312[1]), 
         .Z(n356[1])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i12673_4_lut_4_lut.init = 16'h5140;
    LUT4 rst_n_I_0_1_lut_rep_739 (.A(rst_reg_n), .Z(clk_c_enable_341)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam rst_n_I_0_1_lut_rep_739.init = 16'h5555;
    LUT4 i1_3_lut_rep_640_4_lut_4_lut (.A(rst_reg_n), .B(n27344), .C(n27357), 
         .D(\addr[27] ), .Z(n27265)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_3_lut_rep_640_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_457 (.A(rst_reg_n), .B(n23376), .C(stop_txn_now_N_2363), 
         .D(n27253), .Z(n23033)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_457.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_458 (.A(rst_reg_n), .B(stop_txn_reg), .C(n27299), 
         .D(stop_txn_now_N_2363), .Z(clk_c_enable_349)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_458.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_459 (.A(rst_reg_n), .B(next_bit), .C(n27210), 
         .D(uart_txd_N_2596), .Z(clk_c_enable_426)) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_459.init = 16'hfdf5;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(n27271), .C(n27273), 
         .D(n27272), .Z(n8804)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hff7f;
    LUT4 i1_4_lut_4_lut_adj_460 (.A(rst_reg_n), .B(n24376), .C(n22303), 
         .D(n44), .Z(clk_c_enable_273)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_460.init = 16'h5d55;
    LUT4 rstn_N_2029_I_0_2_lut_2_lut (.A(rst_reg_n), .B(debug_stop_txn), 
         .Z(instr_active_N_2106)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam rstn_N_2029_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_2_lut (.A(rst_reg_n), .B(n805), .Z(clk_c_enable_420)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut_adj_461 (.A(rst_reg_n), .B(n27093), .C(n22344), 
         .D(n27272), .Z(qspi_data_byte_idx_1__N_2025)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_461.init = 16'h55df;
    LUT4 i1_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n27345), .C(n27344), 
         .D(n27298), .Z(n22180)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_2_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i12266_2_lut_2_lut (.A(rst_reg_n), .B(qspi_data_in[1]), .Z(qspi_data_out_3__N_5_c[1])) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i12266_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_rep_458_3_lut (.A(rst_reg_n), .B(stop_txn_reg), .C(stop_txn_now_N_2363), 
         .Z(n27083)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_3_lut_rep_458_3_lut.init = 16'hfdfd;
    LUT4 i1_4_lut_4_lut_adj_462 (.A(rst_reg_n), .B(stop_txn_reg), .C(stop_txn_now_N_2363), 
         .D(n27299), .Z(n6930)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_462.init = 16'hfdff;
    LUT4 i1_2_lut_4_lut_4_lut_adj_463 (.A(rst_reg_n), .B(n1102), .C(stop_txn_reg), 
         .D(stop_txn_now_N_2363), .Z(clk_c_enable_97)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_2_lut_4_lut_4_lut_adj_463.init = 16'hfffd;
    LUT4 i13_3_lut_rep_740 (.A(fsm_state[2]), .B(\fsm_state[0] ), .C(fsm_state[1]), 
         .Z(n27365)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam i13_3_lut_rep_740.init = 16'h1c1c;
    LUT4 i1_2_lut_4_lut (.A(fsm_state[2]), .B(\fsm_state[0] ), .C(fsm_state[1]), 
         .D(\qspi_data_oe[3] ), .Z(n22097)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C (D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h1c00;
    LUT4 mux_2641_i1_4_lut_4_lut (.A(nibbles_remaining[0]), .B(is_writing), 
         .C(fsm_state[2]), .D(\instr_data[12] ), .Z(n4309)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A ((C (D))+!B)) */ ;
    defparam mux_2641_i1_4_lut_4_lut.init = 16'hf131;
    LUT4 i1_3_lut_adj_464 (.A(debug_stop_txn), .B(stop_txn_now_N_2363), 
         .C(stop_txn_reg), .Z(stop_txn_reg_N_2360)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut_adj_464.init = 16'h0202;
    LUT4 is_writing_I_0_1_lut_rep_745 (.A(is_writing), .Z(n27370)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[52:63])
    defparam is_writing_I_0_1_lut_rep_745.init = 16'h5555;
    LUT4 i12361_2_lut_2_lut (.A(is_writing), .B(delay_cycles_cfg[1]), .Z(n4760[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[52:63])
    defparam i12361_2_lut_2_lut.init = 16'h4444;
    LUT4 mux_180_i8_3_lut_3_lut (.A(is_writing), .B(\instr_data[11] ), .C(n24709), 
         .Z(data_out_7__N_2273[7])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[52:63])
    defparam mux_180_i8_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i5_3_lut_3_lut (.A(is_writing), .B(\instr_data[8] ), .C(n24700), 
         .Z(data_out_7__N_2273[4])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[52:63])
    defparam mux_180_i5_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i6_3_lut_3_lut (.A(is_writing), .B(\instr_data[9] ), .C(n24703), 
         .Z(data_out_7__N_2273[5])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[52:63])
    defparam mux_180_i6_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i7_3_lut_3_lut (.A(is_writing), .B(\instr_data[10] ), .C(n24706), 
         .Z(data_out_7__N_2273[6])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[52:63])
    defparam mux_180_i7_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_114_i1_3_lut_3_lut (.A(read_cycles_count[0]), .B(n1183), .C(n333[0]), 
         .Z(n381[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam mux_114_i1_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_60_i1_4_lut_4_lut_4_lut_4_lut (.A(read_cycles_count[0]), .B(n27100), 
         .C(delay_cycles_cfg[0]), .D(is_writing), .Z(n181[0])) /* synthesis lut_function=(!(A (B+((D)+!C))+!A !(B+!((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam mux_60_i1_4_lut_4_lut_4_lut_4_lut.init = 16'h4474;
    LUT4 i1_2_lut_rep_748 (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .Z(n27373)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_748.init = 16'h8888;
    LUT4 i12667_2_lut_3_lut_4_lut_2_lut (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .Z(n181[1])) /* synthesis lut_function=(A (B)) */ ;
    defparam i12667_2_lut_3_lut_4_lut_2_lut.init = 16'h8888;
    LUT4 mux_674_i2_3_lut_4_lut (.A(\addr[24] ), .B(n28559), .C(n1102), 
         .D(n1072), .Z(n1086)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;
    defparam mux_674_i2_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i12424_2_lut_rep_753 (.A(\writing_N_164[3] ), .B(is_writing), .Z(n27378)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12424_2_lut_rep_753.init = 16'heeee;
    LUT4 mux_95_i1_3_lut_4_lut_4_lut_4_lut (.A(\writing_N_164[3] ), .B(is_writing), 
         .C(n27281), .D(\fsm_state[0] ), .Z(n312[0])) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A (B (C (D))+!B (D)))) */ ;
    defparam mux_95_i1_3_lut_4_lut_4_lut_4_lut.init = 16'h0cfd;
    LUT4 i11072_4_lut (.A(\data_to_write[26] ), .B(\instr_data[10] ), .C(qspi_data_ready), 
         .D(n27325), .Z(\instr_data_7__N_1969[26] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i11072_4_lut.init = 16'hca0a;
    LUT4 i11074_4_lut (.A(\data_to_write[25] ), .B(\instr_data[9] ), .C(qspi_data_ready), 
         .D(n27325), .Z(\instr_data_7__N_1969[25] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i11074_4_lut.init = 16'hca0a;
    LUT4 i7306_1_lut (.A(\write_qspi_data_byte_idx_1__N_2021[0] ), .Z(n9653)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i7306_1_lut.init = 16'h5555;
    LUT4 addr_23__bdd_3_lut_24114 (.A(addr[23]), .B(n26710), .C(\fsm_state[0] ), 
         .Z(n26711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam addr_23__bdd_3_lut_24114.init = 16'hcaca;
    LUT4 i1_4_lut_adj_465 (.A(is_writing), .B(\fsm_state[0] ), .C(n24484), 
         .D(n27312), .Z(clk_c_enable_355)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_465.init = 16'h1000;
    LUT4 i1_2_lut_adj_466 (.A(read_cycles_count[0]), .B(\read_cycles_count[1] ), 
         .Z(n24484)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_466.init = 16'h4444;
    LUT4 i2890_4_lut (.A(n27253), .B(n27081), .C(n27299), .D(n5), .Z(n5508)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i2890_4_lut.init = 16'hac0c;
    LUT4 i12393_4_lut (.A(nibbles_remaining[0]), .B(n1102), .C(n24382), 
         .D(n8989), .Z(n1094)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i12393_4_lut.init = 16'hcddd;
    LUT4 i23161_3_lut_4_lut (.A(\instr_data[9] ), .B(n27225), .C(n27221), 
         .D(n24704), .Z(instr_data_15__N_1959[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(231[22] 237[16])
    defparam i23161_3_lut_4_lut.init = 16'h8f80;
    LUT4 i23163_3_lut_4_lut (.A(\instr_data[10] ), .B(n27225), .C(n27221), 
         .D(n24707), .Z(instr_data_15__N_1959[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(231[22] 237[16])
    defparam i23163_3_lut_4_lut.init = 16'h8f80;
    LUT4 i2891_4_lut (.A(n27253), .B(n5501), .C(n27299), .D(n5), .Z(n5505)) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i2891_4_lut.init = 16'haccc;
    LUT4 mux_674_i1_4_lut (.A(n356[0]), .B(\addr_in[24] ), .C(n1102), 
         .D(n14701), .Z(n1085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam mux_674_i1_4_lut.init = 16'hcfca;
    LUT4 i23537_4_lut (.A(n5), .B(debug_stall_txn), .C(\read_cycles_count[1] ), 
         .D(data_stall), .Z(n14701)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i23537_4_lut.init = 16'h0001;
    LUT4 i20_4_lut (.A(n27285), .B(n27221), .C(is_writing), .D(n6), 
         .Z(clk_c_enable_415)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;
    defparam i20_4_lut.init = 16'hf535;
    LUT4 i23613_4_lut (.A(is_writing), .B(n27221), .C(qspi_data_byte_idx[1]), 
         .D(n5909), .Z(n25112)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(238[18] 244[12])
    defparam i23613_4_lut.init = 16'h7557;
    PFUMX data_out_7__I_0_242_i8 (.BLUT(instr_data_15__N_1959[31]), .ALUT(data_out_7__N_2273[7]), 
          .C0(n25112), .Z(data_out_7__N_2177[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i7 (.BLUT(instr_data_15__N_1959[30]), .ALUT(data_out_7__N_2273[6]), 
          .C0(n25112), .Z(data_out_7__N_2177[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i6 (.BLUT(instr_data_15__N_1959[29]), .ALUT(data_out_7__N_2273[5]), 
          .C0(n25112), .Z(data_out_7__N_2177[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i5 (.BLUT(instr_data_15__N_1959[28]), .ALUT(data_out_7__N_2273[4]), 
          .C0(n25112), .Z(data_out_7__N_2177[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 i1_4_lut_adj_467 (.A(n4772[1]), .B(n22112), .C(n8989), .D(n5), 
         .Z(n22992)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(209[30] 211[24])
    defparam i1_4_lut_adj_467.init = 16'h8000;
    LUT4 i23540_4_lut (.A(n5), .B(stop_txn_now_N_2363), .C(n23358), .D(rst_reg_n), 
         .Z(n23078)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i23540_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_468 (.A(spi_clk_pos), .B(n27313), .C(n14670), 
         .D(n27284), .Z(n22112)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[25:140])
    defparam i1_2_lut_4_lut_adj_468.init = 16'h00a3;
    LUT4 i23159_3_lut_4_lut (.A(\instr_data[8] ), .B(n27264), .C(n27221), 
         .D(n24701), .Z(instr_data_15__N_1959[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam i23159_3_lut_4_lut.init = 16'h8f80;
    LUT4 i23165_3_lut_4_lut (.A(\instr_data[11] ), .B(n27264), .C(n27221), 
         .D(n24710), .Z(instr_data_15__N_1959[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam i23165_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_4_lut_adj_469 (.A(\fsm_state[0] ), .B(stop_txn_reg), .C(fsm_state[1]), 
         .D(fsm_state[2]), .Z(n23376)) /* synthesis lut_function=(A (B)+!A (B+(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam i1_4_lut_adj_469.init = 16'hdccd;
    LUT4 i12844_3_lut_rep_596_4_lut_3_lut (.A(n27284), .B(n5), .C(spi_clk_pos), 
         .Z(n27221)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(231[22] 237[16])
    defparam i12844_3_lut_rep_596_4_lut_3_lut.init = 16'h8c8c;
    LUT4 n9_bdd_3_lut_24317_4_lut (.A(fsm_state[1]), .B(n27285), .C(spi_in_buffer[1]), 
         .D(qspi_data_out_3__N_5_c[1]), .Z(n26948)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[102:126])
    defparam n9_bdd_3_lut_24317_4_lut.init = 16'hf1e0;
    LUT4 n15156_bdd_3_lut_24256_4_lut (.A(n27283), .B(n27284), .C(rst_reg_n), 
         .D(qspi_data_in[2]), .Z(n26944)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam n15156_bdd_3_lut_24256_4_lut.init = 16'h4000;
    LUT4 n15156_bdd_3_lut_24247_4_lut (.A(n27283), .B(n27284), .C(rst_reg_n), 
         .D(qspi_data_in[3]), .Z(n26938)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam n15156_bdd_3_lut_24247_4_lut.init = 16'h4000;
    LUT4 n15156_bdd_3_lut_23773_4_lut (.A(n27283), .B(n27284), .C(rst_reg_n), 
         .D(qspi_data_in[0]), .Z(n26129)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam n15156_bdd_3_lut_23773_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_470 (.A(n10), .B(debug_stall_txn), .C(is_writing), 
         .D(data_stall), .Z(data_ready_N_2338)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_470.init = 16'h0002;
    LUT4 i21_4_lut (.A(n27310), .B(\read_cycles_count[1] ), .C(n5), .D(n22112), 
         .Z(n10)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A !(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(165[26] 212[20])
    defparam i21_4_lut.init = 16'ha303;
    PFUMX i24356 (.BLUT(n27410), .ALUT(n27411), .C0(n27378), .Z(n27412));
    L6MUX21 i24265 (.D0(n26952), .D1(n26949), .SD(n25112), .Z(data_out_7__N_2177[1]));
    PFUMX i24263 (.BLUT(n26951), .ALUT(n26950), .C0(n27221), .Z(n26952));
    PFUMX i24261 (.BLUT(n24691), .ALUT(n26948), .C0(n27370), .Z(n26949));
    L6MUX21 i24259 (.D0(n26946), .D1(n26943), .SD(n25112), .Z(data_out_7__N_2177[2]));
    PFUMX i24257 (.BLUT(n26945), .ALUT(n26944), .C0(n27221), .Z(n26946));
    PFUMX i24253 (.BLUT(n24694), .ALUT(n26942), .C0(n27370), .Z(n26943));
    L6MUX21 i24250 (.D0(n26940), .D1(n26937), .SD(n25112), .Z(data_out_7__N_2177[3]));
    PFUMX i24248 (.BLUT(n26939), .ALUT(n26938), .C0(n27221), .Z(n26940));
    PFUMX i24245 (.BLUT(n24697), .ALUT(n26936), .C0(n27370), .Z(n26937));
    
endmodule
//
// Verilog Description of module tinyqv_cpu
//

module tinyqv_cpu (clk_c, instr_len, VCC_net, interrupt_core, data_to_write, 
            n2055, qv_data_read_n, \instr_addr_23__N_318[0] , addr, 
            debug_data_continue, counter_hi, debug_instr_valid, was_early_branch, 
            n2035, \pc[2] , \pc[10] , mem_data_ready, n27106, data_ready_sync, 
            \pc[1] , n2096, n2101, n28575, rst_reg_n, instr_data, 
            \data_txn_len[0] , \qspi_data_buf[12] , n27150, \qspi_data_buf[8] , 
            \qspi_data_buf[14] , \qspi_data_buf[10] , \imm[23] , n4057, 
            n26794, n26793, n27298, \imm[22] , \imm[1] , \imm[10] , 
            instr_fetch_running, \imm[21] , \imm[20] , \imm[6] , \imm[19] , 
            \imm[18] , \imm[17] , qv_data_write_n, \imm[16] , \imm[15] , 
            \imm[14] , \imm[13] , \imm[12] , \imm[11] , \imm[9] , 
            \imm[8] , \imm[7] , \imm[5] , \imm[4] , \imm[3] , \imm[2] , 
            is_timer_addr, n27354, n27342, \addr_out[1] , \instr_write_offset[3] , 
            \next_instr_write_offset[3] , n27297, n26730, \mem_data_from_read[4] , 
            mem_op_increment_reg, n24804, n26714, \mem_data_from_read[6] , 
            \mem_data_from_read[27] , \mem_data_from_read[31] , \pc[23] , 
            debug_stop_txn_N_2148, debug_stop_txn_N_2147, \next_pc_for_core[6] , 
            n24747, n24753, \next_pc_for_core[4] , \next_pc_for_core[9] , 
            \next_pc_for_core[13] , n24778, n25239, \pc[8] , \pc[12] , 
            \next_pc_for_core[3] , \next_pc_for_core[5] , \pc[4] , \next_pc_for_core[7] , 
            \next_pc_for_core[8] , \next_pc_for_core[10] , \next_pc_for_core[12] , 
            \next_pc_for_core[11] , \next_pc_for_core[14] , \next_pc_for_core[15] , 
            \next_pc_for_core[16] , \next_pc_for_core[17] , \next_pc_for_core[18] , 
            \next_pc_for_core[19] , \next_pc_for_core[20] , \next_pc_for_core[21] , 
            \next_pc_for_core[22] , \next_pc_for_core[23] , \pc[22] , 
            \pc[21] , \pc[20] , \pc[19] , \pc[18] , \pc[17] , \pc[16] , 
            \pc[15] , \pc[14] , \pc[13] , \pc[11] , \pc[9] , \pc[7] , 
            \pc[6] , \pc[5] , \pc[3] , \mem_data_from_read[19] , \mem_data_from_read[23] , 
            n24757, n27327, \mem_data_from_read[16] , \mem_data_from_read[20] , 
            n24745, \mem_data_from_read[18] , \mem_data_from_read[22] , 
            n24751, n27127, n27333, n27334, n27110, n27341, cycle, 
            n27227, start_instr, n23432, n27350, \early_branch_addr[3] , 
            \early_branch_addr[6] , \early_branch_addr[2] , \early_branch_addr[5] , 
            \early_branch_addr[4] , \early_branch_addr[7] , \early_branch_addr[8] , 
            \early_branch_addr[9] , \early_branch_addr[10] , \early_branch_addr[11] , 
            \early_branch_addr[12] , \early_branch_addr[13] , \early_branch_addr[14] , 
            \early_branch_addr[15] , \early_branch_addr[16] , \early_branch_addr[17] , 
            \early_branch_addr[18] , \early_branch_addr[19] , \early_branch_addr[20] , 
            \early_branch_addr[21] , \early_branch_addr[22] , \early_branch_addr[23] , 
            n44, \data_from_read[2] , n27294, n10, n27093, n27277, 
            n23526, n22591, n9091, n23532, n27306, n24742, n24743, 
            n24744, n23536, \mem_data_from_read[1] , \mem_data_from_read[5] , 
            \mem_data_from_read[9] , \mem_data_from_read[13] , \data_from_read[6] , 
            instr_fetch_running_N_945, instr_fetch_stopped, \instr_addr[2] , 
            n24759, n27268, \mem_data_from_read[24] , \mem_data_from_read[28] , 
            \mem_data_from_read[26] , \mem_data_from_read[30] , n24126, 
            n27241, n27255, \qspi_data_buf[25] , \qspi_data_buf[29] , 
            \mem_data_from_read[17] , \mem_data_from_read[21] , n27233, 
            n8869, n27279, n23908, n27358, n27220, mem_op_increment_reg_de, 
            n27218, \next_fsm_state_3__N_2499[3] , clk_c_enable_350, clk_c_enable_367, 
            \debug_branch_N_840[29] , \mul_out[2] , \mul_out[3] , \mul_out[1] , 
            \ui_in_sync[1] , n1167, debug_rd, accum, d_3__N_1868, 
            n4577, n26802, n27223, \next_accum[5] , \next_accum[6] , 
            \next_accum[7] , GND_net, \next_accum[8] , \next_accum[9] , 
            \next_accum[10] , \next_accum[11] , \next_accum[12] , \next_accum[13] , 
            \next_accum[14] , \next_accum[15] , \next_accum[16] , \next_accum[17] , 
            \next_accum[18] , \next_accum[19] , \next_accum[4] ) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output [2:1]instr_len;
    input VCC_net;
    output interrupt_core;
    output [31:0]data_to_write;
    input n2055;
    output [1:0]qv_data_read_n;
    output \instr_addr_23__N_318[0] ;
    output [27:0]addr;
    output debug_data_continue;
    output [4:2]counter_hi;
    output debug_instr_valid;
    output was_early_branch;
    input n2035;
    output \pc[2] ;
    output \pc[10] ;
    input mem_data_ready;
    output n27106;
    output data_ready_sync;
    output \pc[1] ;
    output n2096;
    output n2101;
    input n28575;
    input rst_reg_n;
    input [15:0]instr_data;
    input \data_txn_len[0] ;
    input \qspi_data_buf[12] ;
    input n27150;
    input \qspi_data_buf[8] ;
    input \qspi_data_buf[14] ;
    input \qspi_data_buf[10] ;
    output \imm[23] ;
    output n4057;
    input n26794;
    input n26793;
    input n27298;
    output \imm[22] ;
    output \imm[1] ;
    output \imm[10] ;
    output instr_fetch_running;
    output \imm[21] ;
    output \imm[20] ;
    output \imm[6] ;
    output \imm[19] ;
    output \imm[18] ;
    output \imm[17] ;
    output [1:0]qv_data_write_n;
    output \imm[16] ;
    output \imm[15] ;
    output \imm[14] ;
    output \imm[13] ;
    output \imm[12] ;
    output \imm[11] ;
    output \imm[9] ;
    output \imm[8] ;
    output \imm[7] ;
    output \imm[5] ;
    output \imm[4] ;
    output \imm[3] ;
    output \imm[2] ;
    output is_timer_addr;
    output n27354;
    output n27342;
    output \addr_out[1] ;
    output \instr_write_offset[3] ;
    output \next_instr_write_offset[3] ;
    output n27297;
    input n26730;
    input \mem_data_from_read[4] ;
    output mem_op_increment_reg;
    input n24804;
    input n26714;
    input \mem_data_from_read[6] ;
    input \mem_data_from_read[27] ;
    input \mem_data_from_read[31] ;
    output \pc[23] ;
    input debug_stop_txn_N_2148;
    output debug_stop_txn_N_2147;
    input \next_pc_for_core[6] ;
    input n24747;
    input n24753;
    input \next_pc_for_core[4] ;
    input \next_pc_for_core[9] ;
    input \next_pc_for_core[13] ;
    input n24778;
    output n25239;
    output \pc[8] ;
    output \pc[12] ;
    input \next_pc_for_core[3] ;
    input \next_pc_for_core[5] ;
    output \pc[4] ;
    input \next_pc_for_core[7] ;
    input \next_pc_for_core[8] ;
    input \next_pc_for_core[10] ;
    input \next_pc_for_core[12] ;
    input \next_pc_for_core[11] ;
    input \next_pc_for_core[14] ;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[16] ;
    input \next_pc_for_core[17] ;
    input \next_pc_for_core[18] ;
    input \next_pc_for_core[19] ;
    input \next_pc_for_core[20] ;
    input \next_pc_for_core[21] ;
    input \next_pc_for_core[22] ;
    input \next_pc_for_core[23] ;
    output \pc[22] ;
    output \pc[21] ;
    output \pc[20] ;
    output \pc[19] ;
    output \pc[18] ;
    output \pc[17] ;
    output \pc[16] ;
    output \pc[15] ;
    output \pc[14] ;
    output \pc[13] ;
    output \pc[11] ;
    output \pc[9] ;
    output \pc[7] ;
    output \pc[6] ;
    output \pc[5] ;
    output \pc[3] ;
    input \mem_data_from_read[19] ;
    input \mem_data_from_read[23] ;
    output n24757;
    output n27327;
    input \mem_data_from_read[16] ;
    input \mem_data_from_read[20] ;
    output n24745;
    input \mem_data_from_read[18] ;
    input \mem_data_from_read[22] ;
    output n24751;
    input n27127;
    output n27333;
    output n27334;
    output n27110;
    output n27341;
    output [1:0]cycle;
    input n27227;
    output start_instr;
    input n23432;
    output n27350;
    input \early_branch_addr[3] ;
    input \early_branch_addr[6] ;
    input \early_branch_addr[2] ;
    input \early_branch_addr[5] ;
    input \early_branch_addr[4] ;
    input \early_branch_addr[7] ;
    input \early_branch_addr[8] ;
    input \early_branch_addr[9] ;
    input \early_branch_addr[10] ;
    input \early_branch_addr[11] ;
    input \early_branch_addr[12] ;
    input \early_branch_addr[13] ;
    input \early_branch_addr[14] ;
    input \early_branch_addr[15] ;
    input \early_branch_addr[16] ;
    input \early_branch_addr[17] ;
    input \early_branch_addr[18] ;
    input \early_branch_addr[19] ;
    input \early_branch_addr[20] ;
    input \early_branch_addr[21] ;
    input \early_branch_addr[22] ;
    input \early_branch_addr[23] ;
    input n44;
    input \data_from_read[2] ;
    input n27294;
    input n10;
    output n27093;
    input n27277;
    input n23526;
    output n22591;
    input n9091;
    input n23532;
    output n27306;
    input n24742;
    input n24743;
    output n24744;
    input n23536;
    input \mem_data_from_read[1] ;
    input \mem_data_from_read[5] ;
    input \mem_data_from_read[9] ;
    input \mem_data_from_read[13] ;
    input \data_from_read[6] ;
    input instr_fetch_running_N_945;
    input instr_fetch_stopped;
    output \instr_addr[2] ;
    input n24759;
    input n27268;
    input \mem_data_from_read[24] ;
    input \mem_data_from_read[28] ;
    input \mem_data_from_read[26] ;
    input \mem_data_from_read[30] ;
    input n24126;
    input n27241;
    input n27255;
    input \qspi_data_buf[25] ;
    input \qspi_data_buf[29] ;
    input \mem_data_from_read[17] ;
    input \mem_data_from_read[21] ;
    output n27233;
    input n8869;
    output n27279;
    output n23908;
    input n27358;
    input n27220;
    output mem_op_increment_reg_de;
    output n27218;
    input \next_fsm_state_3__N_2499[3] ;
    input clk_c_enable_350;
    input clk_c_enable_367;
    input \debug_branch_N_840[29] ;
    input \mul_out[2] ;
    input \mul_out[3] ;
    input \mul_out[1] ;
    input \ui_in_sync[1] ;
    output n1167;
    output [3:0]debug_rd;
    output [15:0]accum;
    output [19:0]d_3__N_1868;
    input n4577;
    input n26802;
    input n27223;
    input \next_accum[5] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input GND_net;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[4] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [3:0]rs1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(117[15:18])
    
    wire clk_c_enable_282;
    wire [3:0]n2175;
    wire [2:0]mem_op;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(115[15:21])
    wire [2:0]mem_op_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(65[16:25])
    
    wire clk_c_enable_26, n27151;
    wire [3:0]rd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(119[15:17])
    
    wire clk_c_enable_372;
    wire [3:0]n2386;
    wire [3:0]alu_op;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    
    wire n27326;
    wire [3:0]alu_op_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(64[16:25])
    
    wire data_ready_latch, clk_c_enable_14, n23201, load_started, address_ready, 
        n856, clk_c_enable_90, n27112, clk_c_enable_20, n27214;
    wire [31:0]imm;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(100[16:19])
    
    wire clk_c_enable_227;
    wire [31:0]n3438;
    wire [3:0]data_out_slice;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(230[16:30])
    
    wire n27222, clk_c_enable_31;
    wire [15:0]n1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]n5;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]n1735;
    
    wire clk_c_enable_67, clk_c_enable_40;
    wire [2:1]instr_len_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(113[15:24])
    
    wire clk_c_enable_34, n27147, clk_c_enable_280, n22867, clk_c_enable_49;
    wire [2:0]additional_mem_ops;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(120[15:33])
    wire [2:0]additional_mem_ops_2__N_749;
    
    wire clk_c_enable_175;
    wire [63:0]instr_data_0__15__N_638;
    wire [2:0]instr_write_offset_3__N_934;
    
    wire clk_c_enable_272;
    wire [27:0]addr_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(131[17:25])
    
    wire n27145, n26874, n4075, n26875, clk_c_enable_56, clk_c_enable_53, 
        data_continue_N_963, clk_c_enable_60, clk_c_enable_64, n27338, 
        n26868, n26867, n25707, n26869;
    wire [3:2]addr_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(121[15:26])
    wire [1:0]n21;
    
    wire debug_instr_valid_N_436, n26857, n26856, n25708, n22, is_alu_imm, 
        clk_c_enable_242, is_alu_imm_de, n26854, n26853, n26855, is_jalr, 
        is_jalr_de, clk_c_enable_100, debug_early_branch;
    wire [15:0]n31;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]n33;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire n24629, n26197, n26819, n26818, n26820, is_system, n27276, 
        n27231, n23682, n27209, n27109, n24817, data_ready_core;
    wire [17:16]mip_reg;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(321[17:24])
    wire [3:0]csr_read_3__N_1459;
    
    wire n27211, n27198, n23698, clk_c_enable_115;
    wire [31:0]n3397;
    
    wire n26263, n4079, n26264, clk_c_enable_117, clk_c_enable_142, 
        n27396, n27395, n26807, n26806, n28564, n19, n27400, n23506, 
        n27096, n10_c, n27095, n26804, n26803, n27212, n26805, 
        n27399;
    wire [31:0]instr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(47[17:22])
    
    wire n27131;
    wire [30:0]n4703;
    
    wire n27403, n27402;
    wire [31:0]n3350;
    
    wire n26304, n23608, n6, n27103, n23614, n27099, n27260, n24998, 
        is_alu_reg, is_alu_reg_de, n23618, n23624, clk_c_enable_144, 
        clk_c_enable_158, clk_c_enable_160, clk_c_enable_174, n26277, 
        n26280, n26795, n23628, n23634, n24666, is_auipc, is_auipc_de, 
        n26282, n26283, n27330, n24360, n23498, n27123, n27101, 
        clk_c_enable_209, n5590, n26289, n26292, n4073, n4065, n27085, 
        is_system_de;
    wire [31:0]n3163;
    wire [31:0]n2874;
    wire [31:0]n3314;
    
    wire n27374, n27287, n27247, n27, n2700, n26300, n26295, n8900, 
        n22088, n24160, n22178, n22090, n23544, n16, n2029;
    wire [15:0]n1715;
    
    wire n22534, n27086, n24976, clk_c_enable_278;
    wire [1:0]data_write_n_1__N_369;
    
    wire is_lui, is_lui_de, is_store, is_store_de, n23638, n23644, 
        clk_c_enable_229, n27108, n27114, no_write_in_progress, clk_c_enable_231, 
        no_write_in_progress_N_471, is_branch, is_branch_de, n24668;
    wire [3:0]rs2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(118[15:18])
    wire [3:0]n1815;
    
    wire clk_c_enable_245, n22885, n26294, n27102, is_load, is_load_de, 
        is_jal, is_jal_de, n25199, n25198, n25197, n25196, n26119, 
        n26297, n25192, n25191, n26202, n26201, n26203;
    wire [59:0]debug_branch_N_840;
    wire [3:0]timer_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(143[16:26])
    wire [3:0]debug_branch_N_450;
    
    wire n23980, n23087, n27289, n12, stall_core, n27288, n14783, 
        n25190, n25189, n23838, n2704, n25185, n26732, n26728, 
        n26733, n23045;
    wire [1:0]n699;
    
    wire n22226;
    wire [22:0]instr_addr_23__N_318;
    
    wire n26299, n27355, n4, n25184, n25183, n2, n9, n26731, 
        n23398, n23402, instr_complete_N_1647, n25182, n25178, n25177, 
        n25176, n25175, n27347, n27302, n15_adj_2637, n25132, n27142, 
        n28563, n28140, clk_c_enable_275, n27111, n27107;
    wire [15:0]n2036;
    wire [15:0]n2056;
    
    wire n28142, n27148, n29, n27226, n26196, n26198, n26716, 
        n26712, n26717, n26317, n24752, load_top_bit, data_out_3__N_1385, 
        n24664, n24746, n27023;
    wire [59:0]debug_rd_3__N_405;
    
    wire n27319, n7717;
    wire [59:0]debug_branch_N_446;
    
    wire n24658, n22898, n23600, n8, n22816, n26316, clk_c_enable_424;
    wire [6:0]cycle_count_wide;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(279[16:32])
    wire [2:0]time_hi;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(292[15:22])
    
    wire n26926, n22499, n23928, n26715, n22369, n27113, n22866, 
        instr_fetch_restart_N_947, n27179, n4_adj_2638, n8274, n23690;
    wire [3:0]time_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(299[16:26])
    
    wire mstatus_mie, interrupt_pending_N_1671, n23292, any_additional_mem_ops;
    wire [2:0]n4116;
    
    wire n26345, n26346, n26932, n26177, n26176, n26178;
    wire [16:0]mie;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(323[16:19])
    
    wire n26336;
    wire [3:0]n5167;
    
    wire n26335, n22080, n24, n23894;
    wire [31:0]n3273;
    
    wire n24505;
    wire [2:0]n34;
    
    wire n24625, n24900, n24627, n24635, n27163, n27167, n23602;
    wire [3:1]next_pc_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[16:30])
    
    wire n24633, n24641, n24758, clk_c_enable_423;
    wire [20:0]pc_23__N_911;
    
    wire n22592, n27097, n26, n24984, n24509, n27353, n24775, 
        debug_ret;
    wire [23:1]return_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(135[17:28])
    wire [1:0]n1768;
    
    wire n9111, n27190, n27132, is_lui_N_1365;
    wire [12:0]n4745;
    
    wire n9115, n27205, n27191, n23462, n27160, n22671, n23470, 
        n22667, n23478, n22663, n28562, n27189, n27135, n27203, 
        n25083, n27084, n4071, n22745, n23522, n27204, n23516, 
        n24631, n26432, n27202, n26433, n23848, n2031, n22704, 
        n22_adj_2640;
    wire [31:0]n3087;
    
    wire n26434, n23656, n2702, n27199, n23868, n24030, n23738, 
        n149, n24642, n27200, n26116, n24773, n27201, n27175, 
        n15_adj_2641, n25142;
    wire [3:0]n234;
    wire [3:0]debug_rd_3__N_1567;
    wire [1:0]pc_2__N_932;
    
    wire n22715, n25, n24638, n24780, n14587, n37, n22700, n24637, 
        n209, n27293, n24959, n24616, n27140, debug_rd_3__N_413;
    wire [31:0]n3196;
    
    wire n22748;
    wire [3:0]n2161;
    
    wire n2330, n27092, n25237, n26822, n27376, n27305, n27332, 
        n27256, n24612;
    wire [3:0]data_rs1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(83[16:24])
    
    wire alu_a_in_3__N_1552;
    wire [59:0]debug_branch_N_442;
    
    wire cy, n27228, cy_adj_2642, instr_retired, n27246, n157, n35, 
        n27128, n26028, n26027, n4063, n26029;
    wire [4:0]increment_result_3__N_1911;
    
    wire n27124;
    wire [20:0]n36;
    
    wire n26976;
    wire [3:0]n1794;
    wire [5:0]mcause;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(325[15:21])
    
    wire n26930, n149_adj_2643, n26927, n27329, n157_adj_2644, n16_adj_2645, 
        cy_adj_2646, n27267, n27252, n22637, n22721, n27343;
    wire [5:0]n611;
    
    wire n23412, n27088, n23856, n22733, n28, n824, n22559;
    wire [31:0]n3126;
    
    wire n27185, n27184, n7, n24583, n22551, n27197, n26117;
    wire [15:0]n4625;
    
    wire n24_adj_2656, n27372, n27304, n5839;
    wire [31:0]n3232;
    
    wire n24632, n24634, n5868, n22887, n27371, n22888, n22889;
    wire [3:0]n2368;
    wire [3:0]n2376;
    
    wire n25066, n27349, n25069;
    wire [3:0]n2152;
    
    wire n27321, load_done, instr_complete_N_1651, n27170, n22100, 
        n13, n27178, n8_adj_2657, n15_adj_2658, n17, n26_adj_2659, 
        n24525, n22674, n2328, n20, n8486, n16_adj_2660, n11, 
        n2326, n27157;
    wire [2:0]additional_mem_ops_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(70[16:37])
    wire [3:0]n2120;
    wire [3:0]n2128;
    
    wire n23564, n22784, n27152;
    wire [3:0]n2342;
    
    wire n27206, n24624, n30, n25004, n5160, n27207, n30_adj_2661, 
        n30_adj_2662;
    wire [3:0]n2133;
    
    wire n23594, n23726, n24601, n26118, n23572, n23580, n2322;
    wire [3:0]data_rs2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(84[16:24])
    wire [3:0]n92;
    
    wire n28571, n28573, clk_c_enable_276, n27263, n24216, n25702, 
        n25703, n25704, n9124;
    wire [3:0]n2138;
    
    wire n25705, n9675, n27300, n25706, n22121;
    wire [3:0]n1804;
    wire [23:0]mepc;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(68[16:20])
    wire [3:0]csr_read_3__N_1451;
    wire [3:0]n2347;
    
    wire is_ret_de, n23238, n23558, n22909;
    wire [3:0]n2352;
    
    wire n27156, n24640, n24988, n7711;
    wire [3:0]instrret_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(301[16:30])
    wire [3:0]n5114;
    
    wire n6985, debug_reg_wen_N_1692, n27266, n24838, n27270, n27274, 
        n27129, n27292, n27348, n27130, n23658, n23662;
    wire [3:0]alu_b_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[16:24])
    
    wire n27181, n27183;
    wire [3:0]alu_op_3__N_1337;
    
    wire n15_adj_2663, n23678, n27126;
    wire [20:0]n1222;
    
    wire n22739, n27322, n6982, n27138, n32, n27187, n27188, n27215, 
        n27238;
    wire [1:0]n4575;
    
    wire n27158, n26779, n22101, n22_adj_2664, n25179, n25180, n25186, 
        n25187, n25193, n25194, n25200, n25201, n27_adj_2665;
    wire [31:0]data_from_read;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(59[16:30])
    
    wire n27290, n27296, n26435, n26436, n27169, n27173, n24772, 
        n225, n18144, n8_adj_2666, n926, n27362, n24822, n893, 
        n24611, n860, n22164, n8123, n793, n27174, n26175, n27171, 
        n26206, n27176, n27172, n27122, n23792, n24398, n24404, 
        n212, n9117, n27366, n27368, n27275, n27249, n27248, n27367, 
        n27369, n27166, n27390, n27186, n8_adj_2668, n3, n27177;
    wire [31:0]tmp_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(88[16:24])
    
    wire n226, n24774, n25126, n27159, n28141, n27164, n225_adj_2669, 
        n26348, timer_interrupt, load_top_bit_next_N_1731, n15206, mstatus_mte, 
        n5434, n25233, n25234, clk_c_enable_71, clk_c_enable_422, 
        n27245, n27309;
    wire [3:0]csr_read_3__N_1443;
    
    wire n27377;
    wire [5:0]shift_amt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[16:25])
    
    wire n7278;
    wire [3:0]shift_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(132[16:25])
    
    wire n62, n25292, n8153, n8157, n26049, n26685, n26686;
    wire [31:0]a_for_shift_right;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[17:34])
    
    wire n63, n27168, n25014, n24_adj_2670, n25057, n27401, instr_fetch_running_N_943, 
        n27192, n27162, n26195, n23588, n26347, n27121, n26745, 
        n27389, n10_adj_2671, n23, n24599, n24210, n23140, n24198, 
        n24202, n24200, n24182, n24174, n27397, n27244, n23756, 
        n23820, n23824;
    wire [31:0]mtimecmp;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(30[16:24])
    
    wire mtimecmp_2__N_1939, mtimecmp_0__N_1943, n26200, n22778, n23870;
    wire [2:0]n1764;
    
    wire n26318, n28143, n23450, n23804, n23744, n26298, n26296, 
        n23712, debug_rd_3__N_1575, n26821, n27196, n26293, n26290, 
        n24605, n20_adj_2672, n14, n24124, n23768, cmp;
    wire [3:0]alu_a_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[16:24])
    
    wire n23342;
    wire [3:0]mtime_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(29[16:25])
    
    wire n27257, cy_adj_2673, n27219, time_pulse_r, n27236;
    wire [3:0]tmp_data_in_3__N_1514;
    
    wire n8162, n27154;
    wire [4:0]increment_result_3__N_1925;
    
    wire n27229, mstatus_mpie;
    wire [3:0]csr_read_3__N_1439;
    
    wire n26281, n26278, n27391, mtimecmp_1__N_1941, mtimecmp_3__N_1935, 
        n27180, clk_c_enable_73;
    wire [3:0]\reg_access[4] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(30[16:26])
    wire [3:0]\reg_access[3] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(30[16:26])
    
    wire n23750, n23842, n23798, n23810, n24516, n23650, n23718, 
        n23762, n23774, n23598, n12_adj_2674, n23704;
    
    FD1P3AX rs1_i0_i1 (.D(n2175[1]), .SP(clk_c_enable_282), .CK(clk_c), 
            .Q(rs1[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i1.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i2 (.D(mem_op_de[2]), .SP(clk_c_enable_282), .CK(clk_c), 
            .Q(mem_op[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i2.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i1 (.D(mem_op_de[1]), .SP(clk_c_enable_282), .CK(clk_c), 
            .Q(mem_op[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i1.GSR = "DISABLED";
    FD1P3AX instr_len_i2 (.D(n27151), .SP(clk_c_enable_26), .CK(clk_c), 
            .Q(instr_len[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_len_i2.GSR = "DISABLED";
    FD1P3AX rd_i0_i3 (.D(n2386[3]), .SP(clk_c_enable_372), .CK(clk_c), 
            .Q(rd[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i3.GSR = "DISABLED";
    FD1P3AX rd_i0_i2 (.D(n2386[2]), .SP(clk_c_enable_372), .CK(clk_c), 
            .Q(rd[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i2.GSR = "DISABLED";
    FD1P3AX rd_i0_i1 (.D(n2386[1]), .SP(clk_c_enable_372), .CK(clk_c), 
            .Q(rd[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i1.GSR = "DISABLED";
    FD1P3IX alu_op__i3 (.D(alu_op_de[3]), .SP(clk_c_enable_26), .CD(n27326), 
            .CK(clk_c), .Q(alu_op[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i3.GSR = "DISABLED";
    FD1P3IX alu_op__i2 (.D(alu_op_de[2]), .SP(clk_c_enable_26), .CD(n27326), 
            .CK(clk_c), .Q(alu_op[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i2.GSR = "DISABLED";
    FD1P3IX alu_op__i1 (.D(alu_op_de[1]), .SP(clk_c_enable_26), .CD(n27326), 
            .CK(clk_c), .Q(alu_op[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i1.GSR = "DISABLED";
    FD1P3AX data_ready_latch_416 (.D(n23201), .SP(clk_c_enable_14), .CK(clk_c), 
            .Q(data_ready_latch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(235[12] 256[8])
    defparam data_ready_latch_416.GSR = "DISABLED";
    FD1P3IX load_started_422 (.D(VCC_net), .SP(address_ready), .CD(n856), 
            .CK(clk_c), .Q(load_started)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam load_started_422.GSR = "DISABLED";
    FD1P3IX interrupt_core_408 (.D(n27112), .SP(clk_c_enable_90), .CD(n27326), 
            .CK(clk_c), .Q(interrupt_core)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam interrupt_core_408.GSR = "DISABLED";
    FD1P3IX data_out__i31 (.D(n27214), .SP(clk_c_enable_20), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i31.GSR = "DISABLED";
    FD1P3AX imm_i0_i0 (.D(n3438[0]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(imm[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i0.GSR = "DISABLED";
    FD1P3IX data_out__i30 (.D(data_out_slice[2]), .SP(clk_c_enable_20), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i30.GSR = "DISABLED";
    FD1P3IX data_out__i29 (.D(n27222), .SP(clk_c_enable_20), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i29.GSR = "DISABLED";
    FD1P3IX data_out__i28 (.D(data_out_slice[0]), .SP(clk_c_enable_20), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i28.GSR = "DISABLED";
    FD1P3IX data_out__i27 (.D(n27214), .SP(clk_c_enable_31), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i27.GSR = "DISABLED";
    LUT4 mux_1077_i5_3_lut (.A(n1[4]), .B(n5[4]), .C(n2055), .Z(n1735[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i5_3_lut.init = 16'hcaca;
    FD1P3IX data_out__i0 (.D(data_out_slice[0]), .SP(clk_c_enable_67), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i0.GSR = "DISABLED";
    FD1P3IX alu_op__i0 (.D(alu_op_de[0]), .SP(clk_c_enable_26), .CD(n27326), 
            .CK(clk_c), .Q(alu_op[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i0.GSR = "DISABLED";
    FD1P3IX data_out__i26 (.D(data_out_slice[2]), .SP(clk_c_enable_31), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i26.GSR = "DISABLED";
    FD1P3AX rd_i0_i0 (.D(n2386[0]), .SP(clk_c_enable_372), .CK(clk_c), 
            .Q(rd[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i0.GSR = "DISABLED";
    FD1P3IX data_out__i25 (.D(n27222), .SP(clk_c_enable_31), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i25.GSR = "DISABLED";
    FD1P3IX data_out__i24 (.D(data_out_slice[0]), .SP(clk_c_enable_31), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i24.GSR = "DISABLED";
    FD1P3IX data_out__i23 (.D(n27214), .SP(clk_c_enable_40), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[23])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i23.GSR = "DISABLED";
    FD1P3IX data_out__i22 (.D(data_out_slice[2]), .SP(clk_c_enable_40), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[22])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i22.GSR = "DISABLED";
    FD1P3IX instr_len_i1 (.D(n27147), .SP(clk_c_enable_34), .CD(n27326), 
            .CK(clk_c), .Q(instr_len_c[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_len_i1.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i0 (.D(mem_op_de[0]), .SP(clk_c_enable_282), .CK(clk_c), 
            .Q(mem_op[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i0.GSR = "DISABLED";
    FD1P3AX rs1_i0_i0 (.D(n2175[0]), .SP(clk_c_enable_282), .CK(clk_c), 
            .Q(rs1[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i0.GSR = "DISABLED";
    FD1P3AX data_read_n_i0_i0 (.D(n22867), .SP(clk_c_enable_280), .CK(clk_c), 
            .Q(qv_data_read_n[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_read_n_i0_i0.GSR = "DISABLED";
    FD1P3IX data_out__i21 (.D(n27222), .SP(clk_c_enable_40), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[21])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i21.GSR = "DISABLED";
    FD1P3IX data_out__i20 (.D(data_out_slice[0]), .SP(clk_c_enable_40), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[20])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i20.GSR = "DISABLED";
    FD1P3IX data_out__i19 (.D(n27214), .SP(clk_c_enable_49), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[19])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i19.GSR = "DISABLED";
    FD1P3IX data_out__i18 (.D(data_out_slice[2]), .SP(clk_c_enable_49), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[18])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i18.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i0 (.D(additional_mem_ops_2__N_749[0]), .CK(clk_c), 
            .CD(n27326), .Q(additional_mem_ops[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i0.GSR = "DISABLED";
    FD1P3AX instr_data_3__i1 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_175), 
            .CK(clk_c), .Q(n1[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i1.GSR = "DISABLED";
    FD1P3IX data_out__i17 (.D(n27222), .SP(clk_c_enable_49), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[17])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i17.GSR = "DISABLED";
    FD1P3IX data_out__i16 (.D(data_out_slice[0]), .SP(clk_c_enable_49), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[16])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i16.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i1 (.D(instr_write_offset_3__N_934[0]), .CK(clk_c), 
            .CD(n27326), .Q(\instr_addr_23__N_318[0] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i1.GSR = "DISABLED";
    FD1P3IX data_addr__i0 (.D(addr_out[0]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i0.GSR = "DISABLED";
    PFUMX i24215 (.BLUT(n27145), .ALUT(n26874), .C0(n4075), .Z(n26875));
    FD1P3IX data_out__i15 (.D(n27214), .SP(clk_c_enable_56), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i15.GSR = "DISABLED";
    FD1P3IX data_out__i14 (.D(data_out_slice[2]), .SP(clk_c_enable_56), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i14.GSR = "DISABLED";
    FD1P3AX data_continue_420 (.D(data_continue_N_963), .SP(clk_c_enable_53), 
            .CK(clk_c), .Q(debug_data_continue)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_continue_420.GSR = "DISABLED";
    FD1P3IX data_out__i13 (.D(n27222), .SP(clk_c_enable_56), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i13.GSR = "DISABLED";
    FD1P3IX data_out__i12 (.D(data_out_slice[0]), .SP(clk_c_enable_56), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i12.GSR = "DISABLED";
    FD1P3IX data_out__i11 (.D(n27214), .SP(clk_c_enable_60), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i11.GSR = "DISABLED";
    FD1P3IX data_out__i10 (.D(data_out_slice[2]), .SP(clk_c_enable_60), 
            .CD(n27326), .CK(clk_c), .Q(data_to_write[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i10.GSR = "DISABLED";
    FD1P3IX data_out__i9 (.D(n27222), .SP(clk_c_enable_60), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i9.GSR = "DISABLED";
    FD1P3IX data_out__i8 (.D(data_out_slice[0]), .SP(clk_c_enable_60), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i8.GSR = "DISABLED";
    FD1P3IX data_out__i7 (.D(n27214), .SP(clk_c_enable_64), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i7.GSR = "DISABLED";
    FD1P3IX data_out__i6 (.D(data_out_slice[2]), .SP(clk_c_enable_64), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i6.GSR = "DISABLED";
    FD1P3IX data_out__i5 (.D(n27222), .SP(clk_c_enable_64), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i5.GSR = "DISABLED";
    FD1P3IX data_out__i4 (.D(data_out_slice[0]), .SP(clk_c_enable_64), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i4.GSR = "DISABLED";
    FD1P3IX data_out__i3 (.D(n27214), .SP(clk_c_enable_67), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i3.GSR = "DISABLED";
    FD1S3IX counter_hi_3236__i2 (.D(n27338), .CK(clk_c), .CD(n27326), 
            .Q(counter_hi[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3236__i2.GSR = "DISABLED";
    FD1P3IX data_out__i2 (.D(data_out_slice[2]), .SP(clk_c_enable_67), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i2.GSR = "DISABLED";
    FD1P3IX data_out__i1 (.D(n27222), .SP(clk_c_enable_67), .CD(n27326), 
            .CK(clk_c), .Q(data_to_write[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i1.GSR = "DISABLED";
    PFUMX i24211 (.BLUT(n26868), .ALUT(n26867), .C0(n25707), .Z(n26869));
    FD1S3IX addr_offset_3237__i2 (.D(n21[0]), .CK(clk_c), .CD(n27326), 
            .Q(addr_offset[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam addr_offset_3237__i2.GSR = "DISABLED";
    FD1P3IX instr_valid_392 (.D(debug_instr_valid_N_436), .SP(clk_c_enable_90), 
            .CD(n27326), .CK(clk_c), .Q(debug_instr_valid)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_valid_392.GSR = "DISABLED";
    PFUMX i24203 (.BLUT(n26857), .ALUT(n26856), .C0(n25708), .Z(n22));
    FD1P3IX is_alu_imm_394 (.D(is_alu_imm_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_alu_imm)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_alu_imm_394.GSR = "DISABLED";
    PFUMX i24200 (.BLUT(n26854), .ALUT(n26853), .C0(counter_hi[2]), .Z(n26855));
    FD1P3IX is_jalr_400 (.D(is_jalr_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_jalr)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_jalr_400.GSR = "DISABLED";
    FD1P3IX was_early_branch_424 (.D(debug_early_branch), .SP(clk_c_enable_100), 
            .CD(n27326), .CK(clk_c), .Q(was_early_branch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(315[12] 320[8])
    defparam was_early_branch_424.GSR = "DISABLED";
    LUT4 mux_1073_i5_rep_86_3_lut (.A(n31[4]), .B(n33[4]), .C(n2035), 
         .Z(n24629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i5_rep_86_3_lut.init = 16'hcaca;
    LUT4 pc_2__bdd_3_lut_24466 (.A(\pc[2] ), .B(\pc[10] ), .C(counter_hi[3]), 
         .Z(n26197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_2__bdd_3_lut_24466.init = 16'hcaca;
    PFUMX i24176 (.BLUT(n26819), .ALUT(n26818), .C0(mem_data_ready), .Z(n26820));
    LUT4 is_csr_I_0_573_2_lut_rep_651_3_lut_4_lut_3_lut_4_lut (.A(alu_op[1]), 
         .B(alu_op[0]), .C(is_system), .D(debug_instr_valid), .Z(n27276)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_csr_I_0_573_2_lut_rep_651_3_lut_4_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i7286_2_lut_rep_606_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut (.A(alu_op[1]), 
         .B(alu_op[0]), .C(is_system), .D(debug_instr_valid), .Z(n27231)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i7286_2_lut_rep_606_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h6000;
    LUT4 i23467_2_lut_3_lut_4_lut (.A(n23682), .B(n27106), .C(n27209), 
         .D(n27109), .Z(n24817)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i23467_2_lut_3_lut_4_lut.init = 16'hffbf;
    FD1S3IX data_ready_sync_415 (.D(data_ready_core), .CK(clk_c), .CD(n27326), 
            .Q(data_ready_sync)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(235[12] 256[8])
    defparam data_ready_sync_415.GSR = "DISABLED";
    LUT4 i1339_2_lut_3_lut_4_lut_4_lut (.A(instr_len[2]), .B(\pc[2] ), .C(\pc[1] ), 
         .D(instr_len_c[1]), .Z(n2096)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A ((C (D)+!C !(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1339_2_lut_3_lut_4_lut_4_lut.init = 16'h0660;
    LUT4 i1344_2_lut_3_lut_4_lut_4_lut (.A(instr_len[2]), .B(\pc[2] ), .C(\pc[1] ), 
         .D(instr_len_c[1]), .Z(n2101)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (B+(C (D)+!C !(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1344_2_lut_3_lut_4_lut_4_lut.init = 16'h0990;
    LUT4 i12308_2_lut_3_lut_4_lut_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .D(mip_reg[17]), .Z(csr_read_3__N_1459[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i12308_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 i12348_2_lut_3_lut_4_lut_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .D(mip_reg[16]), .Z(csr_read_3__N_1459[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i12348_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 i442_2_lut_rep_469_3_lut_4_lut (.A(n23682), .B(n27106), .C(n28575), 
         .D(n27109), .Z(clk_c_enable_282)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i442_2_lut_rep_469_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_3_lut (.A(n27211), .B(n27198), .C(rst_reg_n), .Z(n23698)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4040;
    FD1P3AX instr_data_3__i64 (.D(instr_data[15]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i64.GSR = "DISABLED";
    LUT4 n3412_bdd_3_lut_23858 (.A(n3397[17]), .B(n26263), .C(n4079), 
         .Z(n26264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3412_bdd_3_lut_23858.init = 16'hcaca;
    FD1P3AX instr_data_3__i63 (.D(instr_data[14]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i63.GSR = "DISABLED";
    FD1P3AX instr_data_3__i62 (.D(instr_data[13]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i62.GSR = "DISABLED";
    FD1P3AX instr_data_3__i61 (.D(instr_data[12]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i61.GSR = "DISABLED";
    FD1P3AX instr_data_3__i60 (.D(instr_data[11]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i60.GSR = "DISABLED";
    FD1P3AX instr_data_3__i59 (.D(instr_data[10]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i59.GSR = "DISABLED";
    FD1P3AX instr_data_3__i58 (.D(instr_data[9]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i58.GSR = "DISABLED";
    FD1P3AX instr_data_3__i57 (.D(instr_data[8]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i57.GSR = "DISABLED";
    FD1P3AX instr_data_3__i56 (.D(instr_data[7]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i56.GSR = "DISABLED";
    FD1P3AX instr_data_3__i55 (.D(instr_data[6]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i55.GSR = "DISABLED";
    FD1P3AX instr_data_3__i54 (.D(instr_data[5]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i54.GSR = "DISABLED";
    FD1P3AX instr_data_3__i53 (.D(instr_data[4]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i53.GSR = "DISABLED";
    FD1P3AX instr_data_3__i52 (.D(instr_data[3]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i52.GSR = "DISABLED";
    FD1P3AX instr_data_3__i51 (.D(instr_data[2]), .SP(clk_c_enable_115), 
            .CK(clk_c), .Q(n5[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i51.GSR = "DISABLED";
    FD1P3AX instr_data_3__i50 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_117), 
            .CK(clk_c), .Q(n5[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i50.GSR = "DISABLED";
    FD1P3AX instr_data_3__i49 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_117), 
            .CK(clk_c), .Q(n5[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i49.GSR = "DISABLED";
    FD1P3AX instr_data_3__i48 (.D(instr_data[15]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i48.GSR = "DISABLED";
    FD1P3AX instr_data_3__i47 (.D(instr_data[14]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i47.GSR = "DISABLED";
    LUT4 mem_data_from_read_4__bdd_3_lut_24122_then_4_lut (.A(\data_txn_len[0] ), 
         .B(\qspi_data_buf[12] ), .C(instr_data[12]), .D(n27150), .Z(n27396)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B)) */ ;
    defparam mem_data_from_read_4__bdd_3_lut_24122_then_4_lut.init = 16'he4cc;
    FD1P3AX instr_data_3__i46 (.D(instr_data[13]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i46.GSR = "DISABLED";
    FD1P3AX instr_data_3__i45 (.D(instr_data[12]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i45.GSR = "DISABLED";
    FD1P3AX instr_data_3__i44 (.D(instr_data[11]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i44.GSR = "DISABLED";
    FD1P3AX instr_data_3__i43 (.D(instr_data[10]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i43.GSR = "DISABLED";
    FD1P3AX instr_data_3__i42 (.D(instr_data[9]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i42.GSR = "DISABLED";
    FD1P3AX instr_data_3__i41 (.D(instr_data[8]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i41.GSR = "DISABLED";
    FD1P3AX instr_data_3__i40 (.D(instr_data[7]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i40.GSR = "DISABLED";
    FD1P3AX instr_data_3__i39 (.D(instr_data[6]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i39.GSR = "DISABLED";
    FD1P3AX instr_data_3__i38 (.D(instr_data[5]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i38.GSR = "DISABLED";
    FD1P3AX instr_data_3__i37 (.D(instr_data[4]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i37.GSR = "DISABLED";
    FD1P3AX instr_data_3__i36 (.D(instr_data[3]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i36.GSR = "DISABLED";
    LUT4 mem_data_from_read_4__bdd_3_lut_24122_else_4_lut (.A(\data_txn_len[0] ), 
         .B(n27150), .C(instr_data[8]), .D(\qspi_data_buf[8] ), .Z(n27395)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mem_data_from_read_4__bdd_3_lut_24122_else_4_lut.init = 16'hf780;
    PFUMX i24165 (.BLUT(n26807), .ALUT(n26806), .C0(n28564), .Z(n19));
    LUT4 mem_data_from_read_6__bdd_3_lut_24109_then_4_lut (.A(\data_txn_len[0] ), 
         .B(\qspi_data_buf[14] ), .C(instr_data[14]), .D(n27150), .Z(n27400)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B)) */ ;
    defparam mem_data_from_read_6__bdd_3_lut_24109_then_4_lut.init = 16'he4cc;
    LUT4 i1_4_lut_rep_470_4_lut (.A(n27109), .B(n23506), .C(n27096), .D(n10_c), 
         .Z(n27095)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_rep_470_4_lut.init = 16'h4000;
    PFUMX i24163 (.BLUT(n26804), .ALUT(n26803), .C0(n27212), .Z(n26805));
    LUT4 mem_data_from_read_6__bdd_3_lut_24109_else_4_lut (.A(\data_txn_len[0] ), 
         .B(n27150), .C(instr_data[10]), .D(\qspi_data_buf[10] ), .Z(n27399)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mem_data_from_read_6__bdd_3_lut_24109_else_4_lut.init = 16'hf780;
    LUT4 instr_27__bdd_4_lut (.A(instr[27]), .B(n27131), .C(n4075), .D(n4703[27]), 
         .Z(n26263)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam instr_27__bdd_4_lut.init = 16'hef20;
    LUT4 mux_1083_i16_3_lut_then_3_lut (.A(n5[15]), .B(n1[15]), .C(n2055), 
         .Z(n27403)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i16_3_lut_then_3_lut.init = 16'hacac;
    LUT4 mux_1083_i16_3_lut_else_3_lut (.A(n31[15]), .B(n33[15]), .C(n2035), 
         .Z(n27402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i16_3_lut_else_3_lut.init = 16'hcaca;
    FD1P3AX imm_i0_i31 (.D(n3350[24]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(imm[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i31.GSR = "DISABLED";
    FD1P3AX imm_i0_i30 (.D(n26304), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(imm[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i30.GSR = "DISABLED";
    FD1P3AX imm_i0_i29 (.D(n3438[29]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(imm[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i29.GSR = "DISABLED";
    FD1P3AX imm_i0_i28 (.D(n3438[28]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(imm[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i28.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut (.A(n27109), .B(n23608), .C(n6), .D(n27103), 
         .Z(n23614)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h4000;
    FD1P3AX imm_i0_i27 (.D(n26264), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(imm[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i27.GSR = "DISABLED";
    FD1P3AX imm_i0_i26 (.D(n3438[26]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(imm[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i26.GSR = "DISABLED";
    LUT4 i23696_3_lut (.A(n4075), .B(n27099), .C(n27260), .Z(n24998)) /* synthesis lut_function=(A+!((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23696_3_lut.init = 16'haeae;
    FD1P3AX imm_i0_i25 (.D(n3438[25]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(imm[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i25.GSR = "DISABLED";
    FD1P3AX imm_i0_i24 (.D(n3438[24]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(imm[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i24.GSR = "DISABLED";
    FD1P3IX is_alu_reg_397 (.D(is_alu_reg_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_alu_reg)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_alu_reg_397.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_adj_316 (.A(n27109), .B(n23618), .C(n6), .D(n27103), 
         .Z(n23624)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_316.init = 16'h4000;
    FD1P3AX imm_i0_i23 (.D(n3438[23]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i23.GSR = "DISABLED";
    FD1P3AX instr_data_3__i35 (.D(instr_data[2]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(n31[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i35.GSR = "DISABLED";
    FD1P3AX instr_data_3__i34 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_144), 
            .CK(clk_c), .Q(n31[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i34.GSR = "DISABLED";
    FD1P3AX instr_data_3__i33 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_144), 
            .CK(clk_c), .Q(n31[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i33.GSR = "DISABLED";
    FD1P3AX instr_data_3__i32 (.D(instr_data[15]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i32.GSR = "DISABLED";
    FD1P3AX instr_data_3__i31 (.D(instr_data[14]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i31.GSR = "DISABLED";
    FD1P3AX instr_data_3__i30 (.D(instr_data[13]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i30.GSR = "DISABLED";
    FD1P3AX instr_data_3__i29 (.D(instr_data[12]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i29.GSR = "DISABLED";
    FD1P3AX instr_data_3__i28 (.D(instr_data[11]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i28.GSR = "DISABLED";
    FD1P3AX instr_data_3__i27 (.D(instr_data[10]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i27.GSR = "DISABLED";
    FD1P3AX instr_data_3__i26 (.D(instr_data[9]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i26.GSR = "DISABLED";
    FD1P3AX instr_data_3__i25 (.D(instr_data[8]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i25.GSR = "DISABLED";
    FD1P3AX instr_data_3__i24 (.D(instr_data[7]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i24.GSR = "DISABLED";
    FD1P3AX instr_data_3__i23 (.D(instr_data[6]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i23.GSR = "DISABLED";
    FD1P3AX instr_data_3__i22 (.D(instr_data[5]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i22.GSR = "DISABLED";
    FD1P3AX instr_data_3__i21 (.D(instr_data[4]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i21.GSR = "DISABLED";
    FD1P3AX instr_data_3__i20 (.D(instr_data[3]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i20.GSR = "DISABLED";
    FD1P3AX instr_data_3__i19 (.D(instr_data[2]), .SP(clk_c_enable_158), 
            .CK(clk_c), .Q(n33[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i19.GSR = "DISABLED";
    FD1P3AX instr_data_3__i18 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_160), 
            .CK(clk_c), .Q(n33[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i18.GSR = "DISABLED";
    FD1P3AX instr_data_3__i17 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_160), 
            .CK(clk_c), .Q(n33[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i17.GSR = "DISABLED";
    FD1P3AX instr_data_3__i16 (.D(instr_data[15]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i16.GSR = "DISABLED";
    FD1P3AX instr_data_3__i15 (.D(instr_data[14]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i15.GSR = "DISABLED";
    FD1P3AX instr_data_3__i14 (.D(instr_data[13]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i14.GSR = "DISABLED";
    FD1P3AX instr_data_3__i13 (.D(instr_data[12]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i13.GSR = "DISABLED";
    FD1P3AX instr_data_3__i12 (.D(instr_data[11]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i12.GSR = "DISABLED";
    FD1P3AX instr_data_3__i11 (.D(instr_data[10]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i11.GSR = "DISABLED";
    FD1P3AX instr_data_3__i10 (.D(instr_data[9]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i10.GSR = "DISABLED";
    FD1P3AX instr_data_3__i9 (.D(instr_data[8]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i9.GSR = "DISABLED";
    FD1P3AX instr_data_3__i8 (.D(instr_data[7]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i8.GSR = "DISABLED";
    FD1P3AX instr_data_3__i7 (.D(instr_data[6]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i7.GSR = "DISABLED";
    FD1P3AX instr_data_3__i6 (.D(instr_data[5]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i6.GSR = "DISABLED";
    FD1P3AX instr_data_3__i5 (.D(instr_data[4]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i5.GSR = "DISABLED";
    FD1P3AX instr_data_3__i4 (.D(instr_data[3]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i4.GSR = "DISABLED";
    FD1P3AX instr_data_3__i3 (.D(instr_data[2]), .SP(clk_c_enable_174), 
            .CK(clk_c), .Q(n1[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i3.GSR = "DISABLED";
    FD1P3AX instr_data_3__i2 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_175), 
            .CK(clk_c), .Q(n1[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i2.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i2 (.D(additional_mem_ops_2__N_749[2]), .CK(clk_c), 
            .CD(n27326), .Q(additional_mem_ops[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i2.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i1 (.D(additional_mem_ops_2__N_749[1]), .CK(clk_c), 
            .CD(n27326), .Q(additional_mem_ops[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i1.GSR = "DISABLED";
    LUT4 n26279_bdd_3_lut (.A(n26277), .B(instr[31]), .C(n4057), .Z(n26280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26279_bdd_3_lut.init = 16'hcaca;
    PFUMX i24159 (.BLUT(n26794), .ALUT(n26793), .C0(n27298), .Z(n26795));
    LUT4 i1_4_lut_4_lut_adj_317 (.A(n27109), .B(n23628), .C(n6), .D(n27103), 
         .Z(n23634)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_317.init = 16'h4000;
    LUT4 n1750_bdd_3_lut (.A(n1735[1]), .B(n27260), .C(n24666), .Z(n26277)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n1750_bdd_3_lut.init = 16'hb8b8;
    FD1P3AX imm_i0_i22 (.D(n3438[22]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i22.GSR = "DISABLED";
    FD1P3IX is_auipc_395 (.D(is_auipc_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_auipc)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_auipc_395.GSR = "DISABLED";
    LUT4 n3412_bdd_3_lut_23867 (.A(n3397[17]), .B(n26282), .C(n4079), 
         .Z(n26283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3412_bdd_3_lut_23867.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n27330), .B(imm[0]), .C(\imm[1] ), .D(\imm[10] ), 
         .Z(n24360)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i3_rep_476_4_lut (.A(n27109), .B(n27106), .C(n23498), .D(n27123), 
         .Z(n27101)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_rep_476_4_lut.init = 16'h4000;
    FD1P3AX instr_fetch_running_429 (.D(n5590), .SP(clk_c_enable_209), .CK(clk_c), 
            .Q(instr_fetch_running)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_fetch_running_429.GSR = "DISABLED";
    LUT4 n26291_bdd_3_lut (.A(n26289), .B(instr[31]), .C(n4057), .Z(n26292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26291_bdd_3_lut.init = 16'hcaca;
    LUT4 i23702_2_lut_rep_460 (.A(n4073), .B(n4065), .Z(n27085)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23702_2_lut_rep_460.init = 16'hbbbb;
    FD1P3AX imm_i0_i21 (.D(n3438[21]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i21.GSR = "DISABLED";
    FD1P3IX is_system_402 (.D(is_system_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_system)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_system_402.GSR = "DISABLED";
    FD1P3AX imm_i0_i20 (.D(n3438[20]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i20.GSR = "DISABLED";
    LUT4 i23390_3_lut_4_lut (.A(n4073), .B(n4065), .C(n3163[8]), .D(n2874[8]), 
         .Z(n3314[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23390_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_622_4_lut (.A(n27374), .B(n27287), .C(n24360), .D(\imm[6] ), 
         .Z(n27247)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_2_lut_rep_622_4_lut.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_318 (.A(n27109), .B(rst_reg_n), .C(n27), .D(n27103), 
         .Z(n2700)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_318.init = 16'h4000;
    FD1P3AX imm_i0_i19 (.D(n26300), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i19.GSR = "DISABLED";
    FD1P3AX imm_i0_i18 (.D(n26295), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i18.GSR = "DISABLED";
    FD1P3AX imm_i0_i17 (.D(n26283), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[17] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i17.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_319 (.A(n8900), .B(n22088), .C(n24160), .D(n22178), 
         .Z(n22090)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_4_lut_adj_319.init = 16'hc888;
    LUT4 i1_4_lut_4_lut_adj_320 (.A(n27109), .B(n23544), .C(n16), .D(n27103), 
         .Z(n2029)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_320.init = 16'h4000;
    LUT4 mux_1077_i12_3_lut (.A(n1[11]), .B(n5[11]), .C(n2055), .Z(n1735[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1073_i12_3_lut (.A(n31[11]), .B(n33[11]), .C(n2035), .Z(n1715[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i12_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_321 (.A(n27109), .B(n28575), .C(n27096), .D(n10_c), 
         .Z(n22534)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_321.init = 16'h4000;
    LUT4 mux_1956_i10_3_lut_4_lut (.A(n4073), .B(n4065), .C(n3163[9]), 
         .D(n2874[9]), .Z(n3314[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1956_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i23703_2_lut_3_lut_4_lut (.A(n4073), .B(n4065), .C(n4079), .D(n27086), 
         .Z(n24976)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23703_2_lut_3_lut_4_lut.init = 16'hf4f0;
    FD1P3AX data_write_n_i1 (.D(data_write_n_1__N_369[1]), .SP(clk_c_enable_278), 
            .CK(clk_c), .Q(qv_data_write_n[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_write_n_i1.GSR = "DISABLED";
    FD1P3AX imm_i0_i16 (.D(n3438[16]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[16] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i16.GSR = "DISABLED";
    FD1P3AX imm_i0_i15 (.D(n3438[15]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[15] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i15.GSR = "DISABLED";
    FD1P3AX imm_i0_i14 (.D(n3438[14]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[14] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i14.GSR = "DISABLED";
    FD1P3AX imm_i0_i13 (.D(n3438[13]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[13] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i13.GSR = "DISABLED";
    FD1P3AX imm_i0_i12 (.D(n3438[12]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[12] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i12.GSR = "DISABLED";
    FD1P3AX imm_i0_i11 (.D(n3438[11]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[11] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i11.GSR = "DISABLED";
    FD1P3IX is_lui_398 (.D(is_lui_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_lui)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_lui_398.GSR = "DISABLED";
    FD1P3IX is_store_396 (.D(is_store_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_store)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_store_396.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_adj_322 (.A(n27109), .B(n23638), .C(n6), .D(n27103), 
         .Z(n23644)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_322.init = 16'h4000;
    FD1P3AX imm_i0_i10 (.D(n3438[10]), .SP(clk_c_enable_227), .CK(clk_c), 
            .Q(\imm[10] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i10.GSR = "DISABLED";
    LUT4 mux_1077_i4_3_lut (.A(n1[3]), .B(n5[3]), .C(n2055), .Z(n1735[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1073_i4_3_lut (.A(n31[3]), .B(n33[3]), .C(n2035), .Z(n1715[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1077_i9_3_lut (.A(n1[8]), .B(n5[8]), .C(n2055), .Z(n1735[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1073_i9_3_lut (.A(n31[8]), .B(n33[8]), .C(n2035), .Z(n1715[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i9_3_lut.init = 16'hcaca;
    FD1P3AX imm_i0_i9 (.D(n3438[9]), .SP(clk_c_enable_229), .CK(clk_c), 
            .Q(\imm[9] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i9.GSR = "DISABLED";
    FD1P3AX imm_i0_i8 (.D(n3438[8]), .SP(clk_c_enable_229), .CK(clk_c), 
            .Q(\imm[8] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i8.GSR = "DISABLED";
    LUT4 mux_1077_i10_3_lut (.A(n1[9]), .B(n5[9]), .C(n2055), .Z(n1735[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1073_i10_3_lut (.A(n31[9]), .B(n33[9]), .C(n2035), .Z(n1715[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1077_i13_3_lut (.A(n1[12]), .B(n5[12]), .C(n2055), .Z(n1735[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1073_i13_3_lut (.A(n31[12]), .B(n33[12]), .C(n2035), .Z(n1715[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1077_i14_3_lut (.A(n1[13]), .B(n5[13]), .C(n2055), .Z(n1735[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1073_i14_3_lut (.A(n31[13]), .B(n33[13]), .C(n2035), .Z(n1715[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i14_3_lut.init = 16'hcaca;
    LUT4 i12432_2_lut_rep_471_3_lut_4_lut (.A(n27108), .B(n27114), .C(n27109), 
         .D(n23682), .Z(n27096)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i12432_2_lut_rep_471_3_lut_4_lut.init = 16'hf0fe;
    FD1P3JX no_write_in_progress_419 (.D(no_write_in_progress_N_471), .SP(clk_c_enable_231), 
            .PD(n27326), .CK(clk_c), .Q(no_write_in_progress)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam no_write_in_progress_419.GSR = "DISABLED";
    FD1P3IX is_branch_399 (.D(is_branch_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_branch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_branch_399.GSR = "DISABLED";
    LUT4 n1749_bdd_3_lut (.A(n1735[2]), .B(n27260), .C(n24668), .Z(n26289)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n1749_bdd_3_lut.init = 16'hb8b8;
    FD1P3AX rs2_i0_i0 (.D(n1815[0]), .SP(clk_c_enable_372), .CK(clk_c), 
            .Q(rs2[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i0.GSR = "DISABLED";
    FD1P3AX imm_i0_i7 (.D(n3438[7]), .SP(clk_c_enable_245), .CK(clk_c), 
            .Q(\imm[7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i7.GSR = "DISABLED";
    FD1P3AX imm_i0_i6 (.D(n3438[6]), .SP(clk_c_enable_245), .CK(clk_c), 
            .Q(\imm[6] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i6.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n27108), .B(n27114), .C(n22885), .D(n23682), 
         .Z(clk_c_enable_242)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i440_2_lut_rep_473_3_lut_4_lut (.A(n27108), .B(n27114), .C(n27109), 
         .D(n23682), .Z(clk_c_enable_34)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i440_2_lut_rep_473_3_lut_4_lut.init = 16'h000e;
    LUT4 n3412_bdd_3_lut_23872 (.A(n3397[17]), .B(n26294), .C(n4079), 
         .Z(n26295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3412_bdd_3_lut_23872.init = 16'hcaca;
    LUT4 i1_3_lut_rep_477_4_lut (.A(n27108), .B(n27114), .C(n23682), .D(n27109), 
         .Z(n27102)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i1_3_lut_rep_477_4_lut.init = 16'hfff1;
    FD1P3AX imm_i0_i5 (.D(n3438[5]), .SP(clk_c_enable_245), .CK(clk_c), 
            .Q(\imm[5] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i5.GSR = "DISABLED";
    FD1P3AX imm_i0_i4 (.D(n3438[4]), .SP(clk_c_enable_245), .CK(clk_c), 
            .Q(\imm[4] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i4.GSR = "DISABLED";
    FD1P3IX is_load_393 (.D(is_load_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_load)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_load_393.GSR = "DISABLED";
    LUT4 mux_1975_i12_3_lut_4_lut (.A(n27086), .B(n27085), .C(n3314[11]), 
         .D(n2874[9]), .Z(n3397[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1975_i12_3_lut_4_lut.init = 16'hf2d0;
    FD1P3IX is_jal_401 (.D(is_jal_de), .SP(clk_c_enable_242), .CD(n27326), 
            .CK(clk_c), .Q(is_jal)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_jal_401.GSR = "DISABLED";
    LUT4 i22856_3_lut (.A(imm[27]), .B(imm[31]), .C(counter_hi[2]), .Z(n25199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22856_3_lut.init = 16'hcaca;
    LUT4 i22855_3_lut (.A(\imm[19] ), .B(\imm[23] ), .C(counter_hi[2]), 
         .Z(n25198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22855_3_lut.init = 16'hcaca;
    LUT4 i22854_3_lut (.A(\imm[11] ), .B(\imm[15] ), .C(counter_hi[2]), 
         .Z(n25197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22854_3_lut.init = 16'hcaca;
    LUT4 i22853_3_lut (.A(\imm[3] ), .B(\imm[7] ), .C(counter_hi[2]), 
         .Z(n25196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22853_3_lut.init = 16'hcaca;
    FD1P3AX imm_i0_i3 (.D(n3438[3]), .SP(clk_c_enable_245), .CK(clk_c), 
            .Q(\imm[3] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i3.GSR = "DISABLED";
    FD1P3AX imm_i0_i2 (.D(n26119), .SP(clk_c_enable_245), .CK(clk_c), 
            .Q(\imm[2] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i2.GSR = "DISABLED";
    LUT4 n4069_bdd_3_lut_24230 (.A(n4057), .B(instr[31]), .C(instr[19]), 
         .Z(n26297)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n4069_bdd_3_lut_24230.init = 16'hd8d8;
    LUT4 i22849_3_lut (.A(imm[26]), .B(imm[30]), .C(counter_hi[2]), .Z(n25192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22849_3_lut.init = 16'hcaca;
    FD1P3AX imm_i0_i1 (.D(n3438[1]), .SP(clk_c_enable_245), .CK(clk_c), 
            .Q(\imm[1] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i1.GSR = "DISABLED";
    LUT4 i22848_3_lut (.A(\imm[18] ), .B(\imm[22] ), .C(counter_hi[2]), 
         .Z(n25191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22848_3_lut.init = 16'hcaca;
    PFUMX i23813 (.BLUT(n26202), .ALUT(n26201), .C0(counter_hi[2]), .Z(n26203));
    LUT4 debug_branch_I_48_i4_3_lut (.A(debug_branch_N_840[31]), .B(timer_data[3]), 
         .C(is_timer_addr), .Z(debug_branch_N_450[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_48_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_323 (.A(n23980), .B(n23087), .C(n27289), .D(n27354), 
         .Z(n12)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !((C (D)+!C !(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[82:120])
    defparam i1_4_lut_adj_323.init = 16'h8448;
    LUT4 stall_core_I_0_438_2_lut_rep_663 (.A(stall_core), .B(interrupt_core), 
         .Z(n27288)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(340[19:48])
    defparam stall_core_I_0_438_2_lut_rep_663.init = 16'h2222;
    LUT4 i12481_2_lut_3_lut (.A(stall_core), .B(interrupt_core), .C(n27342), 
         .Z(n14783)) /* synthesis lut_function=(!(A (B (C))+!A (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(340[19:48])
    defparam i12481_2_lut_3_lut.init = 16'h2f2f;
    LUT4 i22847_3_lut (.A(\imm[10] ), .B(\imm[14] ), .C(counter_hi[2]), 
         .Z(n25190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22847_3_lut.init = 16'hcaca;
    LUT4 i22846_3_lut (.A(\imm[2] ), .B(\imm[6] ), .C(counter_hi[2]), 
         .Z(n25189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22846_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_324 (.A(clk_c_enable_372), .B(n27109), .C(n23838), 
         .D(n27106), .Z(n2704)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_324.init = 16'ha888;
    FD1P3IX data_addr__i27 (.D(addr_out[27]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i27.GSR = "DISABLED";
    LUT4 i22842_3_lut (.A(imm[25]), .B(imm[29]), .C(counter_hi[2]), .Z(n25185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22842_3_lut.init = 16'hcaca;
    FD1P3IX data_addr__i26 (.D(addr_out[26]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i26.GSR = "DISABLED";
    FD1P3IX data_addr__i25 (.D(addr_out[25]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i25.GSR = "DISABLED";
    FD1P3IX data_addr__i24 (.D(addr_out[24]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i24.GSR = "DISABLED";
    FD1P3IX data_addr__i23 (.D(addr_out[23]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[23])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i23.GSR = "DISABLED";
    FD1P3IX data_addr__i22 (.D(addr_out[22]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[22])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i22.GSR = "DISABLED";
    FD1P3IX data_addr__i21 (.D(addr_out[21]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[21])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i21.GSR = "DISABLED";
    FD1P3IX data_addr__i20 (.D(addr_out[20]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[20])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i20.GSR = "DISABLED";
    FD1P3IX data_addr__i19 (.D(addr_out[19]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[19])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i19.GSR = "DISABLED";
    FD1P3IX data_addr__i18 (.D(addr_out[18]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[18])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i18.GSR = "DISABLED";
    FD1P3IX data_addr__i17 (.D(addr_out[17]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[17])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i17.GSR = "DISABLED";
    PFUMX i24125 (.BLUT(n26732), .ALUT(n26728), .C0(n27298), .Z(n26733));
    FD1P3IX data_addr__i16 (.D(addr_out[16]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[16])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i16.GSR = "DISABLED";
    FD1P3IX data_addr__i15 (.D(addr_out[15]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i15.GSR = "DISABLED";
    FD1P3IX data_addr__i14 (.D(addr_out[14]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i14.GSR = "DISABLED";
    FD1P3IX data_addr__i13 (.D(addr_out[13]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i13.GSR = "DISABLED";
    FD1P3IX data_addr__i12 (.D(addr_out[12]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i12.GSR = "DISABLED";
    FD1P3IX data_addr__i11 (.D(addr_out[11]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i11.GSR = "DISABLED";
    FD1P3IX data_addr__i10 (.D(addr_out[10]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i10.GSR = "DISABLED";
    FD1P3IX data_addr__i9 (.D(addr_out[9]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i9.GSR = "DISABLED";
    FD1P3IX data_addr__i8 (.D(addr_out[8]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i8.GSR = "DISABLED";
    FD1P3IX data_addr__i7 (.D(addr_out[7]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i7.GSR = "DISABLED";
    FD1P3IX data_addr__i6 (.D(addr_out[6]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i6.GSR = "DISABLED";
    FD1P3IX data_addr__i5 (.D(addr_out[5]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i5.GSR = "DISABLED";
    FD1P3IX data_addr__i4 (.D(addr_out[4]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i4.GSR = "DISABLED";
    FD1P3IX data_addr__i3 (.D(n23045), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i3.GSR = "DISABLED";
    FD1P3IX data_addr__i2 (.D(n699[0]), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i2.GSR = "DISABLED";
    FD1P3IX data_addr__i1 (.D(\addr_out[1] ), .SP(clk_c_enable_272), .CD(n27326), 
            .CK(clk_c), .Q(addr[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i1.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i3 (.D(\next_instr_write_offset[3] ), .CK(clk_c), 
            .CD(n22226), .Q(\instr_write_offset[3] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i3.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i2 (.D(instr_write_offset_3__N_934[1]), .CK(clk_c), 
            .CD(n27326), .Q(instr_addr_23__N_318[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i2.GSR = "DISABLED";
    LUT4 n3412_bdd_3_lut_23874 (.A(n3397[17]), .B(n26299), .C(n4079), 
         .Z(n26300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3412_bdd_3_lut_23874.init = 16'hcaca;
    LUT4 i4019_3_lut_4_lut (.A(\instr_addr_23__N_318[0] ), .B(n27355), .C(n27297), 
         .D(instr_addr_23__N_318[1]), .Z(n4)) /* synthesis lut_function=(A ((D)+!C)+!A !(B (C+!(D))+!B !((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i4019_3_lut_4_lut.init = 16'hbf0b;
    LUT4 i22841_3_lut (.A(\imm[17] ), .B(\imm[21] ), .C(counter_hi[2]), 
         .Z(n25184)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22841_3_lut.init = 16'hcaca;
    LUT4 i22840_3_lut (.A(\imm[9] ), .B(\imm[13] ), .C(counter_hi[2]), 
         .Z(n25183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22840_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_325 (.A(\instr_write_offset[3] ), .B(instr_addr_23__N_318[1]), 
         .C(\pc[2] ), .D(n2), .Z(n9)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A !(B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam i1_4_lut_4_lut_adj_325.init = 16'h4124;
    PFUMX i24123 (.BLUT(n26730), .ALUT(\mem_data_from_read[4] ), .C0(counter_hi[2]), 
          .Z(n26731));
    LUT4 i1_4_lut_adj_326 (.A(n23398), .B(n23402), .C(instr_complete_N_1647), 
         .D(stall_core), .Z(\next_instr_write_offset[3] )) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i1_4_lut_adj_326.init = 16'haa6a;
    LUT4 i22839_3_lut (.A(\imm[1] ), .B(\imm[5] ), .C(counter_hi[2]), 
         .Z(n25182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22839_3_lut.init = 16'hcaca;
    LUT4 i22835_3_lut (.A(imm[24]), .B(imm[28]), .C(counter_hi[2]), .Z(n25178)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22835_3_lut.init = 16'hcaca;
    LUT4 i22834_3_lut (.A(\imm[16] ), .B(\imm[20] ), .C(counter_hi[2]), 
         .Z(n25177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22834_3_lut.init = 16'hcaca;
    LUT4 i22833_3_lut (.A(\imm[8] ), .B(\imm[12] ), .C(counter_hi[2]), 
         .Z(n25176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22833_3_lut.init = 16'hcaca;
    LUT4 i22832_3_lut (.A(imm[0]), .B(\imm[4] ), .C(counter_hi[2]), .Z(n25175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22832_3_lut.init = 16'hcaca;
    LUT4 i23593_3_lut_4_lut (.A(n27347), .B(alu_op[2]), .C(n27302), .D(n15_adj_2637), 
         .Z(n25132)) /* synthesis lut_function=(A (C+!(D))+!A (B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i23593_3_lut_4_lut.init = 16'hf4ff;
    LUT4 n27211_bdd_4_lut_24741 (.A(n27211), .B(n27142), .C(n27212), .D(n28563), 
         .Z(n28140)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D))+!B (C)))) */ ;
    defparam n27211_bdd_4_lut_24741.init = 16'h0fe5;
    FD1P3AX mem_op_increment_reg_413 (.D(n24804), .SP(clk_c_enable_275), 
            .CK(clk_c), .Q(mem_op_increment_reg)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_increment_reg_413.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_482 (.A(address_ready), .B(n27111), .C(is_load), 
         .Z(n27107)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(291[13:39])
    defparam i1_3_lut_rep_482.init = 16'h2020;
    LUT4 n3412_bdd_3_lut (.A(n3397[17]), .B(n26875), .C(n4079), .Z(n26304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3412_bdd_3_lut.init = 16'hcaca;
    LUT4 n27211_bdd_4_lut_24826 (.A(n27212), .B(n2036[0]), .C(n2056[0]), 
         .D(n27260), .Z(n28142)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam n27211_bdd_4_lut_24826.init = 16'h5044;
    LUT4 i12829_3_lut_4_lut (.A(n27148), .B(n28563), .C(n27212), .D(n27211), 
         .Z(n29)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (D)))) */ ;
    defparam i12829_3_lut_4_lut.init = 16'h001f;
    LUT4 i1_2_lut_4_lut (.A(address_ready), .B(n27111), .C(is_load), .D(n27226), 
         .Z(clk_c_enable_53)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(291[13:39])
    defparam i1_2_lut_4_lut.init = 16'hff20;
    PFUMX i23809 (.BLUT(n26197), .ALUT(n26196), .C0(counter_hi[2]), .Z(n26198));
    PFUMX i24112 (.BLUT(n26716), .ALUT(n26712), .C0(n27298), .Z(n26717));
    LUT4 imm_1__bdd_3_lut_24030 (.A(\imm[4] ), .B(\imm[8] ), .C(\imm[9] ), 
         .Z(n26317)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam imm_1__bdd_3_lut_24030.init = 16'h0101;
    LUT4 shift_right_317_i271_3_lut (.A(n24752), .B(load_top_bit), .C(data_out_3__N_1385), 
         .Z(debug_branch_N_840[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam shift_right_317_i271_3_lut.init = 16'hcaca;
    LUT4 mux_1073_i1_rep_121_3_lut (.A(n31[0]), .B(n33[0]), .C(n2035), 
         .Z(n24664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i1_rep_121_3_lut.init = 16'hcaca;
    LUT4 shift_right_317_i269_3_lut (.A(n24746), .B(load_top_bit), .C(data_out_3__N_1385), 
         .Z(debug_branch_N_840[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam shift_right_317_i269_3_lut.init = 16'hcaca;
    LUT4 next_pc_for_core_23__I_0_i271_4_lut (.A(n27023), .B(debug_rd_3__N_405[30]), 
         .C(n27319), .D(n7717), .Z(debug_branch_N_446[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i271_4_lut.init = 16'hcac0;
    LUT4 mux_1083_i1_rep_115_3_lut (.A(n1735[0]), .B(instr[31]), .C(n4057), 
         .Z(n24658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i1_rep_115_3_lut.init = 16'hcaca;
    LUT4 mux_1077_i1_3_lut (.A(n1[0]), .B(n5[0]), .C(n2055), .Z(n1735[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1083_i1_3_lut (.A(n24664), .B(n1735[0]), .C(n27260), .Z(instr[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1077_i6_3_lut (.A(n1[5]), .B(n5[5]), .C(n2055), .Z(n1735[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i6_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(n22898), .B(n27111), .C(n23600), .D(n8), 
         .Z(n22816)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[22:78])
    defparam i1_3_lut_4_lut.init = 16'h00d0;
    LUT4 imm_1__bdd_4_lut_24066 (.A(imm[0]), .B(\imm[4] ), .C(\imm[8] ), 
         .D(\imm[9] ), .Z(n26316)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam imm_1__bdd_4_lut_24066.init = 16'h8001;
    LUT4 csr_read_3__N_1463_1__bdd_3_lut_24239_4_lut (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(cycle_count_wide[4]), .D(time_hi[0]), .Z(n26926)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam csr_read_3__N_1463_1__bdd_3_lut_24239_4_lut.init = 16'hf2d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_327 (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(n22898), .D(n22499), .Z(n23928)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_327.init = 16'h2f0f;
    PFUMX i24110 (.BLUT(n26714), .ALUT(\mem_data_from_read[6] ), .C0(counter_hi[2]), 
          .Z(n26715));
    LUT4 i20149_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(rst_reg_n), .D(n22499), .Z(n22369)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;
    defparam i20149_2_lut_3_lut_4_lut.init = 16'hd0f0;
    FD1P3AX data_write_n_i0 (.D(data_write_n_1__N_369[0]), .SP(clk_c_enable_278), 
            .CK(clk_c), .Q(qv_data_write_n[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_write_n_i0.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_488_4_lut (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(instr_complete_N_1647), .D(stall_core), .Z(n27113)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_3_lut_rep_488_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_478_3_lut_4_lut (.A(n22898), .B(n27111), .C(n23682), 
         .D(n27114), .Z(n27103)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[22:78])
    defparam i1_2_lut_rep_478_3_lut_4_lut.init = 16'h0f0d;
    FD1P3AX data_read_n_i0_i1 (.D(n22866), .SP(clk_c_enable_280), .CK(clk_c), 
            .Q(qv_data_read_n[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_read_n_i0_i1.GSR = "DISABLED";
    FD1P3AX rs1_i0_i3 (.D(n2175[3]), .SP(clk_c_enable_282), .CK(clk_c), 
            .Q(rs1[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i3.GSR = "DISABLED";
    LUT4 debug_branch_N_441_I_0_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(was_early_branch), .D(n22499), .Z(instr_fetch_restart_N_947)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam debug_branch_N_441_I_0_2_lut_3_lut_4_lut.init = 16'hfdff;
    FD1P3AX rs1_i0_i2 (.D(n2175[2]), .SP(clk_c_enable_282), .CK(clk_c), 
            .Q(rs1[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i2.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_328 (.A(n27179), .B(rst_reg_n), .C(n4_adj_2638), 
         .D(n8274), .Z(n23690)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_328.init = 16'h0040;
    LUT4 cycle_count_wide_6__I_0_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(time_hi[2]), .D(cycle_count_wide[6]), .Z(time_count[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam cycle_count_wide_6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_4_lut_adj_329 (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(mstatus_mie), .D(interrupt_pending_N_1671), .Z(n23292)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_329.init = 16'h2000;
    LUT4 i1_2_lut_3_lut (.A(any_additional_mem_ops), .B(n27113), .C(n4116[0]), 
         .Z(additional_mem_ops_2__N_749[0])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(149[27:88])
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 gnd_bdd_2_lut_23906_2_lut_3_lut (.A(any_additional_mem_ops), .B(n27113), 
         .C(n26345), .Z(n26346)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(149[27:88])
    defparam gnd_bdd_2_lut_23906_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_3_lut_4_lut_adj_330 (.A(any_additional_mem_ops), .B(n27113), 
         .C(n4116[0]), .D(n4116[1]), .Z(additional_mem_ops_2__N_749[1])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(149[27:88])
    defparam i1_3_lut_4_lut_adj_330.init = 16'hf708;
    LUT4 next_pc_for_core_23__I_0_i270_4_lut (.A(n26932), .B(debug_rd_3__N_405[29]), 
         .C(n27319), .D(n7717), .Z(debug_branch_N_446[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i270_4_lut.init = 16'hcac0;
    PFUMX i23801 (.BLUT(n26177), .ALUT(n26176), .C0(counter_hi[2]), .Z(n26178));
    LUT4 cycle_count_wide_5__I_0_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(time_hi[1]), .D(cycle_count_wide[5]), .Z(time_count[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam cycle_count_wide_5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 mie_9__bdd_4_lut (.A(mie[9]), .B(counter_hi[3]), .C(mie[1]), 
         .D(counter_hi[4]), .Z(n26336)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B+!(C (D)))) */ ;
    defparam mie_9__bdd_4_lut.init = 16'hb8aa;
    LUT4 next_pc_for_core_23__I_0_i272_4_lut (.A(n5167[3]), .B(debug_rd_3__N_405[31]), 
         .C(n27319), .D(n7717), .Z(debug_branch_N_446[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i272_4_lut.init = 16'hcac0;
    LUT4 mie_9__bdd_4_lut_23894 (.A(mie[5]), .B(mie[13]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n26335)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mie_9__bdd_4_lut_23894.init = 16'hcac0;
    LUT4 i43_3_lut (.A(n27209), .B(n27211), .C(n22080), .Z(n24)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;
    defparam i43_3_lut.init = 16'h6464;
    LUT4 i1_4_lut_adj_331 (.A(n22), .B(n8274), .C(n4_adj_2638), .D(n27151), 
         .Z(n23894)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_331.init = 16'h0002;
    L6MUX21 mux_1984_i1 (.D0(n3397[0]), .D1(n3350[0]), .SD(n4079), .Z(n3438[0]));
    PFUMX mux_1975_i1 (.BLUT(n3273[0]), .ALUT(n24505), .C0(n27086), .Z(n3397[0]));
    FD1S3IX counter_hi_3236__i3 (.D(n34[1]), .CK(clk_c), .CD(n27326), 
            .Q(counter_hi[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3236__i3.GSR = "DISABLED";
    LUT4 mux_1083_i3_3_lut (.A(n24668), .B(n1735[2]), .C(n27260), .Z(instr[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i3_3_lut.init = 16'hcaca;
    L6MUX21 mux_1984_i5 (.D0(n3397[4]), .D1(n3350[4]), .SD(n4079), .Z(n3438[4]));
    PFUMX mux_1984_i21 (.BLUT(n24625), .ALUT(n3350[20]), .C0(n24900), 
          .Z(n3438[20]));
    PFUMX mux_1984_i22 (.BLUT(n24627), .ALUT(n3350[21]), .C0(n24900), 
          .Z(n3438[21]));
    PFUMX mux_1984_i23 (.BLUT(n24635), .ALUT(n3350[22]), .C0(n24900), 
          .Z(n3438[22]));
    LUT4 i1_4_lut_adj_332 (.A(n27163), .B(n27211), .C(n27167), .D(n28575), 
         .Z(n23506)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_332.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_333 (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(n23600), .D(n22499), .Z(n23602)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_333.init = 16'hd0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_334 (.A(counter_hi[2]), .B(clk_c_enable_424), 
         .C(next_pc_offset[3]), .D(any_additional_mem_ops), .Z(n23402)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_334.init = 16'h0020;
    PFUMX mux_1984_i24 (.BLUT(n24633), .ALUT(n3350[23]), .C0(n24900), 
          .Z(n3438[23]));
    LUT4 i1_3_lut_4_lut_adj_335 (.A(n27179), .B(n27163), .C(rst_reg_n), 
         .D(instr[20]), .Z(n23638)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_335.init = 16'hb000;
    LUT4 i1_3_lut_4_lut_adj_336 (.A(n27179), .B(n27163), .C(rst_reg_n), 
         .D(instr[23]), .Z(n23628)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_336.init = 16'hb000;
    PFUMX mux_1984_i27 (.BLUT(n24641), .ALUT(n3350[26]), .C0(n24900), 
          .Z(n3438[26]));
    LUT4 i23192_3_lut (.A(\mem_data_from_read[27] ), .B(\mem_data_from_read[31] ), 
         .C(counter_hi[2]), .Z(n24758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam i23192_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_337 (.A(n27179), .B(n27163), .C(n28575), .D(instr[22]), 
         .Z(n23608)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_337.init = 16'hb000;
    FD1P3IX pc_offset__i23 (.D(pc_23__N_911[20]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[23] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i23.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_338 (.A(n27179), .B(n27163), .C(n28575), .D(instr[21]), 
         .Z(n23618)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_338.init = 16'hb000;
    LUT4 i1_4_lut_adj_339 (.A(n22592), .B(n27097), .C(debug_stop_txn_N_2148), 
         .D(instr_fetch_restart_N_947), .Z(debug_stop_txn_N_2147)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(435[34:115])
    defparam i1_4_lut_adj_339.init = 16'h1000;
    L6MUX21 mux_1975_i6 (.D0(n3273[5]), .D1(n3314[5]), .SD(n27086), .Z(n3397[5]));
    PFUMX mux_1975_i5 (.BLUT(n3273[4]), .ALUT(n3314[4]), .C0(n27086), 
          .Z(n3397[4]));
    FD1S3IX counter_hi_3236__i4 (.D(n34[2]), .CK(clk_c), .CD(n27326), 
            .Q(counter_hi[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3236__i4.GSR = "DISABLED";
    LUT4 i23699_2_lut_3_lut_4_lut (.A(clk_c_enable_282), .B(n27179), .C(n4079), 
         .D(n26), .Z(n24984)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i23699_2_lut_3_lut_4_lut.init = 16'hfdff;
    FD1S3IX addr_offset_3237__i3 (.D(n24509), .CK(clk_c), .CD(n27326), 
            .Q(addr_offset[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam addr_offset_3237__i3.GSR = "DISABLED";
    LUT4 i22432_3_lut_4_lut (.A(n27354), .B(n27353), .C(counter_hi[2]), 
         .D(\next_pc_for_core[6] ), .Z(n24775)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i22432_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_347_i2_3_lut_4_lut (.A(n27354), .B(n27353), .C(debug_ret), 
         .D(return_addr[2]), .Z(n1768[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam mux_347_i2_3_lut_4_lut.init = 16'hf606;
    LUT4 i23199_3_lut (.A(n24747), .B(timer_data[0]), .C(is_timer_addr), 
         .Z(n9111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam i23199_3_lut.init = 16'hcaca;
    L6MUX21 mux_1984_i8 (.D0(n3397[7]), .D1(n3350[7]), .SD(n4079), .Z(n3438[7]));
    LUT4 i1_4_lut_adj_340 (.A(n27190), .B(n27167), .C(n27132), .D(n28563), 
         .Z(is_lui_N_1365)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_340.init = 16'h8000;
    PFUMX mux_1984_i9 (.BLUT(n3314[8]), .ALUT(n3397[8]), .C0(n24984), 
          .Z(n3438[8]));
    LUT4 mux_2857_i9_3_lut (.A(n27212), .B(instr[31]), .C(n4057), .Z(n4745[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2857_i9_3_lut.init = 16'hcaca;
    LUT4 mux_2857_i8_3_lut (.A(n28563), .B(instr[31]), .C(n4057), .Z(n4745[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2857_i8_3_lut.init = 16'hcaca;
    LUT4 i23203_3_lut (.A(n24753), .B(timer_data[2]), .C(is_timer_addr), 
         .Z(n9115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam i23203_3_lut.init = 16'hcaca;
    LUT4 mux_2857_i7_3_lut (.A(n27211), .B(instr[31]), .C(n4057), .Z(n4745[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2857_i7_3_lut.init = 16'hcaca;
    LUT4 mux_2857_i6_3_lut (.A(n27205), .B(instr[31]), .C(n4057), .Z(n4745[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2857_i6_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_341 (.A(n27191), .B(n23462), .C(n27160), .D(n22534), 
         .Z(n22671)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_341.init = 16'h4000;
    PFUMX mux_1984_i10 (.BLUT(n3314[9]), .ALUT(n3397[9]), .C0(n24984), 
          .Z(n3438[9]));
    LUT4 i1_4_lut_4_lut_adj_342 (.A(n27191), .B(n23470), .C(n27160), .D(n22534), 
         .Z(n22667)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_342.init = 16'h4000;
    PFUMX mux_1984_i11 (.BLUT(n3314[10]), .ALUT(n3397[10]), .C0(n24976), 
          .Z(n3438[10]));
    LUT4 i1_4_lut_4_lut_adj_343 (.A(n27191), .B(n23478), .C(n27160), .D(n22534), 
         .Z(n22663)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_343.init = 16'h4000;
    PFUMX mux_1984_i12 (.BLUT(n3397[11]), .ALUT(n3350[11]), .C0(n4079), 
          .Z(n3438[11]));
    PFUMX mux_1984_i13 (.BLUT(n3397[12]), .ALUT(n3350[12]), .C0(n4079), 
          .Z(n3438[12]));
    LUT4 i29_4_lut (.A(n28562), .B(n27189), .C(n27135), .D(n27203), 
         .Z(n16)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)+!B !(C+(D))))) */ ;
    defparam i29_4_lut.init = 16'h3534;
    LUT4 i23648_2_lut_3_lut_4_lut (.A(clk_c_enable_282), .B(n27179), .C(n4073), 
         .D(n26), .Z(n25083)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i23648_2_lut_3_lut_4_lut.init = 16'hfdff;
    LUT4 i23394_3_lut_4_lut (.A(n27203), .B(n27084), .C(n4071), .D(n22745), 
         .Z(n3273[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23394_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_3_lut_4_lut_adj_344 (.A(n27211), .B(n27209), .C(n27198), .D(n28564), 
         .Z(n23522)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_344.init = 16'h0010;
    PFUMX mux_1984_i14 (.BLUT(n3397[13]), .ALUT(n3350[13]), .C0(n4079), 
          .Z(n3438[13]));
    LUT4 i1_3_lut_4_lut_adj_345 (.A(n27211), .B(n27209), .C(n27204), .D(n28564), 
         .Z(n23516)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_345.init = 16'h0010;
    PFUMX mux_1984_i15 (.BLUT(n3397[14]), .ALUT(n3350[14]), .C0(n4079), 
          .Z(n3438[14]));
    PFUMX mux_1984_i16 (.BLUT(n3397[15]), .ALUT(n3350[15]), .C0(n4079), 
          .Z(n3438[15]));
    L6MUX21 mux_1984_i17 (.D0(n3397[16]), .D1(n3350[16]), .SD(n4079), 
            .Z(n3438[16]));
    LUT4 n4057_bdd_3_lut_24136 (.A(n1735[5]), .B(n24631), .C(n27260), 
         .Z(n26432)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n4057_bdd_3_lut_24136.init = 16'hacac;
    LUT4 n26432_bdd_3_lut (.A(n26432), .B(n27202), .C(n4057), .Z(n26433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26432_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_346 (.A(clk_c_enable_372), .B(n27109), .C(n23848), 
         .D(n27106), .Z(n2031)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_346.init = 16'ha888;
    LUT4 i12582_2_lut_3_lut_4_lut (.A(clk_c_enable_282), .B(n27179), .C(n22704), 
         .D(n22_adj_2640), .Z(n3087[1])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i12582_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 is_alu_imm_N_1367_bdd_4_lut_4_lut (.A(n28563), .B(n27211), .C(n27209), 
         .D(n27212), .Z(n26807)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam is_alu_imm_N_1367_bdd_4_lut_4_lut.init = 16'h0040;
    LUT4 n4057_bdd_4_lut_24139 (.A(n27179), .B(n1735[5]), .C(n24631), 
         .D(n27260), .Z(n26434)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n4057_bdd_4_lut_24139.init = 16'h88a0;
    LUT4 i1_4_lut_adj_347 (.A(clk_c_enable_372), .B(n27109), .C(n23656), 
         .D(n27106), .Z(n2702)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_347.init = 16'ha888;
    LUT4 mux_1933_i2_4_lut_4_lut (.A(n28563), .B(n4065), .C(n27212), .D(n27199), 
         .Z(n3163[1])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_1933_i2_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i1_4_lut_4_lut_adj_348 (.A(n28563), .B(n24), .C(n23868), .D(n24030), 
         .Z(n23738)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_4_lut_adj_348.init = 16'hf040;
    LUT4 n25708_bdd_4_lut_24202_4_lut (.A(n28563), .B(n28564), .C(n27211), 
         .D(n27212), .Z(n26856)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam n25708_bdd_4_lut_24202_4_lut.init = 16'h0010;
    LUT4 mux_1073_i6_rep_88_3_lut (.A(n31[5]), .B(n33[5]), .C(n2035), 
         .Z(n24631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i6_rep_88_3_lut.init = 16'hcaca;
    LUT4 i12318_2_lut (.A(\next_pc_for_core[4] ), .B(counter_hi[2]), .Z(n149)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i12318_2_lut.init = 16'h8888;
    LUT4 mux_1083_i5_3_lut (.A(n24629), .B(n1735[4]), .C(n27260), .Z(instr[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1083_i11_3_lut (.A(n24642), .B(n1735[10]), .C(n27260), .Z(instr[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i11_3_lut.init = 16'hcaca;
    LUT4 n3193_bdd_4_lut_23762 (.A(n3163[2]), .B(n4073), .C(n28563), .D(n27200), 
         .Z(n26116)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B (C (D)))) */ ;
    defparam n3193_bdd_4_lut_23762.init = 16'he222;
    LUT4 mux_1933_i3_4_lut_4_lut (.A(n28563), .B(n4065), .C(n27212), .D(n27200), 
         .Z(n3163[2])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_1933_i3_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i22430_3_lut (.A(\next_pc_for_core[9] ), .B(\next_pc_for_core[13] ), 
         .C(counter_hi[2]), .Z(n24773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22430_3_lut.init = 16'hcaca;
    LUT4 i7265_2_lut_rep_459_3_lut_4_lut (.A(clk_c_enable_282), .B(n27179), 
         .C(n22704), .D(n22_adj_2640), .Z(n27084)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i7265_2_lut_rep_459_3_lut_4_lut.init = 16'hfdff;
    LUT4 mux_1933_i6_4_lut_4_lut (.A(n28563), .B(n4065), .C(n27212), .D(n27201), 
         .Z(n3163[5])) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C+(D))+!B (D))) */ ;
    defparam mux_1933_i6_4_lut_4_lut.init = 16'hddc0;
    LUT4 mux_1933_i4_4_lut_4_lut (.A(n28563), .B(n4065), .C(n27212), .D(n27198), 
         .Z(n3163[3])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_1933_i4_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i12703_2_lut_3_lut_4_lut (.A(n28563), .B(n27211), .C(n27200), 
         .D(n27175), .Z(n15_adj_2641)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12703_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23250_4_lut_4_lut (.A(n27319), .B(n25142), .C(n234[0]), .D(debug_branch_N_446[28]), 
         .Z(debug_rd_3__N_1567[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i23250_4_lut_4_lut.init = 16'hf1e0;
    FD1P3IX pc_offset__i1 (.D(pc_2__N_932[0]), .SP(clk_c_enable_423), .CD(n27326), 
            .CK(clk_c), .Q(\pc[1] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i1.GSR = "DISABLED";
    PFUMX mux_1947_i6 (.BLUT(n3087[5]), .ALUT(n22715), .C0(n4071), .Z(n3273[5]));
    LUT4 i31_4_lut_4_lut (.A(n27212), .B(n28563), .C(n22080), .D(n27211), 
         .Z(n25)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(C+(D))))) */ ;
    defparam i31_4_lut_4_lut.init = 16'h11fc;
    LUT4 mux_1083_i8_3_lut (.A(n24638), .B(n1735[7]), .C(n27260), .Z(instr[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i8_3_lut.init = 16'hcaca;
    LUT4 i23237_3_lut (.A(n24778), .B(n26795), .C(counter_hi[2]), .Z(n24780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam i23237_3_lut.init = 16'hcaca;
    LUT4 i52_4_lut_4_lut (.A(n28564), .B(n27211), .C(n14587), .D(n28563), 
         .Z(n37)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (D)+!B !(C+(D))))) */ ;
    defparam i52_4_lut_4_lut.init = 16'h4403;
    LUT4 i2_rep_50_3_lut_4_lut (.A(n28564), .B(n27211), .C(n22700), .D(n27209), 
         .Z(n22704)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_rep_50_3_lut_4_lut.init = 16'h0010;
    LUT4 mux_1077_i7_3_lut (.A(n1[6]), .B(n5[6]), .C(n2055), .Z(n1735[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1083_i7_3_lut (.A(n24637), .B(n1735[6]), .C(n27260), .Z(instr[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1083_i6_3_lut (.A(n24631), .B(n1735[5]), .C(n27260), .Z(instr[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i6_3_lut.init = 16'hcaca;
    LUT4 next_pc_for_core_23__I_0_i269_4_lut (.A(n209), .B(n5167[0]), .C(n27293), 
         .D(n7717), .Z(debug_branch_N_446[28])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i269_4_lut.init = 16'haca0;
    PFUMX mux_1975_i17 (.BLUT(n3163[16]), .ALUT(n3314[16]), .C0(n24959), 
          .Z(n3397[16]));
    LUT4 debug_branch_I_48_i4_rep_73_3_lut (.A(timer_data[3]), .B(load_top_bit), 
         .C(data_out_3__N_1385), .Z(n24616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_48_i4_rep_73_3_lut.init = 16'hcaca;
    LUT4 i12552_2_lut_rep_515_3_lut (.A(n27209), .B(n28563), .C(n27205), 
         .Z(n27140)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12552_2_lut_rep_515_3_lut.init = 16'h4040;
    LUT4 i1_3_lut_adj_349 (.A(no_write_in_progress), .B(debug_instr_valid), 
         .C(is_store), .Z(debug_rd_3__N_413)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_3_lut_adj_349.init = 16'h8080;
    PFUMX mux_1975_i8 (.BLUT(n3273[7]), .ALUT(n3314[7]), .C0(n27086), 
          .Z(n3397[7]));
    L6MUX21 mux_1975_i7 (.D0(n3273[6]), .D1(n3314[6]), .SD(n27086), .Z(n3397[6]));
    LUT4 i12551_2_lut_3_lut (.A(n27209), .B(n28563), .C(n27199), .Z(n3196[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12551_2_lut_3_lut.init = 16'h4040;
    L6MUX21 mux_1975_i4 (.D0(n3273[3]), .D1(n3314[3]), .SD(n27086), .Z(n3397[3]));
    L6MUX21 mux_1975_i2 (.D0(n3273[1]), .D1(n3314[1]), .SD(n27086), .Z(n3397[1]));
    PFUMX mux_1393_i3 (.BLUT(n22748), .ALUT(n2161[2]), .C0(n2330), .Z(n2175[2]));
    LUT4 mux_1933_i12_4_lut_4_lut_4_lut (.A(n27209), .B(n28563), .C(n4073), 
         .D(n27205), .Z(n3163[11])) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (C (D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1933_i12_4_lut_4_lut_4_lut.init = 16'h4300;
    LUT4 i23708_3_lut_4_lut (.A(n26), .B(n27092), .C(n4065), .D(n4073), 
         .Z(n24959)) /* synthesis lut_function=(!(A (B (C+(D))))) */ ;
    defparam i23708_3_lut_4_lut.init = 16'h777f;
    LUT4 i22896_3_lut (.A(n25237), .B(n26822), .C(counter_hi[4]), .Z(n25239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22896_3_lut.init = 16'hcaca;
    LUT4 mux_1073_i7_rep_94_3_lut (.A(n31[6]), .B(n33[6]), .C(n2035), 
         .Z(n24637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i7_rep_94_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_631_3_lut_4_lut (.A(n27376), .B(counter_hi[2]), .C(n27305), 
         .D(n27332), .Z(n27256)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_2_lut_rep_631_3_lut_4_lut.init = 16'h0010;
    PFUMX mux_1956_i7 (.BLUT(n3163[6]), .ALUT(n3196[6]), .C0(n4073), .Z(n3314[6]));
    LUT4 pc_23__I_0_450_i269_3_lut (.A(n24612), .B(data_rs1[0]), .C(alu_a_in_3__N_1552), 
         .Z(debug_branch_N_442[28])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam pc_23__I_0_450_i269_3_lut.init = 16'hacac;
    LUT4 i4078_2_lut_rep_603_3_lut_3_lut_4_lut (.A(n27376), .B(counter_hi[2]), 
         .C(cy), .D(cycle_count_wide[0]), .Z(n27228)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i4078_2_lut_rep_603_3_lut_3_lut_4_lut.init = 16'hf100;
    LUT4 cy_I_0_3_lut_rep_621_3_lut_4_lut (.A(n27376), .B(counter_hi[2]), 
         .C(cy_adj_2642), .D(instr_retired), .Z(n27246)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam cy_I_0_3_lut_rep_621_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_350 (.A(n27111), .B(n22885), .C(n27112), .D(n23928), 
         .Z(clk_c_enable_90)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;
    defparam i1_4_lut_adj_350.init = 16'h3332;
    LUT4 pc_23__I_0_450_i157_3_lut (.A(\pc[8] ), .B(\pc[12] ), .C(counter_hi[2]), 
         .Z(n157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam pc_23__I_0_450_i157_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_351 (.A(clk_c_enable_34), .B(n28575), 
         .C(n35), .D(n27179), .Z(n4071)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i1_2_lut_3_lut_4_lut_adj_351.init = 16'h0080;
    LUT4 i1_3_lut_rep_503_4_lut (.A(n27212), .B(n27211), .C(n28563), .D(n27142), 
         .Z(n27128)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_3_lut_rep_503_4_lut.init = 16'h0002;
    LUT4 mux_1956_i19_3_lut_3_lut_4_lut (.A(n26), .B(n27092), .C(n27140), 
         .D(n3273[10]), .Z(n3314[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1956_i19_3_lut_3_lut_4_lut.init = 16'hf780;
    PFUMX i23726 (.BLUT(n26028), .ALUT(n26027), .C0(n4063), .Z(n26029));
    LUT4 i4076_2_lut_3_lut_3_lut_4_lut (.A(n27376), .B(counter_hi[2]), .C(cy), 
         .D(cycle_count_wide[0]), .Z(increment_result_3__N_1911[0])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i4076_2_lut_3_lut_3_lut_4_lut.init = 16'h0ef1;
    LUT4 i1_3_lut_adj_352 (.A(any_additional_mem_ops), .B(n27113), .C(n28575), 
         .Z(n22885)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(149[27:88])
    defparam i1_3_lut_adj_352.init = 16'h8080;
    LUT4 data_ready_sync_I_0_3_lut_3_lut_4_lut (.A(n27376), .B(counter_hi[2]), 
         .C(data_ready_sync), .D(n27124), .Z(data_ready_core)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam data_ready_sync_I_0_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_461_3_lut_4_lut (.A(clk_c_enable_34), .B(n28575), 
         .C(n26), .D(n27179), .Z(n27086)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i1_2_lut_rep_461_3_lut_4_lut.init = 16'h0080;
    LUT4 mux_345_i1_3_lut (.A(\next_pc_for_core[3] ), .B(return_addr[3]), 
         .C(debug_ret), .Z(n36[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i1_3_lut.init = 16'hcaca;
    LUT4 csr_read_3__N_1463_1__bdd_3_lut_24281_3_lut_4_lut (.A(n27376), .B(counter_hi[2]), 
         .C(cycle_count_wide[3]), .D(\imm[1] ), .Z(n26976)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam csr_read_3__N_1463_1__bdd_3_lut_24281_3_lut_4_lut.init = 16'h11f0;
    PFUMX mux_1956_i6 (.BLUT(n3163[5]), .ALUT(n3196[5]), .C0(n4073), .Z(n3314[5]));
    LUT4 mux_1096_i1_4_lut (.A(n27201), .B(rs2[0]), .C(n27109), .D(mem_op_increment_reg), 
         .Z(n1794[0])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1096_i1_4_lut.init = 16'h3aca;
    LUT4 mux_345_i2_3_lut (.A(\next_pc_for_core[4] ), .B(return_addr[4]), 
         .C(debug_ret), .Z(n36[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i2_3_lut.init = 16'hcaca;
    LUT4 mux_345_i3_3_lut (.A(\next_pc_for_core[5] ), .B(return_addr[5]), 
         .C(debug_ret), .Z(n36[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i3_3_lut.init = 16'hcaca;
    LUT4 csr_read_3__N_1463_1__bdd_3_lut_24280_3_lut_4_lut (.A(n27376), .B(counter_hi[2]), 
         .C(mcause[1]), .D(\imm[1] ), .Z(n26930)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam csr_read_3__N_1463_1__bdd_3_lut_24280_3_lut_4_lut.init = 16'h1000;
    LUT4 i12299_2_lut (.A(\pc[4] ), .B(counter_hi[2]), .Z(n149_adj_2643)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam i12299_2_lut.init = 16'h8888;
    LUT4 mux_345_i4_3_lut (.A(\next_pc_for_core[6] ), .B(return_addr[6]), 
         .C(debug_ret), .Z(n36[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i4_3_lut.init = 16'hcaca;
    PFUMX mux_1956_i4 (.BLUT(n3163[3]), .ALUT(n3196[3]), .C0(n4073), .Z(n3314[3]));
    LUT4 mux_345_i5_3_lut (.A(\next_pc_for_core[7] ), .B(return_addr[7]), 
         .C(debug_ret), .Z(n36[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i5_3_lut.init = 16'hcaca;
    LUT4 n26926_bdd_3_lut_3_lut_4_lut (.A(n27376), .B(counter_hi[2]), .C(n26926), 
         .D(\imm[1] ), .Z(n26927)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam n26926_bdd_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_345_i6_3_lut (.A(\next_pc_for_core[8] ), .B(return_addr[8]), 
         .C(debug_ret), .Z(n36[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i6_3_lut.init = 16'hcaca;
    LUT4 mux_345_i7_3_lut (.A(\next_pc_for_core[9] ), .B(return_addr[9]), 
         .C(debug_ret), .Z(n36[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i7_3_lut.init = 16'hcaca;
    LUT4 mux_345_i8_3_lut (.A(\next_pc_for_core[10] ), .B(return_addr[10]), 
         .C(debug_ret), .Z(n36[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_353 (.A(\imm[1] ), .B(n27329), .C(\imm[2] ), .D(imm[0]), 
         .Z(n8900)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_adj_353.init = 16'h0110;
    LUT4 next_pc_for_core_23__I_0_i157_3_lut (.A(\next_pc_for_core[8] ), .B(\next_pc_for_core[12] ), 
         .C(counter_hi[2]), .Z(n157_adj_2644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i157_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_354 (.A(clk_c_enable_34), .B(rst_reg_n), 
         .C(n16_adj_2645), .D(n27179), .Z(n4073)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i1_2_lut_3_lut_4_lut_adj_354.init = 16'h0080;
    PFUMX mux_1956_i2 (.BLUT(n3163[1]), .ALUT(n3196[1]), .C0(n4073), .Z(n3314[1]));
    LUT4 mux_345_i9_3_lut (.A(\next_pc_for_core[11] ), .B(return_addr[11]), 
         .C(debug_ret), .Z(n36[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i9_3_lut.init = 16'hcaca;
    LUT4 mux_345_i10_3_lut (.A(\next_pc_for_core[12] ), .B(return_addr[12]), 
         .C(debug_ret), .Z(n36[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i10_3_lut.init = 16'hcaca;
    LUT4 cy_I_0_3_lut_rep_627_3_lut_4_lut (.A(n27376), .B(counter_hi[2]), 
         .C(cy_adj_2646), .D(n27267), .Z(n27252)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam cy_I_0_3_lut_rep_627_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_345_i11_3_lut (.A(\next_pc_for_core[13] ), .B(return_addr[13]), 
         .C(debug_ret), .Z(n36[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i11_3_lut.init = 16'hcaca;
    LUT4 mux_345_i12_3_lut (.A(\next_pc_for_core[14] ), .B(return_addr[14]), 
         .C(debug_ret), .Z(n36[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i12_3_lut.init = 16'hcaca;
    PFUMX mux_1947_i9 (.BLUT(n22637), .ALUT(n22721), .C0(n4071), .Z(n3273[8]));
    LUT4 i1_3_lut_4_lut_4_lut (.A(interrupt_core), .B(n27343), .C(n27305), 
         .D(n27332), .Z(n611[1])) /* synthesis lut_function=(A (B)+!A !((D)+!C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h88d8;
    LUT4 i16_4_lut (.A(n23412), .B(clk_c_enable_34), .C(rst_reg_n), .D(n27088), 
         .Z(clk_c_enable_227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i16_4_lut.init = 16'hcfca;
    LUT4 mux_345_i13_3_lut (.A(\next_pc_for_core[15] ), .B(return_addr[15]), 
         .C(debug_ret), .Z(n36[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i13_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_355 (.A(n4079), .B(n23856), .C(n27109), .D(n27106), 
         .Z(n23412)) /* synthesis lut_function=(A+!((C+!(D))+!B)) */ ;
    defparam i1_4_lut_adj_355.init = 16'haeaa;
    LUT4 mux_345_i14_3_lut (.A(\next_pc_for_core[16] ), .B(return_addr[16]), 
         .C(debug_ret), .Z(n36[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i14_3_lut.init = 16'hcaca;
    LUT4 mux_345_i15_3_lut (.A(\next_pc_for_core[17] ), .B(return_addr[17]), 
         .C(debug_ret), .Z(n36[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i15_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_356 (.A(n27112), .B(n35), .C(n23868), .D(n26), 
         .Z(n23856)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_356.init = 16'h5040;
    PFUMX mux_1947_i7 (.BLUT(n3087[6]), .ALUT(n22733), .C0(n4071), .Z(n3273[6]));
    LUT4 mux_345_i16_3_lut (.A(\next_pc_for_core[18] ), .B(return_addr[18]), 
         .C(debug_ret), .Z(n36[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i16_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_357 (.A(n27211), .B(n26869), .C(n28), .Z(n26)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_adj_357.init = 16'hecec;
    LUT4 i1_4_lut_adj_358 (.A(n824), .B(n27111), .C(is_load), .D(mem_op[1]), 
         .Z(n22866)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_4_lut_adj_358.init = 16'hffef;
    PFUMX mux_1947_i4 (.BLUT(n3087[3]), .ALUT(n22559), .C0(n4071), .Z(n3273[3]));
    LUT4 mux_345_i17_3_lut (.A(\next_pc_for_core[19] ), .B(return_addr[19]), 
         .C(debug_ret), .Z(n36[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i17_3_lut.init = 16'hcaca;
    LUT4 mux_1326_i15_3_lut (.A(n5[14]), .B(n31[14]), .C(n2035), .Z(n2036[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i15_3_lut.init = 16'hcaca;
    LUT4 mux_345_i18_3_lut (.A(\next_pc_for_core[20] ), .B(return_addr[20]), 
         .C(debug_ret), .Z(n36[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i15_3_lut (.A(n33[14]), .B(n1[14]), .C(n2055), .Z(n2056[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i15_3_lut.init = 16'hcaca;
    LUT4 mux_345_i19_3_lut (.A(\next_pc_for_core[21] ), .B(return_addr[21]), 
         .C(debug_ret), .Z(n36[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i19_3_lut.init = 16'hcaca;
    LUT4 mux_345_i20_3_lut (.A(\next_pc_for_core[22] ), .B(return_addr[22]), 
         .C(debug_ret), .Z(n36[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i20_3_lut.init = 16'hcaca;
    LUT4 mux_1336_i2_rep_138_3_lut (.A(n2036[1]), .B(n2056[1]), .C(n27260), 
         .Z(n25707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i2_rep_138_3_lut.init = 16'hcaca;
    PFUMX mux_1947_i2 (.BLUT(n3087[1]), .ALUT(n3126[1]), .C0(n4071), .Z(n3273[1]));
    LUT4 i2_4_lut (.A(n27179), .B(clk_c_enable_282), .C(n27185), .D(n27184), 
         .Z(n4079)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'hc888;
    LUT4 i22303_3_lut_4_lut (.A(n27200), .B(n27199), .C(n27201), .D(n7), 
         .Z(n24583)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22303_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_345_i21_3_lut (.A(\next_pc_for_core[23] ), .B(return_addr[23]), 
         .C(debug_ret), .Z(n36[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i21_3_lut.init = 16'hcaca;
    LUT4 mux_1326_i16_3_lut (.A(n5[15]), .B(n31[15]), .C(n2035), .Z(n2036[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i16_3_lut.init = 16'hcaca;
    LUT4 n3193_bdd_4_lut (.A(n27084), .B(n4071), .C(n22551), .D(n27197), 
         .Z(n26117)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (C))) */ ;
    defparam n3193_bdd_4_lut.init = 16'he2c0;
    LUT4 mux_1330_i16_3_lut (.A(n33[15]), .B(n1[15]), .C(n2055), .Z(n2056[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1326_i14_3_lut (.A(n5[13]), .B(n31[13]), .C(n2035), .Z(n2036[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i14_3_lut (.A(n33[13]), .B(n1[13]), .C(n2055), .Z(n2056[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1956_i13_3_lut_3_lut_4_lut (.A(n26), .B(n27092), .C(n4625[11]), 
         .D(n3273[10]), .Z(n3314[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1956_i13_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 i38_3_lut (.A(n28564), .B(n27209), .C(n24_adj_2656), .Z(n22_adj_2640)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;
    defparam i38_3_lut.init = 16'h9898;
    LUT4 mux_1096_i2_4_lut (.A(n27199), .B(rs2[1]), .C(n27109), .D(n27372), 
         .Z(n1794[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1096_i2_4_lut.init = 16'h3aca;
    LUT4 i1_3_lut_adj_359 (.A(additional_mem_ops[1]), .B(additional_mem_ops[0]), 
         .C(additional_mem_ops[2]), .Z(any_additional_mem_ops)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(137[35:63])
    defparam i1_3_lut_adj_359.init = 16'hfefe;
    LUT4 mux_1096_i3_4_lut (.A(n27200), .B(rs2[2]), .C(n27109), .D(n27304), 
         .Z(n1794[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1096_i3_4_lut.init = 16'h3aca;
    LUT4 mux_1096_i4_4_lut (.A(n27198), .B(rs2[3]), .C(n27109), .D(n5839), 
         .Z(n1794[3])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1096_i4_4_lut.init = 16'h3aca;
    LUT4 i5499_4_lut (.A(n24642), .B(instr[26]), .C(n4075), .D(n27131), 
         .Z(n3232[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i5499_4_lut.init = 16'hca0a;
    LUT4 debug_instr_valid_N_433_I_0_4_lut (.A(debug_instr_valid), .B(is_store), 
         .C(no_write_in_progress), .D(is_load), .Z(stall_core)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(148[23:87])
    defparam debug_instr_valid_N_433_I_0_4_lut.init = 16'h5f5d;
    PFUMX mux_1960_i4 (.BLUT(n24632), .ALUT(n3232[3]), .C0(n24998), .Z(n3350[3]));
    LUT4 mux_1336_i2_rep_139_3_lut (.A(n2036[1]), .B(n2056[1]), .C(n27260), 
         .Z(n25708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i2_rep_139_3_lut.init = 16'hcaca;
    FD1P3AX rs2_i0_i1 (.D(n1815[1]), .SP(clk_c_enable_372), .CK(clk_c), 
            .Q(rs2[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i1.GSR = "DISABLED";
    FD1P3AX rs2_i0_i2 (.D(n1815[2]), .SP(clk_c_enable_372), .CK(clk_c), 
            .Q(rs2[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i2.GSR = "DISABLED";
    FD1P3AX rs2_i0_i3 (.D(n1815[3]), .SP(clk_c_enable_372), .CK(clk_c), 
            .Q(rs2[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i3.GSR = "DISABLED";
    PFUMX mux_1960_i3 (.BLUT(n24634), .ALUT(n3232[2]), .C0(n24998), .Z(n3350[2]));
    FD1P3IX pc_offset__i22 (.D(pc_23__N_911[19]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[22] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i22.GSR = "DISABLED";
    FD1P3IX pc_offset__i21 (.D(pc_23__N_911[18]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[21] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i21.GSR = "DISABLED";
    FD1P3IX pc_offset__i20 (.D(pc_23__N_911[17]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[20] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i20.GSR = "DISABLED";
    FD1P3IX pc_offset__i19 (.D(pc_23__N_911[16]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[19] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i19.GSR = "DISABLED";
    FD1P3IX pc_offset__i18 (.D(pc_23__N_911[15]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[18] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i18.GSR = "DISABLED";
    FD1P3IX pc_offset__i17 (.D(pc_23__N_911[14]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[17] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i17.GSR = "DISABLED";
    FD1P3IX pc_offset__i16 (.D(pc_23__N_911[13]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[16] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i16.GSR = "DISABLED";
    FD1P3IX pc_offset__i15 (.D(pc_23__N_911[12]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[15] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i15.GSR = "DISABLED";
    FD1P3IX pc_offset__i14 (.D(pc_23__N_911[11]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[14] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i14.GSR = "DISABLED";
    FD1P3IX pc_offset__i13 (.D(pc_23__N_911[10]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[13] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i13.GSR = "DISABLED";
    FD1P3IX pc_offset__i12 (.D(pc_23__N_911[9]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[12] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i12.GSR = "DISABLED";
    FD1P3IX pc_offset__i11 (.D(pc_23__N_911[8]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[11] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i11.GSR = "DISABLED";
    FD1P3IX pc_offset__i10 (.D(pc_23__N_911[7]), .SP(clk_c_enable_423), 
            .CD(n27326), .CK(clk_c), .Q(\pc[10] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i10.GSR = "DISABLED";
    FD1P3IX pc_offset__i9 (.D(pc_23__N_911[6]), .SP(clk_c_enable_423), .CD(n27326), 
            .CK(clk_c), .Q(\pc[9] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i9.GSR = "DISABLED";
    FD1P3IX pc_offset__i8 (.D(pc_23__N_911[5]), .SP(clk_c_enable_423), .CD(n27326), 
            .CK(clk_c), .Q(\pc[8] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i8.GSR = "DISABLED";
    FD1P3IX pc_offset__i7 (.D(pc_23__N_911[4]), .SP(clk_c_enable_423), .CD(n27326), 
            .CK(clk_c), .Q(\pc[7] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i7.GSR = "DISABLED";
    FD1P3IX pc_offset__i6 (.D(pc_23__N_911[3]), .SP(clk_c_enable_423), .CD(n27326), 
            .CK(clk_c), .Q(\pc[6] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i6.GSR = "DISABLED";
    FD1P3IX pc_offset__i5 (.D(pc_23__N_911[2]), .SP(clk_c_enable_423), .CD(n27326), 
            .CK(clk_c), .Q(\pc[5] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i5.GSR = "DISABLED";
    FD1P3IX pc_offset__i4 (.D(pc_23__N_911[1]), .SP(clk_c_enable_423), .CD(n27326), 
            .CK(clk_c), .Q(\pc[4] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i4.GSR = "DISABLED";
    FD1P3IX pc_offset__i3 (.D(pc_23__N_911[0]), .SP(clk_c_enable_423), .CD(n27326), 
            .CK(clk_c), .Q(\pc[3] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i3.GSR = "DISABLED";
    PFUMX mux_1975_i19 (.BLUT(n3163[29]), .ALUT(n3314[19]), .C0(n25083), 
          .Z(n3397[17]));
    FD1P3IX pc_offset__i2 (.D(pc_2__N_932[1]), .SP(clk_c_enable_423), .CD(n27326), 
            .CK(clk_c), .Q(\pc[2] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i2.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_360 (.A(rd[3]), .B(n27113), .C(any_additional_mem_ops), 
         .D(n5868), .Z(n22887)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(149[27:88])
    defparam i1_4_lut_adj_360.init = 16'h4080;
    LUT4 mux_1956_i17_3_lut_3_lut_4_lut (.A(n26), .B(n27092), .C(n4625[15]), 
         .D(n3273[10]), .Z(n3314[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1956_i17_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1956_i14_3_lut_3_lut_4_lut (.A(n26), .B(n27092), .C(n4625[12]), 
         .D(n3273[10]), .Z(n3314[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1956_i14_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_361 (.A(rd[2]), .B(n27113), .C(any_additional_mem_ops), 
         .D(n27371), .Z(n22888)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(149[27:88])
    defparam i1_4_lut_adj_361.init = 16'h4080;
    LUT4 mux_1077_i8_3_lut (.A(n1[7]), .B(n5[7]), .C(n2055), .Z(n1735[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i8_3_lut.init = 16'hcaca;
    LUT4 is_lui_I_0_473_2_lut_rep_694 (.A(is_lui), .B(debug_instr_valid), 
         .Z(n27319)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam is_lui_I_0_473_2_lut_rep_694.init = 16'h8888;
    LUT4 i1_4_lut_adj_362 (.A(any_additional_mem_ops), .B(n27113), .C(rd[1]), 
         .D(rd[0]), .Z(n22889)) /* synthesis lut_function=(!(((C (D)+!C !(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(149[27:88])
    defparam i1_4_lut_adj_362.init = 16'h0880;
    LUT4 i1_2_lut (.A(n27112), .B(n8274), .Z(n23682)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    L6MUX21 mux_1576_i4 (.D0(n2368[3]), .D1(n2376[3]), .SD(n2704), .Z(n2386[3]));
    LUT4 mux_1073_i8_rep_95_3_lut (.A(n31[7]), .B(n33[7]), .C(n2035), 
         .Z(n24638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i8_rep_95_3_lut.init = 16'hcaca;
    L6MUX21 mux_1576_i3 (.D0(n2368[2]), .D1(n2376[2]), .SD(n2704), .Z(n2386[2]));
    LUT4 i22726_3_lut_4_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(n25066), 
         .D(n27349), .Z(n25069)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i22726_3_lut_4_lut_4_lut.init = 16'h4000;
    L6MUX21 mux_1576_i2 (.D0(n2368[1]), .D1(n2376[1]), .SD(n2704), .Z(n2386[1]));
    LUT4 mux_91_i1_3_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(debug_rd_3__N_405[28]), 
         .D(n157_adj_2644), .Z(n234[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam mux_91_i1_3_lut_4_lut.init = 16'hf780;
    L6MUX21 mux_1393_i2 (.D0(n2152[1]), .D1(n2161[1]), .SD(n2330), .Z(n2175[1]));
    L6MUX21 mux_1576_i1 (.D0(n2368[0]), .D1(n2376[0]), .SD(n2704), .Z(n2386[0]));
    LUT4 mux_1956_i15_3_lut_3_lut_4_lut (.A(n26), .B(n27092), .C(n4625[13]), 
         .D(n3273[10]), .Z(n3314[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1956_i15_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1956_i12_3_lut_3_lut_4_lut (.A(n26), .B(n27092), .C(n3163[11]), 
         .D(n3273[10]), .Z(n3314[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1956_i12_3_lut_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_1393_i1 (.BLUT(n2152[0]), .ALUT(n2161[0]), .C0(n2330), .Z(n2175[0]));
    LUT4 i1_2_lut_rep_696 (.A(debug_instr_valid), .B(no_write_in_progress), 
         .Z(n27321)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_2_lut_rep_696.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_363 (.A(debug_instr_valid), .B(no_write_in_progress), 
         .C(load_done), .D(is_load), .Z(instr_complete_N_1651)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_3_lut_4_lut_adj_363.init = 16'h8000;
    LUT4 i23384_3_lut (.A(n3232[12]), .B(n4703[12]), .C(n4075), .Z(n3350[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23384_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_364 (.A(n27170), .B(n7), .C(n27199), .D(n27209), 
         .Z(n22100)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_364.init = 16'h0100;
    LUT4 i23382_3_lut (.A(n3232[13]), .B(n4703[13]), .C(n4075), .Z(n3350[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23382_3_lut.init = 16'hcaca;
    LUT4 i23380_3_lut (.A(n3232[14]), .B(n4703[14]), .C(n4075), .Z(n3350[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23380_3_lut.init = 16'hcaca;
    LUT4 i23378_3_lut (.A(n3232[15]), .B(n4703[15]), .C(n4075), .Z(n3350[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23378_3_lut.init = 16'hcaca;
    LUT4 i30_3_lut_4_lut_3_lut (.A(n28564), .B(n27212), .C(n27209), .Z(n13)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam i30_3_lut_4_lut_3_lut.init = 16'h1818;
    LUT4 mux_1956_i11_3_lut_3_lut_4_lut (.A(n26), .B(n27092), .C(n3163[10]), 
         .D(n3273[10]), .Z(n3314[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1956_i11_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_365 (.A(clk_c_enable_34), .B(n28575), 
         .C(n19), .D(n27179), .Z(n4065)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i1_2_lut_3_lut_4_lut_adj_365.init = 16'h0080;
    LUT4 mux_1956_i16_3_lut_3_lut_4_lut (.A(n26), .B(n27092), .C(n4625[14]), 
         .D(n3273[10]), .Z(n3314[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1956_i16_3_lut_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_1960_i17 (.BLUT(n3232[16]), .ALUT(n4703[16]), .C0(n4075), 
          .Z(n3350[16]));
    LUT4 i1_2_lut_rep_463_3_lut_4_lut (.A(clk_c_enable_34), .B(rst_reg_n), 
         .C(n22_adj_2640), .D(n27179), .Z(n27088)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i1_2_lut_rep_463_3_lut_4_lut.init = 16'h0080;
    LUT4 mux_1984_i30_3_lut_4_lut (.A(n4079), .B(n4075), .C(n3350[24]), 
         .D(n4703[29]), .Z(n3438[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1984_i30_3_lut_4_lut.init = 16'hf870;
    LUT4 i22_4_lut_4_lut (.A(n27212), .B(n28564), .C(n22100), .D(n27178), 
         .Z(n8_adj_2657)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam i22_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i12351_2_lut_3_lut (.A(n28564), .B(n27209), .C(n15_adj_2658), 
         .Z(mem_op_de[0])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    defparam i12351_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i2_2_lut_3_lut (.A(n28564), .B(n27209), .C(n27211), .Z(n17)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    defparam i2_2_lut_3_lut.init = 16'h4040;
    LUT4 mux_1984_i29_3_lut_4_lut (.A(n4079), .B(n4075), .C(n3350[24]), 
         .D(n4703[28]), .Z(n3438[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1984_i29_3_lut_4_lut.init = 16'hf870;
    PFUMX mux_1960_i5 (.BLUT(n3232[4]), .ALUT(n4703[4]), .C0(n4075), .Z(n3350[4]));
    LUT4 mux_1336_i15_3_lut_rep_759 (.A(n2036[14]), .B(n2056[14]), .C(n27260), 
         .Z(n28563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i15_3_lut_rep_759.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_366 (.A(clk_c_enable_34), .B(n28575), 
         .C(n26_adj_2659), .D(n27179), .Z(n4063)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i1_2_lut_3_lut_4_lut_adj_366.init = 16'h0080;
    LUT4 i22414_3_lut (.A(\mem_data_from_read[19] ), .B(\mem_data_from_read[23] ), 
         .C(counter_hi[2]), .Z(n24757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22414_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_367 (.A(n27191), .B(n22534), .C(n24525), .D(n27211), 
         .Z(n22674)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_367.init = 16'h0004;
    LUT4 mux_1383_i4_4_lut (.A(n4625[8]), .B(instr[18]), .C(n2328), .D(n27179), 
         .Z(n2161[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam mux_1383_i4_4_lut.init = 16'hca0a;
    LUT4 i1_3_lut_4_lut_3_lut (.A(n28564), .B(n27209), .C(n27212), .Z(n20)) /* synthesis lut_function=(A (B+(C))+!A !(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    defparam i1_3_lut_4_lut_3_lut.init = 16'hb9b9;
    LUT4 i1_4_lut_adj_368 (.A(was_early_branch), .B(n8486), .C(n16_adj_2660), 
         .D(n27179), .Z(n8274)) /* synthesis lut_function=(A+(B (C (D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[82:120])
    defparam i1_4_lut_adj_368.init = 16'hfaba;
    LUT4 i2_2_lut_3_lut_adj_369 (.A(n28564), .B(n27209), .C(n27212), .Z(n11)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    defparam i2_2_lut_3_lut_adj_369.init = 16'h4040;
    LUT4 i2_2_lut_3_lut_4_lut (.A(clk_c_enable_34), .B(n28575), .C(n22), 
         .D(n27179), .Z(n2326)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i4694_4_lut_4_lut (.A(clk_c_enable_34), .B(n27157), .C(additional_mem_ops[0]), 
         .D(n27201), .Z(additional_mem_ops_de[0])) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i4694_4_lut_4_lut.init = 16'hd850;
    PFUMX mux_1378_i2 (.BLUT(n2120[1]), .ALUT(n2128[1]), .C0(n2326), .Z(n2152[1]));
    LUT4 i1_2_lut_rep_702 (.A(\instr_addr_23__N_318[0] ), .B(instr_addr_23__N_318[1]), 
         .Z(n27327)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_rep_702.init = 16'hbbbb;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\instr_addr_23__N_318[0] ), .B(instr_addr_23__N_318[1]), 
         .C(n28575), .Z(n23564)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_2_lut_3_lut.init = 16'hbfbf;
    PFUMX mux_1393_i4 (.BLUT(n22784), .ALUT(n2161[3]), .C0(n2330), .Z(n2175[3]));
    LUT4 i5394_4_lut_4_lut (.A(clk_c_enable_34), .B(n27157), .C(additional_mem_ops[1]), 
         .D(n27199), .Z(additional_mem_ops_de[1])) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i5394_4_lut_4_lut.init = 16'hd850;
    LUT4 mux_1984_i25_3_lut_4_lut (.A(n4079), .B(n4075), .C(n3350[24]), 
         .D(n4703[24]), .Z(n3438[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1984_i25_3_lut_4_lut.init = 16'hf870;
    LUT4 i23576_2_lut_rep_527_3_lut (.A(n28564), .B(n28563), .C(n27212), 
         .Z(n27152)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i23576_2_lut_rep_527_3_lut.init = 16'h1010;
    PFUMX mux_1566_i4 (.BLUT(n22674), .ALUT(n2342[3]), .C0(n2700), .Z(n2368[3]));
    LUT4 mux_1938_i5_3_lut (.A(n27203), .B(instr[24]), .C(n27099), .Z(n3232[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1938_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1083_i5_rep_81_3_lut (.A(n1735[4]), .B(n27206), .C(n4057), 
         .Z(n24624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i5_rep_81_3_lut.init = 16'hcaca;
    PFUMX mux_1566_i3 (.BLUT(n22671), .ALUT(n2342[2]), .C0(n2700), .Z(n2368[2]));
    LUT4 i12710_2_lut_3_lut_4_lut (.A(n28564), .B(n28563), .C(n27211), 
         .D(n27212), .Z(n30)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i12710_2_lut_3_lut_4_lut.init = 16'h1000;
    PFUMX mux_1566_i2 (.BLUT(n22667), .ALUT(n2342[1]), .C0(n2700), .Z(n2368[1]));
    LUT4 i49_3_lut_3_lut (.A(n28564), .B(n28563), .C(n27209), .Z(n28)) /* synthesis lut_function=(!(A (C)+!A (B+!(C)))) */ ;
    defparam i49_3_lut_3_lut.init = 16'h1a1a;
    LUT4 i23386_3_lut (.A(n24624), .B(n3232[11]), .C(n25004), .Z(n3350[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23386_3_lut.init = 16'hcaca;
    PFUMX mux_1933_i8 (.BLUT(n4625[6]), .ALUT(n2874[7]), .C0(n4065), .Z(n3163[7]));
    LUT4 i20060_2_lut_rep_705 (.A(\imm[7] ), .B(\imm[11] ), .Z(n27330)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20060_2_lut_rep_705.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_370 (.A(\imm[7] ), .B(\imm[11] ), .C(n8900), 
         .D(n22088), .Z(n5160)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_370.init = 16'h1000;
    LUT4 i12704_2_lut_3_lut_4_lut (.A(n28564), .B(n28563), .C(n27207), 
         .D(n27190), .Z(n30_adj_2661)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i12704_2_lut_3_lut_4_lut.init = 16'h1000;
    PFUMX mux_1566_i1 (.BLUT(n22663), .ALUT(n2342[0]), .C0(n2700), .Z(n2368[0]));
    LUT4 i12708_2_lut_3_lut_4_lut (.A(n28564), .B(n28563), .C(n27202), 
         .D(n27190), .Z(n30_adj_2662)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i12708_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i22402_3_lut (.A(\mem_data_from_read[16] ), .B(\mem_data_from_read[20] ), 
         .C(counter_hi[2]), .Z(n24745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22402_3_lut.init = 16'hcaca;
    LUT4 i22408_3_lut (.A(\mem_data_from_read[18] ), .B(\mem_data_from_read[22] ), 
         .C(counter_hi[2]), .Z(n24751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22408_3_lut.init = 16'hcaca;
    LUT4 mux_1083_i7_rep_91_3_lut_3_lut (.A(n27099), .B(n27207), .C(n1735[6]), 
         .Z(n24634)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1083_i7_rep_91_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_1383_i1_4_lut (.A(n2133[0]), .B(n27212), .C(n2328), .D(n27179), 
         .Z(n2161[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam mux_1383_i1_4_lut.init = 16'hca0a;
    LUT4 mux_1956_i1_4_lut (.A(n23594), .B(n8274), .C(n4073), .D(n23726), 
         .Z(n24601)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1956_i1_4_lut.init = 16'h3a0a;
    LUT4 mux_1083_i8_rep_89_3_lut_3_lut (.A(n27099), .B(n27204), .C(n1735[7]), 
         .Z(n24632)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1083_i8_rep_89_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_1984_i26_3_lut_4_lut (.A(n4079), .B(n4075), .C(n3350[24]), 
         .D(n4703[25]), .Z(n3438[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1984_i26_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_1938_i17_3_lut_4_lut (.A(n27101), .B(n27127), .C(n4745[9]), 
         .D(n24664), .Z(n3232[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1938_i17_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_4_lut_adj_371 (.A(n824), .B(n27111), .C(address_ready), .D(is_load), 
         .Z(clk_c_enable_280)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_371.init = 16'hfeff;
    LUT4 i1_4_lut_adj_372 (.A(n824), .B(n27111), .C(is_load), .D(mem_op[0]), 
         .Z(n22867)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_4_lut_adj_372.init = 16'hffef;
    PFUMX mux_1933_i5 (.BLUT(n4625[3]), .ALUT(n2874[4]), .C0(n4065), .Z(n3163[4]));
    L6MUX21 i23765 (.D0(n26118), .D1(n3350[2]), .SD(n4079), .Z(n26119));
    LUT4 i1_2_lut_rep_708 (.A(\instr_addr_23__N_318[0] ), .B(instr_addr_23__N_318[1]), 
         .Z(n27333)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_rep_708.init = 16'hdddd;
    LUT4 i1_2_lut_2_lut_3_lut_adj_373 (.A(\instr_addr_23__N_318[0] ), .B(instr_addr_23__N_318[1]), 
         .C(n28575), .Z(n23572)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i1_2_lut_2_lut_3_lut_adj_373.init = 16'hdfdf;
    LUT4 i1_2_lut_rep_709 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .Z(n27334)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_709.init = 16'heeee;
    LUT4 i1_2_lut_2_lut_3_lut_adj_374 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .C(n28575), .Z(n23580)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_2_lut_3_lut_adj_374.init = 16'hefef;
    LUT4 i12317_3_lut (.A(n27206), .B(n2326), .C(n2322), .Z(n2152[0])) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam i12317_3_lut.init = 16'hc8c8;
    LUT4 mux_40_i4_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[31]), 
         .D(data_rs2[3]), .Z(n92[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_40_i3_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[30]), 
         .D(data_rs2[2]), .Z(n92[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i3_3_lut_4_lut.init = 16'hf780;
    PFUMX i23763 (.BLUT(n26117), .ALUT(n26116), .C0(n27086), .Z(n26118));
    LUT4 mux_40_i2_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[29]), 
         .D(data_rs2[1]), .Z(n92[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_40_i1_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[28]), 
         .D(data_rs2[0]), .Z(n92[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i23607_2_lut_rep_712 (.A(counter_hi[3]), .B(n28571), .Z(clk_c_enable_424)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i23607_2_lut_rep_712.init = 16'h7777;
    LUT4 i12883_2_lut_rep_670_3_lut (.A(n28573), .B(n28571), .C(counter_hi[2]), 
         .Z(clk_c_enable_276)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i12883_2_lut_rep_670_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_638_3_lut_4_lut (.A(n28573), .B(n28571), .C(any_additional_mem_ops), 
         .D(counter_hi[2]), .Z(n27263)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_638_3_lut_4_lut.init = 16'h0800;
    LUT4 i12232_2_lut_rep_485_3_lut_4_lut (.A(n28573), .B(n28571), .C(instr_complete_N_1647), 
         .D(counter_hi[2]), .Z(n27110)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12232_2_lut_rep_485_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_375 (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(mcause[5]), .D(counter_hi[2]), .Z(n24216)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_375.init = 16'h8000;
    LUT4 i20179_rep_133_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n22499), .D(counter_hi[2]), .Z(n25702)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20179_rep_133_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i20179_rep_134_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n22499), .D(counter_hi[2]), .Z(n25703)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20179_rep_134_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i20179_rep_135_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n22499), .D(counter_hi[2]), .Z(n25704)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20179_rep_135_2_lut_3_lut_4_lut.init = 16'h8000;
    PFUMX mux_1383_i2 (.BLUT(n9124), .ALUT(n2138[1]), .C0(n2328), .Z(n2161[1]));
    LUT4 i20179_rep_136_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n22499), .D(counter_hi[2]), .Z(n25705)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20179_rep_136_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23584_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), .C(rst_reg_n), 
         .Z(n9675)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam i23584_2_lut_3_lut.init = 16'h0707;
    LUT4 i12894_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n27300), .D(counter_hi[2]), .Z(clk_c_enable_20)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12894_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i20179_rep_489_3_lut_4_lut (.A(n28573), .B(n28571), .C(n22499), 
         .D(counter_hi[2]), .Z(n27114)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20179_rep_489_3_lut_4_lut.init = 16'h8000;
    LUT4 i20179_rep_137_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n22499), .D(counter_hi[2]), .Z(n25706)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20179_rep_137_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_376 (.A(n28573), .B(n28571), .C(\imm[6] ), 
         .Z(n22121)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_376.init = 16'h7070;
    PFUMX mux_1109_i4 (.BLUT(n1804[3]), .ALUT(n1794[3]), .C0(n2031), .Z(n1815[3]));
    PFUMX mux_1109_i3 (.BLUT(n1804[2]), .ALUT(n1794[2]), .C0(n2031), .Z(n1815[2]));
    LUT4 i3916_2_lut (.A(\instr_addr_23__N_318[0] ), .B(\pc[1] ), .Z(n2)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i3916_2_lut.init = 16'hbbbb;
    LUT4 mux_1960_i27_3_lut_4_lut (.A(n4079), .B(n4075), .C(n3350[24]), 
         .D(n24642), .Z(n3350[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1960_i27_3_lut_4_lut.init = 16'hf870;
    LUT4 i12261_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), .C(mepc[0]), 
         .Z(csr_read_3__N_1451[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12261_2_lut_3_lut.init = 16'h7070;
    PFUMX mux_1109_i2 (.BLUT(n1804[1]), .ALUT(n1794[1]), .C0(n2031), .Z(n1815[1]));
    LUT4 i1_3_lut_adj_377 (.A(next_pc_offset[3]), .B(n4), .C(\instr_write_offset[3] ), 
         .Z(n23087)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i1_3_lut_adj_377.init = 16'h9696;
    PFUMX mux_1570_i2 (.BLUT(n2347[1]), .ALUT(n22889), .C0(n2702), .Z(n2376[1]));
    LUT4 i1_rep_44_4_lut (.A(is_ret_de), .B(n27108), .C(n8), .D(n22369), 
         .Z(n22592)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[18] 227[12])
    defparam i1_rep_44_4_lut.init = 16'h0800;
    LUT4 i23719_3_lut_4_lut (.A(n27131), .B(n27260), .C(n4075), .D(n4079), 
         .Z(n24900)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23719_3_lut_4_lut.init = 16'h1fff;
    PFUMX mux_1570_i3 (.BLUT(n2347[2]), .ALUT(n22888), .C0(n2702), .Z(n2376[2]));
    LUT4 i1_4_lut_adj_378 (.A(n27108), .B(n8), .C(n27114), .D(n23238), 
         .Z(debug_early_branch)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_378.init = 16'h0200;
    LUT4 i1_2_lut_adj_379 (.A(is_jal_de), .B(n28575), .Z(n23238)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_379.init = 16'h8888;
    LUT4 i1_4_lut_adj_380 (.A(n23292), .B(n27109), .C(n8274), .D(instr_complete_N_1647), 
         .Z(n8)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_380.init = 16'hfefc;
    LUT4 mux_1326_i10_3_lut (.A(n5[9]), .B(n31[9]), .C(n2035), .Z(n2036[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i10_3_lut (.A(n33[9]), .B(n1[9]), .C(n2055), .Z(n2056[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1326_i8_3_lut (.A(n5[7]), .B(n31[7]), .C(n2035), .Z(n2036[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i8_3_lut.init = 16'hcaca;
    PFUMX mux_1570_i4 (.BLUT(n2347[3]), .ALUT(n22887), .C0(n2702), .Z(n2376[3]));
    LUT4 mux_1330_i8_3_lut (.A(n33[7]), .B(n1[7]), .C(n2055), .Z(n2056[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1326_i13_3_lut (.A(n5[12]), .B(n31[12]), .C(n2035), .Z(n2036[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i13_3_lut (.A(n33[12]), .B(n1[12]), .C(n2055), .Z(n2056[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1938_i3_4_lut (.A(n24637), .B(n27207), .C(n4075), .D(n27131), 
         .Z(n3232[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1938_i3_4_lut.init = 16'hca0a;
    LUT4 mux_1326_i11_3_lut (.A(n5[10]), .B(n31[10]), .C(n2035), .Z(n2036[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i11_3_lut (.A(n33[10]), .B(n1[10]), .C(n2055), .Z(n2056[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i11_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_716 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .Z(n27341)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_716.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_381 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .C(n28575), .Z(n23558)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_381.init = 16'h8080;
    LUT4 i22311_3_lut_rep_717 (.A(counter_hi[2]), .B(n28573), .C(n28571), 
         .Z(n27342)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i22311_3_lut_rep_717.init = 16'h8080;
    LUT4 i23441_2_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), .C(counter_hi[4]), 
         .D(rst_reg_n), .Z(clk_c_enable_100)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;
    defparam i23441_2_lut_4_lut.init = 16'h80ff;
    PFUMX mux_1960_i1 (.BLUT(n22909), .ALUT(n4703[0]), .C0(n4075), .Z(n3350[0]));
    PFUMX mux_1109_i1 (.BLUT(n1804[0]), .ALUT(n1794[0]), .C0(n2031), .Z(n1815[0]));
    PFUMX mux_1570_i1 (.BLUT(n2347[0]), .ALUT(n2352[0]), .C0(n2702), .Z(n2376[0]));
    LUT4 mux_1326_i12_3_lut (.A(n5[11]), .B(n31[11]), .C(n2035), .Z(n2036[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i12_3_lut (.A(n33[11]), .B(n1[11]), .C(n2055), .Z(n2056[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i12_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_531_3_lut_4_lut (.A(n27211), .B(n27212), .C(n28563), 
         .D(n28564), .Z(n27156)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i2_2_lut_rep_531_3_lut_4_lut.init = 16'h0002;
    LUT4 mux_1938_i4_4_lut (.A(n24638), .B(n27204), .C(n4075), .D(n27131), 
         .Z(n3232[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1938_i4_4_lut.init = 16'hca0a;
    LUT4 mux_1326_i1_3_lut (.A(n5[0]), .B(n31[0]), .C(n2035), .Z(n2036[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1326_i9_3_lut (.A(n5[8]), .B(n31[8]), .C(n2035), .Z(n2036[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i9_3_lut (.A(n33[8]), .B(n1[8]), .C(n2055), .Z(n2056[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1326_i3_3_lut (.A(n5[2]), .B(n31[2]), .C(n2035), .Z(n2036[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i3_3_lut (.A(n33[2]), .B(n1[2]), .C(n2055), .Z(n2056[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i3_3_lut.init = 16'hcaca;
    PFUMX mux_1960_i7 (.BLUT(n24640), .ALUT(n3232[6]), .C0(n24988), .Z(n3350[6]));
    LUT4 mux_1326_i5_3_lut (.A(n5[4]), .B(n31[4]), .C(n2035), .Z(n2036[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i5_3_lut (.A(n33[4]), .B(n1[4]), .C(n2055), .Z(n2056[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i5_3_lut.init = 16'hcaca;
    PFUMX mux_55_i2 (.BLUT(n7711), .ALUT(additional_mem_ops_de[1]), .C0(n24817), 
          .Z(n4116[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 mux_1326_i4_3_lut (.A(n5[3]), .B(n31[3]), .C(n2035), .Z(n2036[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i4_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_3_lut (.A(imm[0]), .B(\imm[1] ), .C(\imm[6] ), .Z(n24160)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_3_lut.init = 16'h4141;
    LUT4 mux_3182_i4_4_lut_4_lut (.A(imm[0]), .B(\imm[1] ), .C(instrret_count[3]), 
         .D(cycle_count_wide[3]), .Z(n5114[3])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mux_3182_i4_4_lut_4_lut.init = 16'h7340;
    PFUMX mux_55_i1 (.BLUT(n6985), .ALUT(additional_mem_ops_de[0]), .C0(n24817), 
          .Z(n4116[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i23456_2_lut_rep_722 (.A(alu_op[1]), .B(alu_op[3]), .Z(n27347)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i23456_2_lut_rep_722.init = 16'h7777;
    LUT4 i1_3_lut_4_lut_adj_382 (.A(alu_op[1]), .B(alu_op[3]), .C(cycle[0]), 
         .D(alu_op[2]), .Z(debug_reg_wen_N_1692)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_4_lut_adj_382.init = 16'hfff7;
    LUT4 mux_1330_i4_3_lut (.A(n33[3]), .B(n1[3]), .C(n2055), .Z(n2056[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i4_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_642_4_lut_3_lut (.A(alu_op[1]), .B(alu_op[3]), .C(alu_op[2]), 
         .Z(n27267)) /* synthesis lut_function=(!(A (B (C))+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_rep_642_4_lut_3_lut.init = 16'h6e6e;
    LUT4 i12565_2_lut_rep_641_3_lut_3_lut (.A(alu_op[1]), .B(alu_op[3]), 
         .C(alu_op[2]), .Z(n27266)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i12565_2_lut_rep_641_3_lut_3_lut.init = 16'h2a2a;
    LUT4 i23722_2_lut_3_lut_4_lut (.A(alu_op[1]), .B(alu_op[3]), .C(debug_rd_3__N_413), 
         .D(alu_op[2]), .Z(n24838)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i23722_2_lut_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_645_3_lut_4_lut (.A(alu_op[1]), .B(alu_op[3]), .C(alu_op[0]), 
         .D(alu_op[2]), .Z(n27270)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_rep_645_3_lut_4_lut.init = 16'h70f0;
    LUT4 mux_1326_i6_3_lut (.A(n5[5]), .B(n31[5]), .C(n2035), .Z(n2036[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i6_3_lut (.A(n33[5]), .B(n1[5]), .C(n2055), .Z(n2056[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1326_i7_3_lut (.A(n5[6]), .B(n31[6]), .C(n2035), .Z(n2036[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1330_i7_3_lut (.A(n33[6]), .B(n1[6]), .C(n2055), .Z(n2056[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1960_i24_3_lut_4_lut (.A(n4079), .B(n4075), .C(n3350[24]), 
         .D(n24638), .Z(n3350[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1960_i24_3_lut_4_lut.init = 16'hf870;
    LUT4 i12634_1_lut_rep_649_2_lut_3_lut (.A(alu_op[1]), .B(alu_op[3]), 
         .C(alu_op[2]), .Z(n27274)) /* synthesis lut_function=(!(A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i12634_1_lut_rep_649_2_lut_3_lut.init = 16'h7f7f;
    PFUMX mux_1960_i8 (.BLUT(n3232[7]), .ALUT(n4703[7]), .C0(n4075), .Z(n3350[7]));
    LUT4 i1_3_lut_4_lut_adj_383 (.A(n27185), .B(n27128), .C(rst_reg_n), 
         .D(n27129), .Z(n23726)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_383.init = 16'h0080;
    LUT4 i1_4_lut_adj_384 (.A(n22592), .B(n27097), .C(instr_fetch_restart_N_947), 
         .D(n27227), .Z(start_instr)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(435[34:115])
    defparam i1_4_lut_adj_384.init = 16'h0010;
    LUT4 i1_rep_667_3_lut (.A(alu_op[1]), .B(alu_op[3]), .C(alu_op[2]), 
         .Z(n27292)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_rep_667_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_723 (.A(alu_op[1]), .B(alu_op[3]), .C(alu_op[2]), 
         .Z(n27348)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_rep_723.init = 16'h8080;
    PFUMX mux_1960_i6 (.BLUT(n3232[5]), .ALUT(n4703[5]), .C0(n4075), .Z(n3350[5]));
    LUT4 i1_3_lut_4_lut_adj_385 (.A(n27131), .B(n27130), .C(n23658), .D(n8274), 
         .Z(n23662)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_adj_385.init = 16'h0070;
    LUT4 i23436_4_lut (.A(n27114), .B(rst_reg_n), .C(n22592), .D(n23432), 
         .Z(clk_c_enable_175)) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;
    defparam i23436_4_lut.init = 16'h3733;
    LUT4 i12335_3_lut_rep_566 (.A(n27203), .B(n27212), .C(n28563), .Z(n27191)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i12335_3_lut_rep_566.init = 16'hc8c8;
    LUT4 i4523_2_lut_rep_556_4_lut_4_lut (.A(alu_op[1]), .B(alu_op[3]), 
         .C(alu_op[2]), .D(alu_b_in[3]), .Z(n27181)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(B (D)+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i4523_2_lut_rep_556_4_lut_4_lut.init = 16'h916e;
    LUT4 i12713_4_lut_4_lut (.A(n27211), .B(n28563), .C(n27183), .D(alu_op_3__N_1337[2]), 
         .Z(n15_adj_2663)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i12713_4_lut_4_lut.init = 16'hd0c0;
    LUT4 i1_4_lut_adj_386 (.A(n27108), .B(n8), .C(n27114), .D(n23678), 
         .Z(debug_ret)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_386.init = 16'h0200;
    LUT4 i1_3_lut_rep_499 (.A(is_timer_addr), .B(n27126), .C(data_ready_latch), 
         .Z(n27124)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(258[53:106])
    defparam i1_3_lut_rep_499.init = 16'hfbfb;
    PFUMX mux_797_i21 (.BLUT(n36[20]), .ALUT(n1222[20]), .C0(n27114), 
          .Z(pc_23__N_911[20]));
    LUT4 i23367_3_lut_4_lut_4_lut (.A(n27088), .B(n22739), .C(n4071), 
         .D(n27202), .Z(n3273[7])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i23367_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1_2_lut_adj_387 (.A(is_ret_de), .B(n28575), .Z(n23678)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_387.init = 16'h8888;
    LUT4 i1_2_lut_4_lut_adj_388 (.A(is_timer_addr), .B(n27126), .C(data_ready_latch), 
         .D(n27322), .Z(n6982)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(258[53:106])
    defparam i1_2_lut_4_lut_adj_388.init = 16'hfb00;
    LUT4 i23309_3_lut_4_lut (.A(n27201), .B(n28562), .C(n2029), .D(n23644), 
         .Z(n1804[0])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23309_3_lut_4_lut.init = 16'hefe0;
    LUT4 i23434_4_lut (.A(counter_hi[2]), .B(n27300), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(clk_c_enable_56)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam i23434_4_lut.init = 16'h0080;
    LUT4 i12164_3_lut (.A(any_additional_mem_ops), .B(rst_reg_n), .C(n27107), 
         .Z(data_continue_N_963)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i12164_3_lut.init = 16'ha8a8;
    LUT4 i53_4_lut_4_lut (.A(n27211), .B(n27209), .C(n27138), .D(n28564), 
         .Z(n32)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam i53_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i4522_2_lut_rep_562_4_lut_4_lut (.A(alu_op[1]), .B(alu_op[3]), 
         .C(alu_op[2]), .D(alu_b_in[2]), .Z(n27187)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(B (D)+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i4522_2_lut_rep_562_4_lut_4_lut.init = 16'h916e;
    LUT4 i4479_2_lut_rep_563_4_lut_4_lut (.A(alu_op[1]), .B(alu_op[3]), 
         .C(alu_op[2]), .D(alu_b_in[0]), .Z(n27188)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(B (D)+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i4479_2_lut_rep_563_4_lut_4_lut.init = 16'h916e;
    LUT4 i4521_2_lut_rep_590_4_lut_4_lut (.A(alu_op[1]), .B(alu_op[3]), 
         .C(alu_op[2]), .D(alu_b_in[1]), .Z(n27215)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(B (D)+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i4521_2_lut_rep_590_4_lut_4_lut.init = 16'h916e;
    LUT4 is_branch_I_0_475_2_lut_rep_725 (.A(is_branch), .B(debug_instr_valid), 
         .Z(n27350)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam is_branch_I_0_475_2_lut_rep_725.init = 16'h8888;
    LUT4 mux_796_i1_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[3] ), 
         .D(addr_out[3]), .Z(n1222[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i4_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[6] ), 
         .D(addr_out[6]), .Z(n1222[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2792_i2_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[2] ), .D(n27238), .Z(n4575[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_2792_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i3_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[5] ), 
         .D(addr_out[5]), .Z(n1222[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i3_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_797_i20 (.BLUT(n36[19]), .ALUT(n1222[19]), .C0(n25706), 
          .Z(pc_23__N_911[19]));
    LUT4 mux_796_i2_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[4] ), 
         .D(addr_out[4]), .Z(n1222[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1928_i2_4_lut_4_lut (.A(n27211), .B(n4063), .C(n27199), .D(n27198), 
         .Z(n3126[1])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;
    defparam mux_1928_i2_4_lut_4_lut.init = 16'h7340;
    LUT4 mux_796_i5_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[7] ), 
         .D(addr_out[7]), .Z(n1222[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i6_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[8] ), 
         .D(addr_out[8]), .Z(n1222[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 is_alu_imm_N_1367_bdd_3_lut_24161_4_lut_4_lut (.A(n27211), .B(n28563), 
         .C(n27158), .D(n27202), .Z(n26779)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;
    defparam is_alu_imm_N_1367_bdd_3_lut_24161_4_lut_4_lut.init = 16'h5d55;
    LUT4 mux_1921_i4_4_lut (.A(n27198), .B(n23516), .C(n27088), .D(n22700), 
         .Z(n3087[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1921_i4_4_lut.init = 16'hca0a;
    LUT4 mux_796_i7_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[9] ), 
         .D(addr_out[9]), .Z(n1222[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n27211), .B(n22101), .C(n28564), .D(n27209), 
         .Z(n22_adj_2664)) /* synthesis lut_function=(!(A+(B (C (D))+!B ((D)+!C)))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'h0454;
    L6MUX21 i22838 (.D0(n25179), .D1(n25180), .SD(n28571), .Z(debug_rd_3__N_405[28]));
    L6MUX21 i22845 (.D0(n25186), .D1(n25187), .SD(n28571), .Z(debug_rd_3__N_405[29]));
    LUT4 mux_1921_i7_4_lut (.A(n27206), .B(n23522), .C(n27088), .D(n22700), 
         .Z(n3087[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1921_i7_4_lut.init = 16'hca0a;
    PFUMX mux_797_i19 (.BLUT(n36[18]), .ALUT(n1222[18]), .C0(n25706), 
          .Z(pc_23__N_911[18]));
    L6MUX21 i22852 (.D0(n25193), .D1(n25194), .SD(n28571), .Z(debug_rd_3__N_405[30]));
    LUT4 mux_796_i8_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[10] ), 
         .D(addr_out[10]), .Z(n1222[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i9_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[11] ), 
         .D(addr_out[11]), .Z(n1222[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i9_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_797_i18 (.BLUT(n36[17]), .ALUT(n1222[17]), .C0(n25706), 
          .Z(pc_23__N_911[17]));
    LUT4 mux_796_i10_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[12] ), .D(addr_out[12]), .Z(n1222[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i11_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[13] ), .D(addr_out[13]), .Z(n1222[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i11_3_lut_4_lut.init = 16'hf780;
    L6MUX21 i22859 (.D0(n25200), .D1(n25201), .SD(n28571), .Z(debug_rd_3__N_405[31]));
    LUT4 mux_796_i12_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[14] ), .D(addr_out[14]), .Z(n1222[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i12_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_797_i17 (.BLUT(n36[16]), .ALUT(n1222[16]), .C0(n25706), 
          .Z(pc_23__N_911[16]));
    LUT4 i42_4_lut_4_lut (.A(n27211), .B(n28563), .C(n28564), .D(n27209), 
         .Z(n27_adj_2665)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C)))) */ ;
    defparam i42_4_lut_4_lut.init = 16'h404a;
    LUT4 mux_796_i13_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[15] ), .D(addr_out[15]), .Z(n1222[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i14_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[16] ), .D(addr_out[16]), .Z(n1222[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i15_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[17] ), .D(addr_out[17]), .Z(n1222[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1330_i1_3_lut (.A(n33[0]), .B(n1[0]), .C(n2055), .Z(n2056[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1956_i8_3_lut (.A(n3163[7]), .B(n3196[7]), .C(n4073), .Z(n3314[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1956_i8_3_lut.init = 16'hcaca;
    PFUMX mux_797_i16 (.BLUT(n36[15]), .ALUT(n1222[15]), .C0(n25705), 
          .Z(pc_23__N_911[15]));
    LUT4 mux_796_i16_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[18] ), .D(addr_out[18]), .Z(n1222[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i17_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[19] ), .D(addr_out[19]), .Z(n1222[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i18_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[20] ), .D(addr_out[20]), .Z(n1222[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i19_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[21] ), .D(addr_out[21]), .Z(n1222[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i20_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[22] ), .D(addr_out[22]), .Z(n1222[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_796_i21_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[23] ), .D(addr_out[23]), .Z(n1222[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_796_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 i12269_4_lut_4_lut (.A(addr[5]), .B(n44), .C(\data_from_read[2] ), 
         .D(n27294), .Z(data_from_read[0])) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i12269_4_lut_4_lut.init = 16'hf4f0;
    LUT4 i23320_3_lut_4_lut_4_lut (.A(n28562), .B(n23634), .C(n2029), 
         .D(n27198), .Z(n1804[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam i23320_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 i12456_2_lut_rep_472 (.A(instr_fetch_running), .B(debug_early_branch), 
         .Z(n27097)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12456_2_lut_rep_472.init = 16'heeee;
    LUT4 i23458_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n27300), .D(counter_hi[2]), .Z(clk_c_enable_49)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i23458_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i23519_2_lut_rep_665_3_lut (.A(n28573), .B(n28571), .C(counter_hi[2]), 
         .Z(n27290)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i23519_2_lut_rep_665_3_lut.init = 16'h4040;
    LUT4 i23316_3_lut_4_lut_4_lut (.A(n28562), .B(n23624), .C(n2029), 
         .D(n27199), .Z(n1804[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam i23316_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 equal_158_i5_2_lut_rep_671_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(n27296)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam equal_158_i5_2_lut_rep_671_3_lut.init = 16'hfbfb;
    PFUMX mux_797_i15 (.BLUT(n36[14]), .ALUT(n1222[14]), .C0(n25705), 
          .Z(pc_23__N_911[14]));
    LUT4 i23318_3_lut_4_lut_4_lut (.A(n28562), .B(n23614), .C(n2029), 
         .D(n27200), .Z(n1804[2])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam i23318_3_lut_4_lut_4_lut.init = 16'h5c0c;
    PFUMX mux_797_i14 (.BLUT(n36[13]), .ALUT(n1222[13]), .C0(n25705), 
          .Z(pc_23__N_911[13]));
    LUT4 mux_1960_i23_3_lut_4_lut (.A(n4079), .B(n4075), .C(n3350[24]), 
         .D(n24637), .Z(n3350[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1960_i23_3_lut_4_lut.init = 16'hf870;
    PFUMX mux_797_i13 (.BLUT(n36[12]), .ALUT(n1222[12]), .C0(n25705), 
          .Z(pc_23__N_911[12]));
    LUT4 i12465_4_lut (.A(n27204), .B(n28563), .C(n27198), .D(n27209), 
         .Z(n3196[3])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12465_4_lut.init = 16'hc088;
    LUT4 i23472_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n27300), .D(counter_hi[2]), .Z(clk_c_enable_40)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i23472_2_lut_3_lut_4_lut.init = 16'h4000;
    PFUMX mux_797_i12 (.BLUT(n36[11]), .ALUT(n1222[11]), .C0(n25704), 
          .Z(pc_23__N_911[11]));
    PFUMX mux_797_i11 (.BLUT(n36[10]), .ALUT(n1222[10]), .C0(n25704), 
          .Z(pc_23__N_911[10]));
    LUT4 i1_2_lut_rep_728 (.A(instr_len[2]), .B(\pc[2] ), .Z(n27353)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_2_lut_rep_728.init = 16'h6666;
    LUT4 i12464_4_lut (.A(n27203), .B(n28563), .C(n27197), .D(n27209), 
         .Z(n3196[4])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12464_4_lut.init = 16'hc088;
    LUT4 n26435_bdd_3_lut_4_lut (.A(n27131), .B(n27202), .C(n4075), .D(n26435), 
         .Z(n26436)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26435_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i12463_4_lut (.A(n27201), .B(n28563), .C(n27205), .D(n27209), 
         .Z(n3196[5])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12463_4_lut.init = 16'hc088;
    LUT4 i1_2_lut_3_lut_adj_389 (.A(instr_len[2]), .B(\pc[2] ), .C(instr_addr_23__N_318[1]), 
         .Z(n23980)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_2_lut_3_lut_adj_389.init = 16'h9696;
    PFUMX mux_797_i10 (.BLUT(n36[9]), .ALUT(n1222[9]), .C0(n25704), .Z(pc_23__N_911[9]));
    LUT4 mux_1336_i7_3_lut_rep_572 (.A(n2036[6]), .B(n2056[6]), .C(n27260), 
         .Z(n27197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i7_3_lut_rep_572.init = 16'hcaca;
    LUT4 instr_6__I_0_128_i7_2_lut_4_lut (.A(n2036[6]), .B(n2056[6]), .C(n27260), 
         .D(n27198), .Z(n7)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_6__I_0_128_i7_2_lut_4_lut.init = 16'hffca;
    LUT4 i1346_3_lut_rep_635_4_lut_4_lut (.A(instr_len[2]), .B(\pc[2] ), 
         .C(debug_instr_valid), .D(n27354), .Z(n27260)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C (D))+!B !(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1346_3_lut_rep_635_4_lut_4_lut.init = 16'h9c6c;
    LUT4 i3756_2_lut_rep_729 (.A(\pc[1] ), .B(instr_len_c[1]), .Z(n27354)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i3756_2_lut_rep_729.init = 16'h8888;
    LUT4 i2_2_lut_rep_672_3_lut_4_lut (.A(\pc[1] ), .B(instr_len_c[1]), 
         .C(\pc[2] ), .D(instr_len[2]), .Z(n27297)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i2_2_lut_rep_672_3_lut_4_lut.init = 16'h8778;
    PFUMX mux_797_i9 (.BLUT(n36[8]), .ALUT(n1222[8]), .C0(n25704), .Z(pc_23__N_911[8]));
    LUT4 i12501_2_lut_4_lut (.A(n2036[6]), .B(n2056[6]), .C(n27260), .D(n27212), 
         .Z(n2874[4])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12501_2_lut_4_lut.init = 16'hffca;
    LUT4 i3754_2_lut_rep_730 (.A(\pc[1] ), .B(instr_len_c[1]), .Z(n27355)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i3754_2_lut_rep_730.init = 16'h6666;
    LUT4 i12462_4_lut (.A(n27198), .B(n28563), .C(n27201), .D(n27209), 
         .Z(n3196[6])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12462_4_lut.init = 16'hc088;
    LUT4 mux_1326_i2_3_lut (.A(n5[1]), .B(n31[1]), .C(n2035), .Z(n2036[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1326_i2_3_lut.init = 16'hcaca;
    LUT4 i12496_2_lut_2_lut_4_lut (.A(n2036[6]), .B(n2056[6]), .C(n27260), 
         .D(n28563), .Z(n4625[6])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12496_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 n11_bdd_2_lut_4_lut (.A(n2036[6]), .B(n2056[6]), .C(n27260), 
         .D(n27204), .Z(n26028)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam n11_bdd_2_lut_4_lut.init = 16'h00ca;
    PFUMX mux_797_i8 (.BLUT(n36[7]), .ALUT(n1222[7]), .C0(n25703), .Z(pc_23__N_911[7]));
    LUT4 i12401_2_lut_rep_544_4_lut (.A(n2036[6]), .B(n2056[6]), .C(n27260), 
         .D(n27198), .Z(n27169)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12401_2_lut_rep_544_4_lut.init = 16'hca00;
    PFUMX mux_797_i7 (.BLUT(n36[6]), .ALUT(n1222[6]), .C0(n25703), .Z(pc_23__N_911[6]));
    LUT4 instr_6__I_0_129_i7_2_lut_rep_548_4_lut (.A(n2036[6]), .B(n2056[6]), 
         .C(n27260), .D(n27198), .Z(n27173)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_6__I_0_129_i7_2_lut_rep_548_4_lut.init = 16'hcaff;
    LUT4 i22429_3_lut_4_lut (.A(\pc[1] ), .B(instr_len_c[1]), .C(counter_hi[2]), 
         .D(\next_pc_for_core[5] ), .Z(n24772)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i22429_3_lut_4_lut.init = 16'hf606;
    LUT4 i4011_2_lut_rep_664_3_lut (.A(\pc[1] ), .B(instr_len_c[1]), .C(\instr_addr_23__N_318[0] ), 
         .Z(n27289)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i4011_2_lut_rep_664_3_lut.init = 16'hf9f9;
    LUT4 i1_4_lut_4_lut_adj_390 (.A(\pc[1] ), .B(instr_len_c[1]), .C(debug_instr_valid), 
         .D(\instr_addr_23__N_318[0] ), .Z(n8486)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_4_lut_4_lut_adj_390.init = 16'h956a;
    PFUMX mux_797_i6 (.BLUT(n36[5]), .ALUT(n1222[5]), .C0(n25703), .Z(pc_23__N_911[5]));
    LUT4 mux_347_i1_3_lut_4_lut (.A(\pc[1] ), .B(instr_len_c[1]), .C(debug_ret), 
         .D(return_addr[1]), .Z(n1768[0])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam mux_347_i1_3_lut_4_lut.init = 16'hf606;
    PFUMX mux_797_i5 (.BLUT(n36[4]), .ALUT(n1222[4]), .C0(n25703), .Z(pc_23__N_911[4]));
    PFUMX pc_23__I_0_450_i209_rep_69 (.BLUT(n149_adj_2643), .ALUT(n225), 
          .C0(n28571), .Z(n24612)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    PFUMX mux_797_i4 (.BLUT(n36[3]), .ALUT(n1222[3]), .C0(n25702), .Z(pc_23__N_911[3]));
    PFUMX mux_797_i3 (.BLUT(n36[2]), .ALUT(n1222[2]), .C0(n25702), .Z(pc_23__N_911[2]));
    PFUMX mux_797_i2 (.BLUT(n36[1]), .ALUT(n1222[1]), .C0(n25702), .Z(pc_23__N_911[1]));
    LUT4 mux_1933_i7_4_lut (.A(n2133[0]), .B(n27198), .C(n4065), .D(n27212), 
         .Z(n3163[6])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1933_i7_4_lut.init = 16'hfaca;
    LUT4 i1_3_lut_adj_391 (.A(mie[14]), .B(n18144), .C(n8_adj_2666), .Z(n926)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_391.init = 16'hcece;
    LUT4 mux_1336_i6_3_lut_rep_573 (.A(n2036[5]), .B(n2056[5]), .C(n27260), 
         .Z(n27198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i6_3_lut_rep_573.init = 16'hcaca;
    PFUMX mux_797_i1 (.BLUT(n36[0]), .ALUT(n1222[0]), .C0(n25702), .Z(pc_23__N_911[0]));
    LUT4 i12460_4_lut (.A(n27197), .B(n28563), .C(n27199), .D(n27209), 
         .Z(n3196[7])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12460_4_lut.init = 16'hc088;
    LUT4 i20040_3_lut_rep_501 (.A(n10), .B(addr[26]), .C(addr[27]), .Z(n27126)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i20040_3_lut_rep_501.init = 16'heaea;
    LUT4 i22492_2_lut_rep_737 (.A(counter_hi[4]), .B(counter_hi[3]), .Z(n27362)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i22492_2_lut_rep_737.init = 16'h4444;
    LUT4 i22479_2_lut_3_lut (.A(counter_hi[4]), .B(n28573), .C(alu_a_in_3__N_1552), 
         .Z(n24822)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i22479_2_lut_3_lut.init = 16'h4040;
    LUT4 i243_2_lut_4_lut (.A(n10), .B(addr[26]), .C(addr[27]), .D(load_started), 
         .Z(n824)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B !(D)))) */ ;
    defparam i243_2_lut_4_lut.init = 16'h1500;
    LUT4 i1_3_lut_adj_392 (.A(mie[10]), .B(n18144), .C(n8_adj_2666), .Z(n893)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_392.init = 16'hcece;
    LUT4 pc_23__I_0_450_i269_rep_68_3_lut_4_lut (.A(counter_hi[4]), .B(counter_hi[3]), 
         .C(n24612), .D(n157), .Z(n24611)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam pc_23__I_0_450_i269_rep_68_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_3_lut_adj_393 (.A(mie[6]), .B(n18144), .C(n8_adj_2666), .Z(n860)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_393.init = 16'hcece;
    LUT4 i1_2_lut_4_lut_adj_394 (.A(n2036[5]), .B(n2056[5]), .C(n27260), 
         .D(n27200), .Z(n22164)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_394.init = 16'h00ca;
    LUT4 mux_1975_i9_4_lut (.A(n3273[8]), .B(instr[28]), .C(n4079), .D(n8123), 
         .Z(n3397[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1975_i9_4_lut.init = 16'hca0a;
    LUT4 i1_3_lut_adj_395 (.A(mie[2]), .B(n18144), .C(n8_adj_2666), .Z(n793)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_395.init = 16'hcece;
    LUT4 i23637_4_lut (.A(n27114), .B(n27112), .C(n8274), .D(is_ret_de), 
         .Z(debug_instr_valid_N_436)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i23637_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_396 (.A(n2326), .B(n27092), .C(n27207), .D(n4_adj_2638), 
         .Z(n22748)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;
    defparam i1_4_lut_adj_396.init = 16'h20a0;
    LUT4 i23695_3_lut_4_lut (.A(n4057), .B(n27260), .C(n27101), .D(n4075), 
         .Z(n25004)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i23695_3_lut_4_lut.init = 16'hff1f;
    LUT4 mux_1336_i4_3_lut_rep_574 (.A(n2036[3]), .B(n2056[3]), .C(n27260), 
         .Z(n27199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i4_3_lut_rep_574.init = 16'hcaca;
    LUT4 mux_1330_i2_3_lut (.A(n33[1]), .B(n1[1]), .C(n2055), .Z(n2056[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1330_i2_3_lut.init = 16'hcaca;
    LUT4 instr_6__I_0_128_i6_2_lut_rep_549_4_lut (.A(n2036[3]), .B(n2056[3]), 
         .C(n27260), .D(n27201), .Z(n27174)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_6__I_0_128_i6_2_lut_rep_549_4_lut.init = 16'hffca;
    LUT4 n26178_bdd_3_lut (.A(n26178), .B(n26175), .C(n28571), .Z(debug_branch_N_442[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26178_bdd_3_lut.init = 16'hcaca;
    LUT4 i12504_2_lut_4_lut (.A(n2036[3]), .B(n2056[3]), .C(n27260), .D(n27212), 
         .Z(n2874[7])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12504_2_lut_4_lut.init = 16'hffca;
    LUT4 is_jalr_N_1372_bdd_2_lut_23816_4_lut (.A(n27171), .B(n27142), .C(n28563), 
         .D(n27129), .Z(n26206)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam is_jalr_N_1372_bdd_2_lut_23816_4_lut.init = 16'h0002;
    LUT4 i22225_2_lut_rep_551_4_lut (.A(n2036[3]), .B(n2056[3]), .C(n27260), 
         .D(n27200), .Z(n27176)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i22225_2_lut_rep_551_4_lut.init = 16'hffca;
    LUT4 i1_3_lut_rep_468_4_lut (.A(instr_fetch_running), .B(debug_early_branch), 
         .C(instr_fetch_restart_N_947), .D(n22592), .Z(n27093)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_rep_468_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_4_lut_adj_397 (.A(n2036[3]), .B(n2056[3]), .C(n27260), 
         .D(n28564), .Z(n23470)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_397.init = 16'h00ca;
    LUT4 i23525_4_lut (.A(n27114), .B(n22592), .C(n27277), .D(n23580), 
         .Z(clk_c_enable_115)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i23525_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_547_4_lut (.A(n2036[3]), .B(n2056[3]), .C(n27260), 
         .D(n27201), .Z(n27172)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_547_4_lut.init = 16'hcaff;
    LUT4 i23514_4_lut (.A(n27114), .B(rst_reg_n), .C(n22592), .D(n23526), 
         .Z(clk_c_enable_117)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i23514_4_lut.init = 16'h3337;
    LUT4 i1_2_lut_rep_497_4_lut (.A(n27171), .B(n27142), .C(n28563), .D(n27185), 
         .Z(n27122)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_497_4_lut.init = 16'h0200;
    LUT4 i23522_4_lut (.A(n27114), .B(n22592), .C(n27277), .D(n23572), 
         .Z(clk_c_enable_142)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i23522_4_lut.init = 16'h0010;
    LUT4 i1_3_lut_4_lut_adj_398 (.A(instr_fetch_running), .B(debug_early_branch), 
         .C(instr_fetch_restart_N_947), .D(n22592), .Z(n22591)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_adj_398.init = 16'hffef;
    LUT4 mux_1960_i22_3_lut_4_lut (.A(n4079), .B(n4075), .C(n3350[24]), 
         .D(n24631), .Z(n3350[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1960_i22_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_1336_i5_3_lut_rep_575 (.A(n2036[4]), .B(n2056[4]), .C(n27260), 
         .Z(n27200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i5_3_lut_rep_575.init = 16'hcaca;
    LUT4 mux_1956_i5_3_lut (.A(n3163[4]), .B(n3196[4]), .C(n4073), .Z(n3314[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1956_i5_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_399 (.A(n27205), .B(rst_reg_n), .C(n27207), .D(n27211), 
         .Z(n23792)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_399.init = 16'hc088;
    LUT4 i1_2_lut_4_lut_adj_400 (.A(n2036[4]), .B(n2056[4]), .C(n27260), 
         .D(n28564), .Z(n23462)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_400.init = 16'h00ca;
    LUT4 i1_2_lut_rep_545_4_lut (.A(n2036[4]), .B(n2056[4]), .C(n27260), 
         .D(n27201), .Z(n27170)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_545_4_lut.init = 16'hffca;
    LUT4 i1_4_lut_adj_401 (.A(\imm[1] ), .B(n27330), .C(n24398), .D(\imm[2] ), 
         .Z(n24404)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_401.init = 16'h0010;
    LUT4 mux_1336_i3_3_lut_rep_576 (.A(n2036[2]), .B(n2056[2]), .C(n27260), 
         .Z(n27201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i3_3_lut_rep_576.init = 16'hcaca;
    LUT4 n11_bdd_2_lut_23725_2_lut_4_lut (.A(n2036[2]), .B(n2056[2]), .C(n27260), 
         .D(n27211), .Z(n26027)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam n11_bdd_2_lut_23725_2_lut_4_lut.init = 16'h00ca;
    L6MUX21 shift_right_317_i272 (.D0(n212), .D1(n9117), .SD(counter_hi[4]), 
            .Z(debug_branch_N_840[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i1_2_lut_rep_741 (.A(alu_op[1]), .B(alu_op[0]), .Z(n27366)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_rep_741.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_402 (.A(n2036[2]), .B(n2056[2]), .C(n27260), 
         .D(n28564), .Z(n23478)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_402.init = 16'h00ca;
    LUT4 i1_3_lut_rep_680_4_lut (.A(alu_op[1]), .B(alu_op[0]), .C(n27368), 
         .D(alu_op[2]), .Z(n27305)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_rep_680_4_lut.init = 16'h0010;
    LUT4 is_system_I_0_481_2_lut_rep_743 (.A(is_system), .B(debug_instr_valid), 
         .Z(n27368)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam is_system_I_0_481_2_lut_rep_743.init = 16'h8888;
    LUT4 i1_2_lut_rep_650_3_lut_2_lut_3_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[1]), .Z(n27275)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_650_3_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_624_3_lut_4_lut_3_lut_4_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[0]), .D(alu_op[1]), .Z(n27249)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_624_3_lut_4_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_623_3_lut_4_lut_3_lut_4_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[0]), .D(alu_op[1]), .Z(n27248)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_623_3_lut_4_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 is_system_I_0_2_lut_rep_742_4_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[0]), .D(alu_op[1]), .Z(n27367)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam is_system_I_0_2_lut_rep_742_4_lut.init = 16'h8880;
    LUT4 i23588_2_lut_rep_744 (.A(alu_op[1]), .B(alu_op[0]), .Z(n27369)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i23588_2_lut_rep_744.init = 16'h4444;
    LUT4 i1_2_lut_rep_677_3_lut_4_lut (.A(alu_op[1]), .B(alu_op[0]), .C(cycle[0]), 
         .D(cycle[1]), .Z(n27302)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_rep_677_3_lut_4_lut.init = 16'hffbf;
    LUT4 mux_1336_i9_3_lut_rep_577 (.A(n2036[8]), .B(n2056[8]), .C(n27260), 
         .Z(n27202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i9_3_lut_rep_577.init = 16'hcaca;
    LUT4 i1_4_lut_then_4_lut (.A(n27166), .B(n2056[3]), .C(n23658), .D(n27201), 
         .Z(n27390)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h4010;
    LUT4 i12623_2_lut_2_lut_4_lut (.A(n2036[8]), .B(n2056[8]), .C(n27260), 
         .D(n27095), .Z(n2342[1])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12623_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 i12621_2_lut_4_lut (.A(n2036[8]), .B(n2056[8]), .C(n27260), .D(n2322), 
         .Z(n2128[1])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12621_2_lut_4_lut.init = 16'hffca;
    LUT4 i12646_2_lut_2_lut_4_lut (.A(n2036[8]), .B(n2056[8]), .C(n27260), 
         .D(n27209), .Z(n2347[1])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12646_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_1336_i12_3_lut_rep_578 (.A(n2036[11]), .B(n2056[11]), .C(n27260), 
         .Z(n27203)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i12_3_lut_rep_578.init = 16'hcaca;
    LUT4 i1_4_lut_adj_403 (.A(\imm[10] ), .B(imm[0]), .C(n27374), .D(\imm[6] ), 
         .Z(n24398)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_403.init = 16'h4000;
    LUT4 i23533_2_lut_rep_561_4_lut (.A(n2036[11]), .B(n2056[11]), .C(n27260), 
         .D(n27204), .Z(n27186)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i23533_2_lut_rep_561_4_lut.init = 16'h35ff;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(alu_op[1]), .B(alu_op[0]), .C(data_rs1[3]), 
         .D(n27367), .Z(n8_adj_2668)) /* synthesis lut_function=(A (C (D))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'he400;
    PFUMX shift_right_317_i212 (.BLUT(n24780), .ALUT(n9091), .C0(counter_hi[3]), 
          .Z(n212)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 mux_1960_i21_3_lut_4_lut (.A(n4079), .B(n4075), .C(n3350[24]), 
         .D(n24629), .Z(n3350[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1960_i21_3_lut_4_lut.init = 16'hf870;
    LUT4 i12494_2_lut_2_lut_4_lut (.A(n2036[11]), .B(n2056[11]), .C(n27260), 
         .D(n28563), .Z(n4625[3])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12494_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_1336_i11_3_lut_rep_579 (.A(n2036[10]), .B(n2056[10]), .C(n27260), 
         .Z(n27204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i11_3_lut_rep_579.init = 16'hcaca;
    LUT4 i12498_2_lut_4_lut (.A(n2036[10]), .B(n2056[10]), .C(n27260), 
         .D(n28563), .Z(n4625[8])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12498_2_lut_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_467_3_lut_4_lut (.A(n27103), .B(n27109), .C(n27179), 
         .D(rst_reg_n), .Z(n27092)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i1_2_lut_rep_467_3_lut_4_lut.init = 16'h0200;
    LUT4 i3722_2_lut_rep_746 (.A(rd[1]), .B(rd[0]), .Z(n27371)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(180[19:31])
    defparam i3722_2_lut_rep_746.init = 16'h8888;
    LUT4 i3729_2_lut_3_lut (.A(rd[1]), .B(rd[0]), .C(rd[2]), .Z(n5868)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(180[19:31])
    defparam i3729_2_lut_3_lut.init = 16'h8080;
    LUT4 i3685_2_lut_rep_747 (.A(rs2[0]), .B(mem_op_increment_reg), .Z(n27372)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i3685_2_lut_rep_747.init = 16'h8888;
    LUT4 i12625_2_lut_2_lut_4_lut (.A(n2036[10]), .B(n2056[10]), .C(n27260), 
         .D(n27095), .Z(n2342[3])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12625_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 i12648_2_lut_2_lut_4_lut (.A(n2036[10]), .B(n2056[10]), .C(n27260), 
         .D(n27209), .Z(n2347[3])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12648_2_lut_2_lut_4_lut.init = 16'hcaff;
    LUT4 mux_1336_i13_3_lut_rep_580 (.A(n2036[12]), .B(n2056[12]), .C(n27260), 
         .Z(n27205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i13_3_lut_rep_580.init = 16'hcaca;
    LUT4 i3693_2_lut_rep_679_3_lut (.A(rs2[0]), .B(mem_op_increment_reg), 
         .C(rs2[1]), .Z(n27304)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i3693_2_lut_rep_679_3_lut.init = 16'h8080;
    LUT4 i3700_2_lut_3_lut_4_lut (.A(rs2[0]), .B(mem_op_increment_reg), 
         .C(rs2[2]), .D(rs2[1]), .Z(n5839)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i3700_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 equal_25_i3_2_lut_4_lut (.A(n2036[12]), .B(n2056[12]), .C(n27260), 
         .D(n27211), .Z(n3)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam equal_25_i3_2_lut_4_lut.init = 16'hff35;
    LUT4 mux_1336_i8_3_lut_rep_581 (.A(n2036[7]), .B(n2056[7]), .C(n27260), 
         .Z(n27206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i8_3_lut_rep_581.init = 16'hcaca;
    LUT4 i1_4_lut_adj_404 (.A(n27112), .B(n27109), .C(n27106), .D(n23662), 
         .Z(n4075)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_404.init = 16'h1000;
    LUT4 i12290_2_lut_4_lut (.A(n2036[7]), .B(n2056[7]), .C(n27260), .D(n27095), 
         .Z(n2342[0])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12290_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_1077_i11_3_lut (.A(n1[10]), .B(n5[10]), .C(n2055), .Z(n1735[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i11_3_lut.init = 16'hcaca;
    LUT4 i12313_2_lut_4_lut (.A(n2036[7]), .B(n2056[7]), .C(n27260), .D(n27209), 
         .Z(n2347[0])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12313_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_rep_552_4_lut (.A(n2036[7]), .B(n2056[7]), .C(n27260), 
         .D(n27207), .Z(n27177)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_552_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_rep_749 (.A(\imm[9] ), .B(\imm[8] ), .Z(n27374)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_rep_749.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_405 (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[31]), 
         .D(n27305), .Z(addr_out[27])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_3_lut_4_lut_adj_405.init = 16'h70f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_406 (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[29]), 
         .D(n27305), .Z(addr_out[25])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_3_lut_4_lut_adj_406.init = 16'h70f0;
    LUT4 i1_3_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(\imm[4] ), 
         .D(\imm[10] ), .Z(n22088)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_407 (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[30]), 
         .D(n27305), .Z(addr_out[26])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_3_lut_4_lut_adj_407.init = 16'h70f0;
    LUT4 i12212_2_lut_4_lut (.A(n2036[7]), .B(n2056[7]), .C(n27260), .D(n28563), 
         .Z(n2133[0])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12212_2_lut_4_lut.init = 16'h00ca;
    LUT4 i12578_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[28]), 
         .D(n27305), .Z(addr_out[24])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i12578_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 mux_1336_i10_3_lut_rep_582 (.A(n2036[9]), .B(n2056[9]), .C(n27260), 
         .Z(n27207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i10_3_lut_rep_582.init = 16'hcaca;
    LUT4 i12497_2_lut_4_lut (.A(n2036[9]), .B(n2056[9]), .C(n27260), .D(n28563), 
         .Z(n4625[7])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12497_2_lut_4_lut.init = 16'h00ca;
    LUT4 i12647_2_lut_2_lut_4_lut (.A(n2036[9]), .B(n2056[9]), .C(n27260), 
         .D(n27209), .Z(n2347[2])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12647_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 i12624_2_lut_2_lut_4_lut (.A(n2036[9]), .B(n2056[9]), .C(n27260), 
         .D(n27095), .Z(n2342[2])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12624_2_lut_2_lut_4_lut.init = 16'h00ca;
    PFUMX i22431 (.BLUT(n24773), .ALUT(n226), .C0(counter_hi[4]), .Z(n24774));
    LUT4 mux_1975_i16_3_lut (.A(n3163[14]), .B(n3314[15]), .C(n24959), 
         .Z(n3397[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1975_i16_3_lut.init = 16'hcaca;
    LUT4 i23594_2_lut_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), .D(n27209), 
         .Z(n25126)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i23594_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_1975_i15_3_lut (.A(n3163[14]), .B(n3314[14]), .C(n24959), 
         .Z(n3397[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1975_i15_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_560_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n27209), .Z(n27185)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i2_2_lut_rep_560_4_lut.init = 16'h3500;
    LUT4 mux_1336_i1_3_lut_rep_760 (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .Z(n28564)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i1_3_lut_rep_760.init = 16'hcaca;
    LUT4 i23491_2_lut_rep_534_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n27212), .Z(n27159)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i23491_2_lut_rep_534_4_lut.init = 16'h0035;
    LUT4 mux_1975_i14_3_lut (.A(n3163[14]), .B(n3314[13]), .C(n24959), 
         .Z(n3397[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1975_i14_3_lut.init = 16'hcaca;
    LUT4 i22248_2_lut_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), .D(n27209), 
         .Z(n24525)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i22248_2_lut_4_lut.init = 16'hffca;
    LUT4 n28140_bdd_2_lut_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n28140), .Z(n28141)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam n28140_bdd_2_lut_4_lut.init = 16'h3500;
    PFUMX i23947 (.BLUT(n26434), .ALUT(n26433), .C0(n27101), .Z(n26435));
    LUT4 i3767_4_lut_4_lut (.A(\pc[2] ), .B(instr_len[2]), .C(\pc[1] ), 
         .D(instr_len_c[1]), .Z(next_pc_offset[3])) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i3767_4_lut_4_lut.init = 16'he888;
    LUT4 mux_1938_i12_3_lut_4_lut (.A(n4075), .B(n27101), .C(n4745[4]), 
         .D(n24629), .Z(n3232[11])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1938_i12_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i2_2_lut_rep_539_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n27211), .Z(n27164)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i2_2_lut_rep_539_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_rep_550_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n27212), .Z(n27175)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_550_4_lut.init = 16'h3500;
    LUT4 mux_1975_i13_3_lut (.A(n3163[14]), .B(n3314[12]), .C(n24959), 
         .Z(n3397[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1975_i13_3_lut.init = 16'hcaca;
    PFUMX next_pc_for_core_23__I_0_i209 (.BLUT(n149), .ALUT(n225_adj_2669), 
          .C0(counter_hi[4]), .Z(n209)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i166_2_lut_rep_564_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n27209), .Z(n27189)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i166_2_lut_rep_564_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_751 (.A(n28573), .B(n28571), .Z(n27376)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_2_lut_rep_751.init = 16'heeee;
    LUT4 i23498_4_lut (.A(n27114), .B(rst_reg_n), .C(n22592), .D(n23532), 
         .Z(clk_c_enable_144)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i23498_4_lut.init = 16'h3337;
    LUT4 mux_1975_i11_4_lut (.A(n2874[9]), .B(instr[30]), .C(n4079), .D(n8123), 
         .Z(n3397[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1975_i11_4_lut.init = 16'hca0a;
    LUT4 mux_1975_i10_4_lut (.A(n26348), .B(instr[29]), .C(n4079), .D(n8123), 
         .Z(n3397[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1975_i10_4_lut.init = 16'hca0a;
    LUT4 i1_3_lut_4_lut_adj_408 (.A(counter_hi[3]), .B(counter_hi[4]), .C(timer_interrupt), 
         .D(counter_hi[2]), .Z(csr_read_3__N_1459[3])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_3_lut_4_lut_adj_408.init = 16'h1000;
    LUT4 i1_2_lut_rep_558_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n27212), .Z(n27183)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_558_4_lut.init = 16'hca00;
    LUT4 i23646_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_top_bit_next_N_1731), .D(counter_hi[2]), .Z(n15206)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i23646_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i3424_2_lut_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(mstatus_mte), .D(counter_hi[2]), .Z(n5434)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i3424_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    L6MUX21 i22894 (.D0(n25233), .D1(n25234), .SD(n28573), .Z(n25237));
    LUT4 i1_2_lut_rep_681_3_lut (.A(n28573), .B(n28571), .C(counter_hi[2]), 
         .Z(n27306)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_2_lut_rep_681_3_lut.init = 16'hfefe;
    LUT4 i10821_1_lut_rep_633_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(clk_c_enable_71)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i10821_1_lut_rep_633_2_lut_3_lut.init = 16'h0101;
    PFUMX i22401 (.BLUT(n24742), .ALUT(n24743), .C0(counter_hi[2]), .Z(n24744));
    LUT4 i1_2_lut_rep_554_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n27209), .Z(n27179)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_554_4_lut.init = 16'hca00;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_top_bit_next_N_1731), .D(counter_hi[2]), .Z(clk_c_enable_422)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i12429_2_lut_rep_620_2_lut_3_lut_4_lut (.A(n28573), .B(n28571), 
         .C(cy), .D(counter_hi[2]), .Z(n27245)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i12429_2_lut_rep_620_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i23508_4_lut (.A(n27114), .B(n22592), .C(n27277), .D(n23564), 
         .Z(clk_c_enable_158)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i23508_4_lut.init = 16'h0010;
    LUT4 equal_3217_i8_2_lut_rep_684_3_lut (.A(n28573), .B(n28571), .C(counter_hi[2]), 
         .Z(n27309)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam equal_3217_i8_2_lut_rep_684_3_lut.init = 16'hefef;
    LUT4 i23477_4_lut (.A(n27114), .B(rst_reg_n), .C(n22592), .D(n23536), 
         .Z(clk_c_enable_160)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i23477_4_lut.init = 16'h3337;
    LUT4 i12542_2_lut_3_lut_4_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(csr_read_3__N_1443[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i12542_2_lut_3_lut_4_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_752 (.A(alu_op[3]), .B(tmp_data[31]), .Z(n27377)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_rep_752.init = 16'h8888;
    LUT4 i4963_3_lut_4_lut (.A(alu_op[3]), .B(tmp_data[31]), .C(shift_amt[5]), 
         .D(n7278), .Z(shift_out[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i4963_3_lut_4_lut.init = 16'h8f80;
    LUT4 i22949_3_lut_4_lut (.A(alu_op[3]), .B(tmp_data[31]), .C(shift_amt[1]), 
         .D(n62), .Z(n25292)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i22949_3_lut_4_lut.init = 16'h8f80;
    LUT4 i5836_3_lut_4_lut (.A(alu_op[3]), .B(tmp_data[31]), .C(shift_amt[5]), 
         .D(n8153), .Z(shift_out[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i5836_3_lut_4_lut.init = 16'h8f80;
    LUT4 n192_bdd_3_lut_24077_4_lut (.A(alu_op[3]), .B(tmp_data[31]), .C(shift_amt[5]), 
         .D(n8157), .Z(n26049)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam n192_bdd_3_lut_24077_4_lut.init = 16'h8f80;
    LUT4 n26685_bdd_3_lut_4_lut (.A(alu_op[3]), .B(tmp_data[31]), .C(shift_amt[5]), 
         .D(n26685), .Z(n26686)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam n26685_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i22781_2_lut_rep_542_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n27209), .Z(n27167)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i22781_2_lut_rep_542_4_lut.init = 16'h00ca;
    LUT4 top_bit_I_0_i63_3_lut_4_lut (.A(alu_op[3]), .B(tmp_data[31]), .C(shift_amt[0]), 
         .D(a_for_shift_right[31]), .Z(n63)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam top_bit_I_0_i63_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_4_lut_adj_409 (.A(n27114), .B(n22592), .C(n27277), .D(n23558), 
         .Z(clk_c_enable_174)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(410[18] 430[16])
    defparam i1_4_lut_adj_409.init = 16'h1000;
    LUT4 i1_4_lut_adj_410 (.A(n4116[2]), .B(n4116[1]), .C(n4116[0]), .D(n27109), 
         .Z(additional_mem_ops_2__N_749[2])) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_410.init = 16'ha9aa;
    LUT4 i12332_1_lut_rep_522_2_lut_4_lut (.A(n2036[0]), .B(n2056[0]), .C(n27260), 
         .D(n27209), .Z(n27147)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12332_1_lut_rep_522_2_lut_4_lut.init = 16'h35ff;
    LUT4 mux_1336_i2_3_lut_rep_584 (.A(n2036[1]), .B(n2056[1]), .C(n27260), 
         .Z(n27209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i2_3_lut_rep_584.init = 16'hcaca;
    LUT4 i23591_2_lut_rep_535_4_lut (.A(n2036[1]), .B(n2056[1]), .C(n27260), 
         .D(n27211), .Z(n27160)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i23591_2_lut_rep_535_4_lut.init = 16'h0035;
    PFUMX i22890 (.BLUT(\mem_data_from_read[1] ), .ALUT(\mem_data_from_read[5] ), 
          .C0(counter_hi[2]), .Z(n25233));
    LUT4 n26805_bdd_2_lut_4_lut (.A(n2036[1]), .B(n2056[1]), .C(n27260), 
         .D(n26805), .Z(n26806)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam n26805_bdd_2_lut_4_lut.init = 16'h3500;
    LUT4 pc_3__bdd_3_lut_23800 (.A(\pc[7] ), .B(\pc[15] ), .C(counter_hi[3]), 
         .Z(n26176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_3__bdd_3_lut_23800.init = 16'hcaca;
    LUT4 i23578_2_lut_rep_543_4_lut (.A(n2036[1]), .B(n2056[1]), .C(n27260), 
         .D(n28563), .Z(n27168)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i23578_2_lut_rep_543_4_lut.init = 16'h3500;
    LUT4 i23686_2_lut_4_lut (.A(n2036[1]), .B(n2056[1]), .C(n27260), .D(n27212), 
         .Z(n25014)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i23686_2_lut_4_lut.init = 16'hcaff;
    PFUMX i38 (.BLUT(n17), .ALUT(n22_adj_2664), .C0(n27212), .Z(n24_adj_2670));
    LUT4 pc_3__bdd_3_lut_23882 (.A(\pc[3] ), .B(\pc[11] ), .C(counter_hi[3]), 
         .Z(n26177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_3__bdd_3_lut_23882.init = 16'hcaca;
    PFUMX i22891 (.BLUT(\mem_data_from_read[9] ), .ALUT(\mem_data_from_read[13] ), 
          .C0(counter_hi[2]), .Z(n25234));
    PFUMX debug_branch_I_48_i3 (.BLUT(n9115), .ALUT(debug_branch_N_840[30]), 
          .C0(n25057), .Z(debug_branch_N_450[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i12337_2_lut (.A(n26029), .B(n4071), .Z(n3273[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12337_2_lut.init = 16'h8888;
    LUT4 mem_data_from_read_6__bdd_4_lut (.A(counter_hi[3]), .B(\data_from_read[6] ), 
         .C(\data_from_read[2] ), .D(counter_hi[2]), .Z(n26712)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mem_data_from_read_6__bdd_4_lut.init = 16'he4f0;
    LUT4 i17737_2_lut (.A(counter_hi[3]), .B(counter_hi[2]), .Z(n34[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i17737_2_lut.init = 16'h6666;
    PFUMX debug_branch_I_48_i1 (.BLUT(n9111), .ALUT(debug_branch_N_840[28]), 
          .C0(n25057), .Z(debug_branch_N_450[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 mux_1073_i11_rep_99_3_lut (.A(n31[10]), .B(n33[10]), .C(n2035), 
         .Z(n24642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i11_rep_99_3_lut.init = 16'hcaca;
    LUT4 mux_1336_i14_3_lut_rep_586 (.A(n2036[13]), .B(n2056[13]), .C(n27260), 
         .Z(n27211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i14_3_lut_rep_586.init = 16'hcaca;
    LUT4 n26715_bdd_3_lut_24396 (.A(n26715), .B(n27401), .C(counter_hi[3]), 
         .Z(n26716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26715_bdd_3_lut_24396.init = 16'hcaca;
    LUT4 i1_4_lut_adj_411 (.A(n22369), .B(n22816), .C(instr_fetch_running_N_945), 
         .D(instr_fetch_stopped), .Z(clk_c_enable_209)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_411.init = 16'hfffd;
    LUT4 i12172_4_lut (.A(instr_fetch_running_N_943), .B(rst_reg_n), .C(was_early_branch), 
         .D(n27114), .Z(n5590)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam i12172_4_lut.init = 16'hc088;
    LUT4 i12162_4_lut (.A(instr_fetch_running_N_945), .B(n27108), .C(n8), 
         .D(n23602), .Z(instr_fetch_running_N_943)) /* synthesis lut_function=(A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam i12162_4_lut.init = 16'ha2aa;
    LUT4 i1_3_lut_adj_412 (.A(is_jal_de), .B(rst_reg_n), .C(is_ret_de), 
         .Z(n23600)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut_adj_412.init = 16'hc8c8;
    LUT4 instr_addr_23__I_0_i2_3_lut (.A(instr_addr_23__N_318[1]), .B(\early_branch_addr[2] ), 
         .C(was_early_branch), .Z(\instr_addr[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[25:119])
    defparam instr_addr_23__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_2_lut_rep_567_4_lut (.A(n2036[13]), .B(n2056[13]), .C(n27260), 
         .D(n28563), .Z(n27192)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_2_lut_rep_567_4_lut.init = 16'h3500;
    LUT4 i1_4_lut_adj_413 (.A(n27226), .B(n27126), .C(data_ready_sync), 
         .D(clk_c_enable_276), .Z(clk_c_enable_278)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_413.init = 16'hfbbb;
    LUT4 i1_2_lut_rep_546_4_lut (.A(n2036[13]), .B(n2056[13]), .C(n27260), 
         .D(n27212), .Z(n27171)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_546_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_rep_565_4_lut (.A(n2036[13]), .B(n2056[13]), .C(n27260), 
         .D(n27212), .Z(n27190)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_565_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_537_4_lut (.A(n2036[13]), .B(n2056[13]), .C(n27260), 
         .D(n28563), .Z(n27162)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_537_4_lut.init = 16'hca00;
    LUT4 i1_2_lut_rep_553_4_lut (.A(n2036[13]), .B(n2056[13]), .C(n27260), 
         .D(n28563), .Z(n27178)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_553_4_lut.init = 16'hffca;
    LUT4 mux_1336_i16_3_lut_rep_587 (.A(n2036[15]), .B(n2056[15]), .C(n27260), 
         .Z(n27212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1336_i16_3_lut_rep_587.init = 16'hcaca;
    LUT4 pc_2__bdd_3_lut_23808 (.A(\pc[6] ), .B(\pc[14] ), .C(counter_hi[3]), 
         .Z(n26196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_2__bdd_3_lut_23808.init = 16'hcaca;
    PFUMX i6777 (.BLUT(n24758), .ALUT(n24759), .C0(n27268), .Z(n9117));
    PFUMX i54 (.BLUT(n37), .ALUT(n32), .C0(n25014), .Z(n35));
    LUT4 n26198_bdd_3_lut (.A(n26198), .B(n26195), .C(n28571), .Z(debug_branch_N_442[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26198_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_414 (.A(n2036[15]), .B(n2056[15]), .C(n27260), 
         .D(n28575), .Z(n23588)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_414.init = 16'hca00;
    PFUMX i23899 (.BLUT(n26347), .ALUT(n26346), .C0(n4071), .Z(n26348));
    LUT4 i12287_2_lut_rep_538_4_lut (.A(n2036[15]), .B(n2056[15]), .C(n27260), 
         .D(n28563), .Z(n27163)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i12287_2_lut_rep_538_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_rep_559_4_lut (.A(n2036[15]), .B(n2056[15]), .C(n27260), 
         .D(n28563), .Z(n27184)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_559_4_lut.init = 16'hca00;
    LUT4 i22232_4_lut (.A(n27102), .B(addr_offset[3]), .C(n27109), .D(addr_offset[2]), 
         .Z(n24509)) /* synthesis lut_function=(!((B (C (D))+!B !(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i22232_4_lut.init = 16'h2888;
    LUT4 additional_mem_ops_2__N_1132_0__bdd_2_lut_4_lut (.A(n2036[14]), .B(n2056[14]), 
         .C(n27260), .D(n27121), .Z(n26745)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam additional_mem_ops_2__N_1132_0__bdd_2_lut_4_lut.init = 16'h00ca;
    LUT4 i1_4_lut_else_4_lut (.A(n27166), .B(n2036[3]), .C(n23658), .D(n27201), 
         .Z(n27389)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4010;
    LUT4 mem_data_from_read_4__bdd_4_lut (.A(counter_hi[3]), .B(data_from_read[0]), 
         .C(\data_from_read[2] ), .D(counter_hi[2]), .Z(n26728)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam mem_data_from_read_4__bdd_4_lut.init = 16'hf0e4;
    PFUMX i42 (.BLUT(n10_adj_2671), .ALUT(n29), .C0(n28564), .Z(n23));
    LUT4 i1_4_lut_adj_415 (.A(n24599), .B(n24210), .C(n23140), .D(addr[6]), 
         .Z(is_timer_addr)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_415.init = 16'h0040;
    LUT4 i22319_3_lut (.A(addr[3]), .B(addr[5]), .C(addr[4]), .Z(n24599)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22319_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_416 (.A(addr[7]), .B(n24198), .C(n24202), .D(n24200), 
         .Z(n24210)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_416.init = 16'h4000;
    LUT4 i1_4_lut_adj_417 (.A(addr[24]), .B(n24182), .C(n24174), .D(addr[27]), 
         .Z(n23140)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_417.init = 16'h8000;
    PFUMX i22403 (.BLUT(\mem_data_from_read[24] ), .ALUT(\mem_data_from_read[28] ), 
          .C0(counter_hi[2]), .Z(n24746));
    LUT4 pc_1__bdd_3_lut_23812 (.A(\pc[5] ), .B(\pc[13] ), .C(counter_hi[3]), 
         .Z(n26201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_1__bdd_3_lut_23812.init = 16'hcaca;
    LUT4 n26731_bdd_3_lut (.A(n26731), .B(n27397), .C(counter_hi[3]), 
         .Z(n26732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26731_bdd_3_lut.init = 16'hcaca;
    PFUMX i22409 (.BLUT(\mem_data_from_read[26] ), .ALUT(\mem_data_from_read[30] ), 
          .C0(counter_hi[2]), .Z(n24752));
    LUT4 no_write_in_progress_I_42_4_lut (.A(n24126), .B(addr_out[27]), 
         .C(n27244), .D(n27126), .Z(no_write_in_progress_N_471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(279[18] 289[12])
    defparam no_write_in_progress_I_42_4_lut.init = 16'hcacf;
    LUT4 i1_4_lut_adj_418 (.A(n27205), .B(n28575), .C(n27202), .D(n27211), 
         .Z(n23756)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_418.init = 16'hc088;
    LUT4 i1_4_lut_adj_419 (.A(addr[10]), .B(addr[8]), .C(addr[12]), .D(addr[17]), 
         .Z(n24198)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_419.init = 16'h8000;
    LUT4 mux_1933_i11_4_lut (.A(n27202), .B(n27140), .C(n4073), .D(n28563), 
         .Z(n3163[10])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1933_i11_4_lut.init = 16'hc0ca;
    LUT4 pc_1__bdd_3_lut_24428 (.A(\pc[1] ), .B(\pc[9] ), .C(counter_hi[3]), 
         .Z(n26202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_1__bdd_3_lut_24428.init = 16'hcaca;
    LUT4 i1_3_lut_adj_420 (.A(n35), .B(n26_adj_2659), .C(n23820), .Z(n23824)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_420.init = 16'h8080;
    LUT4 i1_4_lut_adj_421 (.A(addr[11]), .B(addr[23]), .C(addr[13]), .D(addr[16]), 
         .Z(n24202)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_421.init = 16'h8000;
    LUT4 mux_1073_i15_3_lut (.A(n31[14]), .B(n33[14]), .C(n2035), .Z(n1715[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1077_i15_3_lut (.A(n1[14]), .B(n5[14]), .C(n2055), .Z(n1735[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i15_3_lut.init = 16'hcaca;
    LUT4 mtimecmp_6__I_0_3_lut_4_lut (.A(addr[2]), .B(n27241), .C(data_out_slice[2]), 
         .D(mtimecmp[6]), .Z(mtimecmp_2__N_1939)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(449[27:65])
    defparam mtimecmp_6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 mtimecmp_4__I_0_3_lut_4_lut (.A(addr[2]), .B(n27241), .C(data_out_slice[0]), 
         .D(mtimecmp[4]), .Z(mtimecmp_0__N_1943)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(449[27:65])
    defparam mtimecmp_4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_422 (.A(addr[19]), .B(addr[21]), .C(addr[26]), .D(addr[25]), 
         .Z(n24200)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_422.init = 16'h8000;
    LUT4 i1_4_lut_adj_423 (.A(addr[18]), .B(addr[14]), .C(addr[22]), .D(addr[9]), 
         .Z(n24182)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_423.init = 16'h8000;
    LUT4 i1_2_lut_adj_424 (.A(addr[20]), .B(addr[15]), .Z(n24174)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_424.init = 16'h8888;
    LUT4 n26203_bdd_3_lut (.A(n26203), .B(n26200), .C(n28571), .Z(debug_branch_N_442[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26203_bdd_3_lut.init = 16'hcaca;
    LUT4 i16_4_lut_adj_425 (.A(n4079), .B(clk_c_enable_34), .C(rst_reg_n), 
         .D(n22778), .Z(clk_c_enable_245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i16_4_lut_adj_425.init = 16'hcfca;
    LUT4 i1_4_lut_adj_426 (.A(n27112), .B(n27109), .C(n27106), .D(n23870), 
         .Z(n22778)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_426.init = 16'h1000;
    LUT4 i1_4_lut_adj_427 (.A(n26), .B(n23868), .C(n35), .D(n22_adj_2640), 
         .Z(n23870)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_427.init = 16'hccc8;
    LUT4 mux_2813_i12_3_lut (.A(n27205), .B(n27201), .C(n28563), .Z(n4625[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2813_i12_3_lut.init = 16'hcaca;
    LUT4 mux_2813_i13_3_lut (.A(n27205), .B(n27199), .C(n28563), .Z(n4625[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2813_i13_3_lut.init = 16'hcaca;
    LUT4 mux_346_i2_3_lut_4_lut (.A(instr_addr_23__N_318[1]), .B(n27255), 
         .C(debug_ret), .D(return_addr[2]), .Z(n1764[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam mux_346_i2_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_2813_i14_3_lut (.A(n27205), .B(n27200), .C(n28563), .Z(n4625[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2813_i14_3_lut.init = 16'hcaca;
    LUT4 mux_2813_i15_3_lut (.A(n27205), .B(n27198), .C(n28563), .Z(n4625[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2813_i15_3_lut.init = 16'hcaca;
    PFUMX i23880 (.BLUT(n26317), .ALUT(n26316), .C0(\imm[1] ), .Z(n26318));
    LUT4 mux_1073_i2_rep_123_3_lut (.A(n31[1]), .B(n33[1]), .C(n2035), 
         .Z(n24666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i2_rep_123_3_lut.init = 16'hcaca;
    LUT4 mux_1984_i7_3_lut (.A(n3397[6]), .B(n3350[6]), .C(n4079), .Z(n3438[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1984_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1984_i6_3_lut (.A(n3397[5]), .B(n3350[5]), .C(n4079), .Z(n3438[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1984_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1077_i2_3_lut (.A(n1[1]), .B(n5[1]), .C(n2055), .Z(n1735[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i2_3_lut.init = 16'hcaca;
    LUT4 mux_1984_i4_3_lut (.A(n3397[3]), .B(n3350[3]), .C(n4079), .Z(n3438[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1984_i4_3_lut.init = 16'hcaca;
    LUT4 i17750_3_lut_4_lut (.A(n27109), .B(n27106), .C(n23682), .D(addr_offset[2]), 
         .Z(n21[0])) /* synthesis lut_function=(!(A (D)+!A !(B (C (D))+!B (D)))) */ ;
    defparam i17750_3_lut_4_lut.init = 16'h51aa;
    PFUMX i24742 (.BLUT(n28142), .ALUT(n28141), .C0(n25707), .Z(n28143));
    LUT4 mux_1073_i3_rep_125_3_lut (.A(n31[2]), .B(n33[2]), .C(n2035), 
         .Z(n24668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1073_i3_rep_125_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_3_lut_4_lut_adj_428 (.A(n22_adj_2640), .B(n27092), .C(n27207), 
         .D(rst_reg_n), .Z(n22637)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam i1_3_lut_3_lut_4_lut_adj_428.init = 16'h7000;
    LUT4 mux_1077_i3_3_lut (.A(n1[2]), .B(n5[2]), .C(n2055), .Z(n1735[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1077_i3_3_lut.init = 16'hcaca;
    LUT4 i23501_2_lut_4_lut (.A(n27109), .B(n27106), .C(n23682), .D(rst_reg_n), 
         .Z(clk_c_enable_229)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B (D)))) */ ;
    defparam i23501_2_lut_4_lut.init = 16'h04ff;
    PFUMX i22836 (.BLUT(n25175), .ALUT(n25176), .C0(counter_hi[3]), .Z(n25179));
    LUT4 mux_1984_i2_3_lut (.A(n3397[1]), .B(n26436), .C(n4079), .Z(n3438[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1984_i2_3_lut.init = 16'hcaca;
    LUT4 i43_3_lut_4_lut (.A(n27159), .B(n27178), .C(n27209), .D(n23), 
         .Z(n26_adj_2659)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam i43_3_lut_4_lut.init = 16'h2f20;
    PFUMX i22837 (.BLUT(n25177), .ALUT(n25178), .C0(counter_hi[3]), .Z(n25180));
    LUT4 n4061_bdd_3_lut_23909_4_lut (.A(n22_adj_2640), .B(n27092), .C(rst_reg_n), 
         .D(n27204), .Z(n26347)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam n4061_bdd_3_lut_23909_4_lut.init = 16'h7000;
    PFUMX i22843 (.BLUT(n25182), .ALUT(n25183), .C0(counter_hi[3]), .Z(n25186));
    LUT4 i12489_2_lut_3_lut_4_lut (.A(n22_adj_2640), .B(n27092), .C(n27205), 
         .D(n22704), .Z(n3087[5])) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i12489_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i1_3_lut_adj_429 (.A(n8274), .B(n28563), .C(n28575), .Z(n23450)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_429.init = 16'h4040;
    PFUMX i22844 (.BLUT(n25184), .ALUT(n25185), .C0(counter_hi[3]), .Z(n25187));
    LUT4 i1_4_lut_adj_430 (.A(n27205), .B(n28575), .C(n27204), .D(n27211), 
         .Z(n23804)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_430.init = 16'hc088;
    LUT4 i1_4_lut_adj_431 (.A(n27197), .B(rst_reg_n), .C(n27203), .D(n27211), 
         .Z(n23744)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_431.init = 16'hc088;
    LUT4 i1_4_lut_adj_432 (.A(addr_out[3]), .B(n27238), .C(addr_offset[3]), 
         .D(addr_offset[2]), .Z(n23045)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(266[43:70])
    defparam i1_4_lut_adj_432.init = 16'h965a;
    PFUMX i29 (.BLUT(n11), .ALUT(n13), .C0(n28563), .Z(n16_adj_2645));
    LUT4 i1_4_lut_adj_433 (.A(n27108), .B(n22369), .C(n8), .D(n23678), 
         .Z(n22226)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B))) */ ;
    defparam i1_4_lut_adj_433.init = 16'h3b33;
    PFUMX i22850 (.BLUT(n25189), .ALUT(n25190), .C0(counter_hi[3]), .Z(n25193));
    PFUMX i29_adj_434 (.BLUT(n9), .ALUT(n12), .C0(debug_instr_valid), 
          .Z(n16_adj_2660));
    PFUMX i23870 (.BLUT(n26298), .ALUT(n26296), .C0(n4075), .Z(n26299));
    LUT4 mux_1933_i15_3_lut_4_lut (.A(n27205), .B(n27168), .C(n4073), 
         .D(n2874[9]), .Z(n3163[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1933_i15_3_lut_4_lut.init = 16'h8f80;
    PFUMX i22851 (.BLUT(n25191), .ALUT(n25192), .C0(counter_hi[3]), .Z(n25194));
    LUT4 mux_1933_i9_3_lut_4_lut (.A(n27205), .B(n27168), .C(n4073), .D(n4625[7]), 
         .Z(n3163[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1933_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_1933_i10_3_lut_4_lut (.A(n27205), .B(n27168), .C(n4073), 
         .D(n4625[8]), .Z(n3163[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1933_i10_3_lut_4_lut.init = 16'h8f80;
    LUT4 mem_data_ready_bdd_3_lut_24175 (.A(counter_hi[2]), .B(instr_data[9]), 
         .C(instr_data[13]), .Z(n26818)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mem_data_ready_bdd_3_lut_24175.init = 16'he4e4;
    LUT4 is_store_I_0_469_2_lut_rep_619 (.A(is_store), .B(address_ready), 
         .Z(n27244)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(275[22:47])
    defparam is_store_I_0_469_2_lut_rep_619.init = 16'h8888;
    LUT4 i23666_2_lut (.A(n28571), .B(counter_hi[3]), .Z(n25066)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i23666_2_lut.init = 16'heeee;
    LUT4 mem_data_ready_bdd_3_lut_24387 (.A(\qspi_data_buf[25] ), .B(\qspi_data_buf[29] ), 
         .C(counter_hi[2]), .Z(n26819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mem_data_ready_bdd_3_lut_24387.init = 16'hcaca;
    PFUMX i22857 (.BLUT(n25196), .ALUT(n25197), .C0(counter_hi[3]), .Z(n25200));
    LUT4 mux_1933_i17_3_lut_4_lut (.A(n27205), .B(n27168), .C(n4073), 
         .D(n2874[16]), .Z(n3163[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1933_i17_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_3_lut_4_lut_adj_435 (.A(is_store), .B(address_ready), 
         .C(mem_op[1]), .D(rst_reg_n), .Z(data_write_n_1__N_369[1])) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(275[22:47])
    defparam i1_2_lut_3_lut_4_lut_adj_435.init = 16'hf7ff;
    LUT4 i1_2_lut_3_lut_4_lut_adj_436 (.A(is_store), .B(address_ready), 
         .C(mem_op[0]), .D(rst_reg_n), .Z(data_write_n_1__N_369[0])) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(275[22:47])
    defparam i1_2_lut_3_lut_4_lut_adj_436.init = 16'hf7ff;
    PFUMX i22858 (.BLUT(n25198), .ALUT(n25199), .C0(counter_hi[3]), .Z(n25201));
    LUT4 i1_3_lut_adj_437 (.A(n27211), .B(n27200), .C(n28575), .Z(n23712)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_437.init = 16'h4040;
    LUT4 i1_4_lut_adj_438 (.A(no_write_in_progress), .B(data_ready_core), 
         .C(debug_instr_valid), .D(is_load), .Z(debug_rd_3__N_1575)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_4_lut_adj_438.init = 16'h8000;
    LUT4 mem_data_from_read_17__bdd_3_lut_24391 (.A(\mem_data_from_read[17] ), 
         .B(counter_hi[2]), .C(\mem_data_from_read[21] ), .Z(n26821)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam mem_data_from_read_17__bdd_3_lut_24391.init = 16'he2e2;
    LUT4 n26821_bdd_3_lut (.A(n26821), .B(n26820), .C(counter_hi[3]), 
         .Z(n26822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26821_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_2813_i16_3_lut (.A(n27205), .B(n27197), .C(n28563), .Z(n4625[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2813_i16_3_lut.init = 16'hcaca;
    LUT4 i12855_2_lut_3_lut_4_lut (.A(n23682), .B(n27106), .C(n28575), 
         .D(n27109), .Z(clk_c_enable_372)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i12855_2_lut_3_lut_4_lut.init = 16'hf040;
    LUT4 i1_4_lut_adj_439 (.A(n27164), .B(n27184), .C(n27163), .D(n27209), 
         .Z(n4_adj_2638)) /* synthesis lut_function=(!((B (C (D))+!B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_439.init = 16'h0a88;
    LUT4 i1_2_lut_rep_571_3_lut_4_lut (.A(alu_op[0]), .B(n27275), .C(data_rs1[3]), 
         .D(n27276), .Z(n27196)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_rep_571_3_lut_4_lut.init = 16'hf040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_440 (.A(alu_op[0]), .B(n27275), .C(data_rs1[2]), 
         .D(n27276), .Z(n18144)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_3_lut_4_lut_adj_440.init = 16'hf040;
    PFUMX i23865 (.BLUT(n26293), .ALUT(n26290), .C0(n4075), .Z(n26294));
    LUT4 i13_3_lut_4_lut (.A(alu_op[0]), .B(n27275), .C(data_rs1[2]), 
         .D(n27276), .Z(n8_adj_2666)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i22324_3_lut_4_lut (.A(alu_op[0]), .B(n27275), .C(data_rs1[0]), 
         .D(n27276), .Z(n24605)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i22324_3_lut_4_lut.init = 16'hff80;
    LUT4 i25_3_lut_4_lut (.A(alu_op[0]), .B(n27275), .C(data_rs1[1]), 
         .D(n27276), .Z(n20_adj_2672)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i25_3_lut_4_lut.init = 16'h8f80;
    LUT4 i20_3_lut_4_lut (.A(alu_op[0]), .B(n27275), .C(data_rs1[3]), 
         .D(n27276), .Z(n14)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i20_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_1083_i2_3_lut (.A(n24666), .B(n1735[1]), .C(n27260), .Z(instr[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1083_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_441 (.A(clk_c_enable_282), .B(n27179), .C(n27185), 
         .D(n27162), .Z(n2328)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_441.init = 16'ha888;
    LUT4 mux_346_i1_3_lut_4_lut (.A(n27277), .B(\instr_addr_23__N_318[0] ), 
         .C(debug_ret), .D(return_addr[1]), .Z(n1764[0])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam mux_346_i1_3_lut_4_lut.init = 16'hf606;
    LUT4 i1_3_lut_4_lut_adj_442 (.A(n27277), .B(\instr_addr_23__N_318[0] ), 
         .C(\instr_write_offset[3] ), .D(instr_addr_23__N_318[1]), .Z(n23398)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i1_3_lut_4_lut_adj_442.init = 16'h78f0;
    LUT4 mie_10__bdd_4_lut (.A(mie[10]), .B(counter_hi[3]), .C(mie[2]), 
         .D(counter_hi[4]), .Z(n26854)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B+!(C (D)))) */ ;
    defparam mie_10__bdd_4_lut.init = 16'hb8aa;
    LUT4 i4140_2_lut_rep_608_3_lut (.A(n27277), .B(\instr_addr_23__N_318[0] ), 
         .C(instr_addr_23__N_318[1]), .Z(n27233)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i4140_2_lut_rep_608_3_lut.init = 16'h7878;
    LUT4 i1_4_lut_adj_443 (.A(clk_c_enable_282), .B(n27179), .C(n20), 
         .D(n25), .Z(n2330)) /* synthesis lut_function=(A (B+!(C+(D)))) */ ;
    defparam i1_4_lut_adj_443.init = 16'h888a;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n27306), .B(alu_b_in[0]), .C(n27267), 
         .D(cy_adj_2646), .Z(n24124)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hc66c;
    LUT4 i1_4_lut_adj_444 (.A(n27205), .B(n28575), .C(n27206), .D(n27211), 
         .Z(n23768)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_444.init = 16'hc088;
    LUT4 mie_10__bdd_4_lut_24199 (.A(mie[6]), .B(mie[14]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n26853)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam mie_10__bdd_4_lut_24199.init = 16'hcac0;
    LUT4 i1_3_lut_4_lut_4_lut_adj_445 (.A(n27306), .B(cmp), .C(alu_b_in[1]), 
         .D(alu_a_in[1]), .Z(n23342)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_3_lut_4_lut_4_lut_adj_445.init = 16'hd00d;
    LUT4 i4155_2_lut_rep_594_4_lut_4_lut (.A(n27306), .B(mtime_out[0]), 
         .C(n27257), .D(cy_adj_2673), .Z(n27219)) /* synthesis lut_function=(A (B (D))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i4155_2_lut_rep_594_4_lut_4_lut.init = 16'hc840;
    PFUMX mux_1083_i14 (.BLUT(n1715[13]), .ALUT(n1735[13]), .C0(n27260), 
          .Z(instr[29]));
    LUT4 cy_I_0_3_lut_rep_611_4_lut_4_lut (.A(n27306), .B(cy_adj_2673), 
         .C(time_pulse_r), .D(n8869), .Z(n27236)) /* synthesis lut_function=(A (B)+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam cy_I_0_3_lut_rep_611_4_lut_4_lut.init = 16'hd8dd;
    LUT4 tmp_data_in_3__I_124_i4_4_lut_4_lut_4_lut (.A(n27306), .B(data_rs1[3]), 
         .C(interrupt_core), .D(n27279), .Z(tmp_data_in_3__N_1514[3])) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam tmp_data_in_3__I_124_i4_4_lut_4_lut_4_lut.init = 16'h505c;
    PFUMX mux_1083_i13 (.BLUT(n1715[12]), .ALUT(n1735[12]), .C0(n27260), 
          .Z(instr[28]));
    LUT4 n25708_bdd_4_lut (.A(n28563), .B(n27212), .C(n27211), .D(n28564), 
         .Z(n26857)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !((C)+!B)) */ ;
    defparam n25708_bdd_4_lut.init = 16'h8c8e;
    LUT4 i1_4_lut_adj_446 (.A(n27212), .B(n27129), .C(n27205), .D(n24583), 
         .Z(n22080)) /* synthesis lut_function=(!((B (C+!(D))+!B (C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_446.init = 16'h0a22;
    LUT4 i12754_4_lut_4_lut (.A(n27306), .B(\imm[1] ), .C(mcause[2]), 
         .D(mstatus_mte), .Z(n8162)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i12754_4_lut_4_lut.init = 16'h5140;
    LUT4 i4052_2_lut_rep_529_3_lut_4_lut_4_lut (.A(n27306), .B(alu_b_in[0]), 
         .C(n27267), .D(cy_adj_2646), .Z(n27154)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i4052_2_lut_rep_529_3_lut_4_lut_4_lut.init = 16'h3810;
    PFUMX mux_1083_i10 (.BLUT(n1715[9]), .ALUT(n1735[9]), .C0(n27260), 
          .Z(instr[25]));
    LUT4 i4104_2_lut_4_lut_4_lut (.A(n27306), .B(instrret_count[0]), .C(instr_retired), 
         .D(cy_adj_2642), .Z(increment_result_3__N_1925[0])) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i4104_2_lut_4_lut_4_lut.init = 16'h369c;
    LUT4 i4106_2_lut_rep_604_4_lut_4_lut (.A(n27306), .B(instrret_count[0]), 
         .C(instr_retired), .D(cy_adj_2642), .Z(n27229)) /* synthesis lut_function=(A (B (D))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i4106_2_lut_rep_604_4_lut_4_lut.init = 16'hc840;
    LUT4 i4084_2_lut_3_lut_4_lut_4_lut (.A(n27306), .B(cycle_count_wide[0]), 
         .C(cycle_count_wide[1]), .D(cy), .Z(increment_result_3__N_1911[1])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i4084_2_lut_3_lut_4_lut_4_lut.init = 16'h3cb4;
    PFUMX mux_1083_i9 (.BLUT(n1715[8]), .ALUT(n1735[8]), .C0(n27260), 
          .Z(instr[24]));
    LUT4 i1_3_lut_4_lut_adj_447 (.A(n27306), .B(rst_reg_n), .C(data_ready_latch), 
         .D(address_ready), .Z(clk_c_enable_14)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_447.init = 16'hff7f;
    LUT4 i1_3_lut_4_lut_adj_448 (.A(n27306), .B(rst_reg_n), .C(data_ready_latch), 
         .D(n27126), .Z(n23201)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_448.init = 16'h0008;
    PFUMX mux_1083_i4 (.BLUT(n1715[3]), .ALUT(n1735[3]), .C0(n27260), 
          .Z(instr[19]));
    LUT4 mux_2835_i2_4_lut_4_lut (.A(n27309), .B(n27306), .C(mstatus_mpie), 
         .D(mstatus_mie), .Z(csr_read_3__N_1439[3])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam mux_2835_i2_4_lut_4_lut.init = 16'h7340;
    LUT4 n3244_bdd_3_lut_23864_4_lut (.A(instr[31]), .B(n27179), .C(n27101), 
         .D(n26280), .Z(n26281)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3244_bdd_3_lut_23864_4_lut.init = 16'hf808;
    LUT4 i3314_2_lut_3_lut_4_lut (.A(n23682), .B(n27106), .C(rst_reg_n), 
         .D(n27109), .Z(clk_c_enable_26)) /* synthesis lut_function=(!(A (C)+!A (B (C (D))+!B (C)))) */ ;
    defparam i3314_2_lut_3_lut_4_lut.init = 16'h0f4f;
    PFUMX mux_1083_i12_rep_127 (.BLUT(n1715[11]), .ALUT(n1735[11]), .C0(n27260), 
          .Z(instr[27]));
    FD1S3IX counter_hi_3236__i3_rep_764 (.D(n34[1]), .CK(clk_c), .CD(n27326), 
            .Q(n28573));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3236__i3_rep_764.GSR = "DISABLED";
    LUT4 mux_2857_i5_4_lut_4_lut (.A(instr[31]), .B(n27179), .C(n27131), 
         .D(n4075), .Z(n4745[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2857_i5_4_lut_4_lut.init = 16'ha088;
    LUT4 n1_bdd_4_lut (.A(n28563), .B(n27212), .C(n27148), .D(n28564), 
         .Z(n26868)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;
    defparam n1_bdd_4_lut.init = 16'hc800;
    LUT4 mux_1938_i16_3_lut_4_lut (.A(instr[31]), .B(n27179), .C(n27101), 
         .D(n4745[8]), .Z(n3232[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1938_i16_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_1938_i15_3_lut_4_lut (.A(instr[31]), .B(n27179), .C(n27101), 
         .D(n4745[7]), .Z(n3232[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1938_i15_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_1938_i14_3_lut_4_lut (.A(instr[31]), .B(n27179), .C(n27101), 
         .D(n4745[6]), .Z(n3232[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1938_i14_3_lut_4_lut.init = 16'hf808;
    LUT4 n14584_bdd_3_lut_24271 (.A(n1715[14]), .B(n1735[14]), .C(n27260), 
         .Z(instr[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n14584_bdd_3_lut_24271.init = 16'hcaca;
    LUT4 i23667_3_lut_4_lut (.A(n27298), .B(counter_hi[3]), .C(is_timer_addr), 
         .D(data_out_3__N_1385), .Z(n25057)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam i23667_3_lut_4_lut.init = 16'hff04;
    LUT4 mux_1938_i13_3_lut_4_lut (.A(instr[31]), .B(n27179), .C(n27101), 
         .D(n4745[5]), .Z(n3232[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1938_i13_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_2857_i10_3_lut_4_lut (.A(instr[31]), .B(n27179), .C(n27101), 
         .D(n24658), .Z(n4745[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2857_i10_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_3_lut_adj_449 (.A(n27112), .B(n8274), .C(n28575), .Z(n23908)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_adj_449.init = 16'h1010;
    PFUMX i23856 (.BLUT(n26281), .ALUT(n26278), .C0(n4075), .Z(n26282));
    LUT4 n3244_bdd_3_lut_23869_4_lut (.A(instr[31]), .B(n27179), .C(n27101), 
         .D(n26292), .Z(n26293)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3244_bdd_3_lut_23869_4_lut.init = 16'hf808;
    LUT4 n3244_bdd_3_lut_23873_4_lut (.A(instr[31]), .B(n27179), .C(n27101), 
         .D(n26297), .Z(n26298)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3244_bdd_3_lut_23873_4_lut.init = 16'hf808;
    LUT4 mux_1984_i32_3_lut_4_lut (.A(instr[31]), .B(n27179), .C(n4079), 
         .D(n3397[17]), .Z(n3350[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1984_i32_3_lut_4_lut.init = 16'h8f80;
    PFUMX i24351 (.BLUT(n27402), .ALUT(n27403), .C0(n27260), .Z(instr[31]));
    PFUMX i24349 (.BLUT(n27399), .ALUT(n27400), .C0(counter_hi[2]), .Z(n27401));
    PFUMX i24347 (.BLUT(n27395), .ALUT(n27396), .C0(counter_hi[2]), .Z(n27397));
    FD1S3IX counter_hi_3236__i4_rep_762 (.D(n34[2]), .CK(clk_c), .CD(n27326), 
            .Q(n28571));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3236__i4_rep_762.GSR = "DISABLED";
    PFUMX i24343 (.BLUT(n27389), .ALUT(n27390), .C0(n27260), .Z(n27391));
    tinyQV_time i_timer (.clk_c(clk_c), .n27326(n27326), .mtimecmp_2__N_1939(mtimecmp_2__N_1939), 
            .mtimecmp_1__N_1941(mtimecmp_1__N_1941), .mtimecmp_0__N_1943(mtimecmp_0__N_1943), 
            .time_pulse_r(time_pulse_r), .clk_c_enable_71(clk_c_enable_71), 
            .n27257(n27257), .\mtimecmp[7] (mtimecmp[7]), .\mtimecmp[6] (mtimecmp[6]), 
            .\mtimecmp[5] (mtimecmp[5]), .\mtimecmp[4] (mtimecmp[4]), .clk_c_enable_276(clk_c_enable_276), 
            .\addr[2] (addr[2]), .timer_data({timer_data}), .\mtime_out[0] (mtime_out[0]), 
            .mtimecmp_3__N_1935(mtimecmp_3__N_1935), .timer_interrupt(timer_interrupt), 
            .n8869(n8869), .cy(cy_adj_2673), .rst_reg_n(rst_reg_n), .n28575(n28575), 
            .\cycle_count_wide[3] (cycle_count_wide[3]), .n27180(n27180), 
            .clk_c_enable_73(clk_c_enable_73), .no_write_in_progress(no_write_in_progress), 
            .is_store(is_store), .n27300(n27300), .\reg_access[4][3] (\reg_access[4] [3]), 
            .clk_c_enable_31(clk_c_enable_31), .address_ready(address_ready), 
            .n27226(n27226), .\instr_data[0] (instr_data[0]), .\instr_data_0__15__N_638[0] (instr_data_0__15__N_638[0]), 
            .clk_c_enable_272(clk_c_enable_272), .\reg_access[3][2] (\reg_access[3] [2]), 
            .clk_c_enable_60(clk_c_enable_60), .n27309(n27309), .clk_c_enable_64(clk_c_enable_64), 
            .n27306(n27306), .clk_c_enable_67(clk_c_enable_67), .clk_c_enable_231(clk_c_enable_231), 
            .\instr_data[1] (instr_data[1]), .\instr_data_0__15__N_638[49] (instr_data_0__15__N_638[49]), 
            .n27358(n27358), .is_timer_addr(is_timer_addr), .n27219(n27219), 
            .n27236(n27236), .\data_out_slice[2] (data_out_slice[2]), .n27220(n27220), 
            .n27222(n27222), .\data_out_slice[0] (data_out_slice[0]), .n27214(n27214)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(450[17] 461[6])
    tinyqv_decoder i_decoder (.n27197(n27197), .\instr[31] (instr[31]), 
            .n27205(n27205), .n4722(n4703[12]), .n28564(n28564), .n26779(n26779), 
            .n27212(n27212), .n26206(n26206), .n27209(n27209), .n27179(n27179), 
            .n28563(n28563), .n27211(n27211), .n26745(n26745), .n23744(n23744), 
            .n8274(n8274), .n26(n26_adj_2659), .n23750(n23750), .n27189(n27189), 
            .n27185(n27185), .n23842(n23842), .n23792(n23792), .n23798(n23798), 
            .n7(n7), .n27172(n27172), .n27200(n27200), .is_auipc_de(is_auipc_de), 
            .n28575(n28575), .n23820(n23820), .n2328(n2328), .\instr[17] (instr[17]), 
            .n4634(n4625[7]), .n2163(n2161[2]), .n23804(n23804), .n23810(n23810), 
            .n27186(n27186), .n26803(n26803), .\mem_op_de[2] (mem_op_de[2]), 
            .n6(n6), .n27174(n27174), .\instr[26] (instr[26]), .n27173(n27173), 
            .n27192(n27192), .n27203(n27203), .n27178(n27178), .n27177(n27177), 
            .n27204(n27204), .n27202(n27202), .n9124(n9124), .n27158(n27158), 
            .n26804(n26804), .n27152(n27152), .n27199(n27199), .n27201(n27201), 
            .n27166(n27166), .n27198(n27198), .is_alu_imm_de(is_alu_imm_de), 
            .n27142(n27142), .n23588(n23588), .n19(n19), .n23594(n23594), 
            .n2898(n2874[8]), .n27131(n27131), .n27130(n27130), .n27157(n27157), 
            .n27206(n27206), .n27207(n27207), .n27132(n27132), .n27138(n27138), 
            .n28562(n28562), .n27(n27_adj_2665), .n24030(n24030), .\instr[25] (instr[25]), 
            .n3259(n3232[5]), .n27101(n27101), .n4057(n4057), .n27099(n27099), 
            .n27260(n27260), .n4075(n4075), .n24988(n24988), .\instr[27] (instr[27]), 
            .n3257(n3232[7]), .n24516(n24516), .n28143(n28143), .n27_adj_7(n27), 
            .n27135(n27135), .n23650(n23650), .\instr[30] (instr[30]), 
            .n3(n3), .n27145(n27145), .n23658(n23658), .n27184(n27184), 
            .n1741(n1735[10]), .n24640(n24640), .n23868(n23868), .\instr[16] (instr[16]), 
            .n2141(n2138[1]), .n4707(n4703[27]), .n27151(n27151), .\instr[20] (instr[20]), 
            .n22909(n22909), .mem_op_increment_reg_de(mem_op_increment_reg_de), 
            .\alu_op_3__N_1337[2] (alu_op_3__N_1337[2]), .n10(n10_adj_2671), 
            .n24(n24_adj_2656), .n23712(n23712), .n23718(n23718), .n23756(n23756), 
            .n23762(n23762), .n27148(n27148), .n14587(n14587), .n27121(n27121), 
            .n27175(n27175), .is_ret_de(is_ret_de), .n27176(n27176), .clk_c_enable_34(clk_c_enable_34), 
            .\additional_mem_ops[2] (additional_mem_ops[2]), .n4117(n4116[2]), 
            .n30(n30), .n30_adj_8(n30_adj_2662), .n7711(n7711), .n27156(n27156), 
            .n6985(n6985), .n26867(n26867), .is_system_de(is_system_de), 
            .n2897(n2874[9]), .n22100(n22100), .n22101(n22101), .n15(n15_adj_2658), 
            .n23768(n23768), .n23774(n23774), .n27128(n27128), .alu_op_de({alu_op_de}), 
            .n25707(n25707), .n26874(n26874), .n4718(n4703[16]), .\instr[24] (instr[24]), 
            .n4710(n4703[24]), .\instr[29] (instr[29]), .n4705(n4703[29]), 
            .n4709(n4703[25]), .n26289(n26289), .n26290(n26290), .n4719(n4703[15]), 
            .n24641(n24641), .n1745(n1735[6]), .n24635(n24635), .n15_adj_9(n15_adj_2663), 
            .n25708(n25708), .n4720(n4703[14]), .\instr[19] (instr[19]), 
            .n26296(n26296), .n27123(n27123), .n26277(n26277), .n26278(n26278), 
            .\instr[28] (instr[28]), .n4706(n4703[28]), .is_alu_reg_de(is_alu_reg_de), 
            .n1744(n1735[7]), .n24633(n24633), .n1746(n1735[5]), .n24627(n24627), 
            .n8123(n8123), .n1747(n1735[4]), .n24625(n24625), .is_jalr_de(is_jalr_de), 
            .is_lui_N_1365(is_lui_N_1365), .is_lui_de(is_lui_de), .n4721(n4703[13]), 
            .is_store_de(is_store_de), .n8(n8_adj_2657), .n25126(n25126), 
            .is_load_de(is_load_de), .n23544(n23544), .n27167(n27167), 
            .is_branch_de(is_branch_de), .n22164(n22164), .n15_adj_10(n15_adj_2641), 
            .n30_adj_11(n30_adj_2661), .n23598(n23598), .n27109(n27109), 
            .n3166(n3163[29]), .is_jal_de(is_jal_de), .n27170(n27170), 
            .n12(n12_adj_2674), .n4729(n4703[5]), .n4727(n4703[7]), .n4734(n4703[0]), 
            .n4730(n4703[4]), .\mem_op_de[1] (mem_op_de[1]), .n2890(n2874[16]), 
            .n23682(n23682), .n27114(n27114), .n27108(n27108), .n10_adj_12(n10_c), 
            .n27169(n27169), .n23698(n23698), .n23704(n23704), .n27129(n27129)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    tinyqv_core i_core (.n26927(n26927), .\imm[0] (imm[0]), .mstatus_mpie(mstatus_mpie), 
            .clk_c(clk_c), .clk_c_enable_424(clk_c_enable_424), .n9675(n9675), 
            .n27218(n27218), .time_hi({time_hi}), .n27326(n27326), .\debug_branch_N_446[31] (debug_branch_N_446[31]), 
            .tmp_data({Open_5, Open_6, tmp_data[29:28], Open_7, Open_8, 
            Open_9, Open_10, Open_11, Open_12, Open_13, Open_14, 
            Open_15, Open_16, Open_17, Open_18, Open_19, Open_20, 
            Open_21, Open_22, Open_23, Open_24, Open_25, Open_26, 
            Open_27, Open_28, Open_29, Open_30, Open_31, Open_32, 
            Open_33, Open_34}), .load_done(load_done), .clk_c_enable_71(clk_c_enable_71), 
            .n6982(n6982), .instr_retired(instr_retired), .n14783(n14783), 
            .instr_complete_N_1647(instr_complete_N_1647), .n27367(n27367), 
            .n27369(n27369), .n24404(n24404), .n27287(n27287), .n27348(n27348), 
            .n15(n15_adj_2637), .cycle({cycle}), .\shift_amt[0] (shift_amt[0]), 
            .n92({n92}), .n5434(n5434), .n27279(n27279), .clk_c_enable_73(clk_c_enable_73), 
            .\mie[14] (mie[14]), .n926(n926), .\mie[13] (mie[13]), .\mie[10] (mie[10]), 
            .n893(n893), .\mie[9] (mie[9]), .\mie[6] (mie[6]), .n860(n860), 
            .\mie[5] (mie[5]), .\mie[2] (mie[2]), .n793(n793), .\mie[1] (mie[1]), 
            .cmp(cmp), .\mepc[0] (mepc[0]), .\next_fsm_state_3__N_2499[3] (\next_fsm_state_3__N_2499[3] ), 
            .cy(cy_adj_2646), .mstatus_mte(mstatus_mte), .n26930(n26930), 
            .\imm[10] (\imm[10] ), .n27374(n27374), .n27305(n27305), .n27238(n27238), 
            .\addr_out[0] (addr_out[0]), .\addr_out[1] (\addr_out[1] ), 
            .\next_pc_for_core[7] (\next_pc_for_core[7] ), .\next_pc_for_core[3] (\next_pc_for_core[3] ), 
            .counter_hi({counter_hi}), .\addr_out[23] (addr_out[23]), .\addr_out[22] (addr_out[22]), 
            .\addr_out[21] (addr_out[21]), .\tmp_data[31] (tmp_data[31]), 
            .alu_op({alu_op}), .\tmp_data[30] (tmp_data[30]), .\addr_out[20] (addr_out[20]), 
            .\addr_out[19] (addr_out[19]), .\addr_out[18] (addr_out[18]), 
            .\addr_out[17] (addr_out[17]), .\next_pc_for_core[15] (\next_pc_for_core[15] ), 
            .\next_pc_for_core[11] (\next_pc_for_core[11] ), .\addr_out[16] (addr_out[16]), 
            .n27309(n27309), .\imm[6] (\imm[6] ), .\imm[2] (\imm[2] ), 
            .\addr_out[15] (addr_out[15]), .\next_pc_for_core[23] (\next_pc_for_core[23] ), 
            .\next_pc_for_core[19] (\next_pc_for_core[19] ), .\addr_out[14] (addr_out[14]), 
            .\addr_out[13] (addr_out[13]), .\addr_out[12] (addr_out[12]), 
            .\addr_out[11] (addr_out[11]), .\addr_out[10] (addr_out[10]), 
            .\addr_out[9] (addr_out[9]), .\addr_out[8] (addr_out[8]), .\addr_out[7] (addr_out[7]), 
            .n27196(n27196), .mstatus_mie(mstatus_mie), .\addr_out[6] (addr_out[6]), 
            .\addr_out[5] (addr_out[5]), .\addr_out[4] (addr_out[4]), .\addr_out[3] (addr_out[3]), 
            .n22121(n22121), .\imm[1] (\imm[1] ), .n27332(n27332), .interrupt_core(interrupt_core), 
            .n27306(n27306), .\csr_read_3__N_1443[0] (csr_read_3__N_1443[0]), 
            .\csr_read_3__N_1451[0] (csr_read_3__N_1451[0]), .n27292(n27292), 
            .\cycle_count_wide[0] (cycle_count_wide[0]), .\instrret_count[0] (instrret_count[0]), 
            .\debug_rd_3__N_405[28] (debug_rd_3__N_405[28]), .\debug_rd_3__N_405[30] (debug_rd_3__N_405[30]), 
            .\debug_rd_3__N_405[29] (debug_rd_3__N_405[29]), .\debug_rd_3__N_405[31] (debug_rd_3__N_405[31]), 
            .\next_pc_for_core[14] (\next_pc_for_core[14] ), .\next_pc_for_core[10] (\next_pc_for_core[10] ), 
            .\time_count[2] (time_count[2]), .mip_reg({mip_reg}), .clk_c_enable_350(clk_c_enable_350), 
            .n24216(n24216), .n8162(n8162), .\next_pc_for_core[22] (\next_pc_for_core[22] ), 
            .\next_pc_for_core[18] (\next_pc_for_core[18] ), .clk_c_enable_367(clk_c_enable_367), 
            .n26855(n26855), .n27112(n27112), .n27106(n27106), .n23738(n23738), 
            .n27109(n27109), .n2123(n2120[1]), .n23798(n23798), .n22721(n22721), 
            .n23750(n23750), .n22745(n22745), .n23718(n23718), .n22551(n22551), 
            .n24822(n24822), .\debug_branch_N_442[28] (debug_branch_N_442[28]), 
            .n157(n157), .n23704(n23704), .n22559(n22559), .n23774(n23774), 
            .n22733(n22733), .n23450(n23450), .n22700(n22700), .n8(n8_adj_2668), 
            .n23820(n23820), .n26(n26_adj_2659), .n26345(n26345), .n23690(n23690), 
            .n2322(n2322), .n23810(n23810), .n22715(n22715), .debug_rd_3__N_1575(debug_rd_3__N_1575), 
            .load_top_bit_next_N_1731(load_top_bit_next_N_1731), .mem_op({mem_op}), 
            .n24516(n24516), .n8274(n8274), .n24(n24_adj_2670), .n23838(n23838), 
            .n23824(n23824), .n3295(n3273[10]), .n23762(n23762), .n22739(n22739), 
            .\imm[4] (\imm[4] ), .n27329(n27329), .n24360(n24360), .n23842(n23842), 
            .n12(n12_adj_2674), .n23848(n23848), .n24601(n24601), .n24505(n24505), 
            .\a_for_shift_right[31] (a_for_shift_right[31]), .data_rs1({data_rs1}), 
            .n23894(n23894), .n22784(n22784), .n23650(n23650), .n27122(n27122), 
            .n23656(n23656), .n27391(n27391), .n23498(n23498), .n23594(n23594), 
            .n27114(n27114), .n27108(n27108), .n23598(n23598), .n27110(n27110), 
            .rst_reg_n(rst_reg_n), .n27342(n27342), .load_top_bit(load_top_bit), 
            .data_out_3__N_1385(data_out_3__N_1385), .alu_a_in_3__N_1552(alu_a_in_3__N_1552), 
            .\debug_branch_N_442[29] (debug_branch_N_442[29]), .\alu_a_in[1] (alu_a_in[1]), 
            .\debug_branch_N_840[29] (\debug_branch_N_840[29] ), .\timer_data[1] (timer_data[1]), 
            .is_timer_addr(is_timer_addr), .n27347(n27347), .\mul_out[2] (\mul_out[2] ), 
            .\mul_out[3] (\mul_out[3] ), .\mul_out[1] (\mul_out[1] ), .n27290(n27290), 
            .\ui_in_sync[1] (\ui_in_sync[1] ), .n1167(n1167), .n27276(n27276), 
            .n27249(n27249), .n27248(n27248), .n26686(n26686), .n27302(n27302), 
            .n25069(n25069), .n26049(n26049), .clk_c_enable_276(clk_c_enable_276), 
            .debug_rd({debug_rd}), .\shift_amt[1] (shift_amt[1]), .stall_core(stall_core), 
            .n27263(n27263), .is_load(is_load), .n856(n856), .n22226(n22226), 
            .clk_c_enable_423(clk_c_enable_423), .n22898(n22898), .any_additional_mem_ops(any_additional_mem_ops), 
            .clk_c_enable_275(clk_c_enable_275), .accum({accum}), .d_3__N_1868({d_3__N_1868}), 
            .\shift_out[1] (shift_out[1]), .n27368(n27368), .n27366(n27366), 
            .\imm[7] (\imm[7] ), .n7717(n7717), .n26733(n26733), .\debug_branch_N_450[0] (debug_branch_N_450[0]), 
            .debug_instr_valid(debug_instr_valid), .n27376(n27376), .n27256(n27256), 
            .data_rs2({data_rs2}), .alu_b_in({alu_b_in}), .is_auipc(is_auipc), 
            .is_jal(is_jal), .n5160(n5160), .n5171(n5167[0]), .n22499(n22499), 
            .n4575({n4575[1], n4577}), .n1766(n1764[1]), .\instr_write_offset_3__N_934[1] (instr_write_offset_3__N_934[1]), 
            .n1767(n1764[0]), .\instr_write_offset_3__N_934[0] (instr_write_offset_3__N_934[0]), 
            .n27111(n27111), .n27288(n27288), .n1768({n1768}), .pc_2__N_932({pc_2__N_932}), 
            .\mcause[1] (mcause[1]), .n616(n611[1]), .\mcause[2] (mcause[2]), 
            .\mcause[5] (mcause[5]), .is_branch(is_branch), .is_jalr(is_jalr), 
            .is_system(is_system), .is_alu_imm(is_alu_imm), .is_alu_reg(is_alu_reg), 
            .clk_c_enable_422(clk_c_enable_422), .n15206(n15206), .\debug_branch_N_450[3] (debug_branch_N_450[3]), 
            .is_lui(is_lui), .n27350(n27350), .\debug_branch_N_442[31] (debug_branch_N_442[31]), 
            .n27293(n27293), .n27322(n27322), .interrupt_pending_N_1671(interrupt_pending_N_1671), 
            .no_write_in_progress(no_write_in_progress), .n5168(n5167[3]), 
            .\imm[3] (\imm[3] ), .\imm[5] (\imm[5] ), .n22178(n22178), 
            .n26802(n26802), .\imm[8] (\imm[8] ), .\imm[9] (\imm[9] ), 
            .\debug_branch_N_442[30] (debug_branch_N_442[30]), .n26318(n26318), 
            .n27338(n27338), .n28573(n28573), .n28571(n28571), .n18(n34[2]), 
            .n27343(n27343), .timer_interrupt(timer_interrupt), .n27349(n27349), 
            .n27362(n27362), .n25142(n25142), .n27231(n27231), .n20(n20_adj_2672), 
            .n14(n14), .n24838(n24838), .debug_rd_3__N_413(debug_rd_3__N_413), 
            .\tmp_data_in_3__N_1514[3] (tmp_data_in_3__N_1514[3]), .n27274(n27274), 
            .\debug_rd_3__N_1567[0] (debug_rd_3__N_1567[0]), .debug_reg_wen_N_1692(debug_reg_wen_N_1692), 
            .\shift_out[0] (shift_out[0]), .n25132(n25132), .\pc[21] (\pc[21] ), 
            .\pc[17] (\pc[17] ), .n26200(n26200), .\next_pc_for_core[20] (\next_pc_for_core[20] ), 
            .\next_pc_for_core[16] (\next_pc_for_core[16] ), .n225(n225_adj_2669), 
            .\pc[23] (\pc[23] ), .\pc[19] (\pc[19] ), .n26175(n26175), 
            .\pc[20] (\pc[20] ), .\pc[16] (\pc[16] ), .n225_adj_4(n225), 
            .\next_pc_for_core[21] (\next_pc_for_core[21] ), .\next_pc_for_core[17] (\next_pc_for_core[17] ), 
            .n226(n226), .\pc[22] (\pc[22] ), .\pc[18] (\pc[18] ), .n26195(n26195), 
            .n26685(n26685), .\data_out_slice[2] (data_out_slice[2]), .n27214(n27214), 
            .n27223(n27223), .\mtimecmp[7] (mtimecmp[7]), .mtimecmp_3__N_1935(mtimecmp_3__N_1935), 
            .n24772(n24772), .\debug_branch_N_446[29] (debug_branch_N_446[29]), 
            .n27222(n27222), .\mtimecmp[5] (mtimecmp[5]), .mtimecmp_1__N_1941(mtimecmp_1__N_1941), 
            .n27247(n27247), .n27296(n27296), .n27321(n27321), .address_ready(address_ready), 
            .n28575(n28575), .n24775(n24775), .\debug_branch_N_446[30] (debug_branch_N_446[30]), 
            .n26336(n26336), .n26335(n26335), .\addr_offset[2] (addr_offset[2]), 
            .n701(n699[0]), .is_store(is_store), .n24611(n24611), .n26717(n26717), 
            .\debug_branch_N_450[2] (debug_branch_N_450[2]), .n24774(n24774), 
            .\csr_read_3__N_1459[0] (csr_read_3__N_1459[0]), .n24616(n24616), 
            .\debug_branch_N_840[31] (debug_branch_N_840[31]), .\data_out_slice[0] (data_out_slice[0]), 
            .\csr_read_3__N_1459[3] (csr_read_3__N_1459[3]), .n27023(n27023), 
            .\csr_read_3__N_1459[1] (csr_read_3__N_1459[1]), .\cycle_count_wide[1] (cycle_count_wide[1]), 
            .\csr_read_3__N_1439[3] (csr_read_3__N_1439[3]), .n22090(n22090), 
            .\imm[11] (\imm[11] ), .n26976(n26976), .instr_complete_N_1651(instr_complete_N_1651), 
            .\time_count[3] (time_count[3]), .n5115(n5114[3]), .n26932(n26932), 
            .\next_accum[5] (\next_accum[5] ), .\next_accum[6] (\next_accum[6] ), 
            .\next_accum[7] (\next_accum[7] ), .GND_net(GND_net), .VCC_net(VCC_net), 
            .\next_accum[8] (\next_accum[8] ), .\next_accum[9] (\next_accum[9] ), 
            .\next_accum[10] (\next_accum[10] ), .\next_accum[11] (\next_accum[11] ), 
            .\next_accum[12] (\next_accum[12] ), .\next_accum[13] (\next_accum[13] ), 
            .\next_accum[14] (\next_accum[14] ), .\next_accum[15] (\next_accum[15] ), 
            .\next_accum[16] (\next_accum[16] ), .\next_accum[17] (\next_accum[17] ), 
            .\next_accum[18] (\next_accum[18] ), .\next_accum[19] (\next_accum[19] ), 
            .\next_accum[4] (\next_accum[4] ), .n62(n62), .n27377(n27377), 
            .n8157(n8157), .n8153(n8153), .n7278(n7278), .n25292(n25292), 
            .n63(n63), .\shift_amt[5] (shift_amt[5]), .rs1({rs1}), .rd({rd}), 
            .rs2({rs2}), .return_addr({return_addr}), .\reg_access[4][3] (\reg_access[4] [3]), 
            .n24605(n24605), .\reg_access[3][2] (\reg_access[3] [2]), .n27205(n27205), 
            .n27113(n27113), .n2356(n2352[0]), .cy_adj_5(cy_adj_2642), 
            .\increment_result_3__N_1925[0] (increment_result_3__N_1925[0]), 
            .\instrret_count[3] (instrret_count[3]), .n27229(n27229), .n27246(n27246), 
            .cy_adj_6(cy), .\increment_result_3__N_1911[1] (increment_result_3__N_1911[1]), 
            .\increment_result_3__N_1911[0] (increment_result_3__N_1911[0]), 
            .\cycle_count_wide[6] (cycle_count_wide[6]), .\cycle_count_wide[5] (cycle_count_wide[5]), 
            .\cycle_count_wide[4] (cycle_count_wide[4]), .\cycle_count_wide[3] (cycle_count_wide[3]), 
            .n27228(n27228), .n27245(n27245), .n27180(n27180), .n27187(n27187), 
            .n24124(n24124), .n27188(n27188), .n27252(n27252), .n27215(n27215), 
            .n27154(n27154), .n27181(n27181), .n23342(n23342), .n27267(n27267), 
            .n27266(n27266), .n27270(n27270)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(322[72] 368[6])
    
endmodule
//
// Verilog Description of module tinyQV_time
//

module tinyQV_time (clk_c, n27326, mtimecmp_2__N_1939, mtimecmp_1__N_1941, 
            mtimecmp_0__N_1943, time_pulse_r, clk_c_enable_71, n27257, 
            \mtimecmp[7] , \mtimecmp[6] , \mtimecmp[5] , \mtimecmp[4] , 
            clk_c_enable_276, \addr[2] , timer_data, \mtime_out[0] , 
            mtimecmp_3__N_1935, timer_interrupt, n8869, cy, rst_reg_n, 
            n28575, \cycle_count_wide[3] , n27180, clk_c_enable_73, 
            no_write_in_progress, is_store, n27300, \reg_access[4][3] , 
            clk_c_enable_31, address_ready, n27226, \instr_data[0] , 
            \instr_data_0__15__N_638[0] , clk_c_enable_272, \reg_access[3][2] , 
            clk_c_enable_60, n27309, clk_c_enable_64, n27306, clk_c_enable_67, 
            clk_c_enable_231, \instr_data[1] , \instr_data_0__15__N_638[49] , 
            n27358, is_timer_addr, n27219, n27236, \data_out_slice[2] , 
            n27220, n27222, \data_out_slice[0] , n27214) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output n27326;
    input mtimecmp_2__N_1939;
    input mtimecmp_1__N_1941;
    input mtimecmp_0__N_1943;
    output time_pulse_r;
    input clk_c_enable_71;
    output n27257;
    output \mtimecmp[7] ;
    output \mtimecmp[6] ;
    output \mtimecmp[5] ;
    output \mtimecmp[4] ;
    input clk_c_enable_276;
    input \addr[2] ;
    output [3:0]timer_data;
    output \mtime_out[0] ;
    input mtimecmp_3__N_1935;
    output timer_interrupt;
    input n8869;
    output cy;
    input rst_reg_n;
    input n28575;
    input \cycle_count_wide[3] ;
    input n27180;
    output clk_c_enable_73;
    input no_write_in_progress;
    input is_store;
    output n27300;
    input \reg_access[4][3] ;
    output clk_c_enable_31;
    input address_ready;
    output n27226;
    input \instr_data[0] ;
    output \instr_data_0__15__N_638[0] ;
    output clk_c_enable_272;
    input \reg_access[3][2] ;
    output clk_c_enable_60;
    input n27309;
    output clk_c_enable_64;
    input n27306;
    output clk_c_enable_67;
    output clk_c_enable_231;
    input \instr_data[1] ;
    output \instr_data_0__15__N_638[49] ;
    input n27358;
    input is_timer_addr;
    input n27219;
    input n27236;
    input \data_out_slice[2] ;
    input n27220;
    input n27222;
    input \data_out_slice[0] ;
    input n27214;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [31:0]mtimecmp;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(30[16:24])
    
    wire cy_c;
    wire [4:0]comparison;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[16:26])
    wire [3:0]mtime_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(29[16:25])
    
    wire timer_interrupt_N_1954, n27380, n27381, n6, n4, n2;
    
    FD1S3IX mtimecmp_2__90 (.D(mtimecmp_2__N_1939), .CK(clk_c), .CD(n27326), 
            .Q(mtimecmp[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_2__90.GSR = "DISABLED";
    FD1S3IX mtimecmp_1__91 (.D(mtimecmp_1__N_1941), .CK(clk_c), .CD(n27326), 
            .Q(mtimecmp[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_1__91.GSR = "DISABLED";
    FD1S3IX mtimecmp_0__92 (.D(mtimecmp_0__N_1943), .CK(clk_c), .CD(n27326), 
            .Q(mtimecmp[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_0__92.GSR = "DISABLED";
    FD1S3IX time_pulse_r_95 (.D(n27257), .CK(clk_c), .CD(clk_c_enable_71), 
            .Q(time_pulse_r)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(82[12] 85[8])
    defparam time_pulse_r_95.GSR = "DISABLED";
    FD1S3AX mtimecmp_30__62 (.D(mtimecmp[2]), .CK(clk_c), .Q(mtimecmp[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_30__62.GSR = "DISABLED";
    FD1S3AX mtimecmp_29__63 (.D(mtimecmp[1]), .CK(clk_c), .Q(mtimecmp[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_29__63.GSR = "DISABLED";
    FD1S3AX mtimecmp_28__64 (.D(mtimecmp[0]), .CK(clk_c), .Q(mtimecmp[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_28__64.GSR = "DISABLED";
    FD1S3AX mtimecmp_27__65 (.D(mtimecmp[31]), .CK(clk_c), .Q(mtimecmp[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_27__65.GSR = "DISABLED";
    FD1S3AX mtimecmp_26__66 (.D(mtimecmp[30]), .CK(clk_c), .Q(mtimecmp[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_26__66.GSR = "DISABLED";
    FD1S3AX mtimecmp_25__67 (.D(mtimecmp[29]), .CK(clk_c), .Q(mtimecmp[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_25__67.GSR = "DISABLED";
    FD1S3AX mtimecmp_24__68 (.D(mtimecmp[28]), .CK(clk_c), .Q(mtimecmp[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_24__68.GSR = "DISABLED";
    FD1S3AX mtimecmp_23__69 (.D(mtimecmp[27]), .CK(clk_c), .Q(mtimecmp[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_23__69.GSR = "DISABLED";
    FD1S3AX mtimecmp_22__70 (.D(mtimecmp[26]), .CK(clk_c), .Q(mtimecmp[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_22__70.GSR = "DISABLED";
    FD1S3AX mtimecmp_21__71 (.D(mtimecmp[25]), .CK(clk_c), .Q(mtimecmp[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_21__71.GSR = "DISABLED";
    FD1S3AX mtimecmp_20__72 (.D(mtimecmp[24]), .CK(clk_c), .Q(mtimecmp[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_20__72.GSR = "DISABLED";
    FD1S3AX mtimecmp_19__73 (.D(mtimecmp[23]), .CK(clk_c), .Q(mtimecmp[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_19__73.GSR = "DISABLED";
    FD1S3AX mtimecmp_18__74 (.D(mtimecmp[22]), .CK(clk_c), .Q(mtimecmp[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_18__74.GSR = "DISABLED";
    FD1S3AX mtimecmp_17__75 (.D(mtimecmp[21]), .CK(clk_c), .Q(mtimecmp[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_17__75.GSR = "DISABLED";
    FD1S3AX mtimecmp_16__76 (.D(mtimecmp[20]), .CK(clk_c), .Q(mtimecmp[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_16__76.GSR = "DISABLED";
    FD1S3AX mtimecmp_15__77 (.D(mtimecmp[19]), .CK(clk_c), .Q(mtimecmp[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_15__77.GSR = "DISABLED";
    FD1S3AX mtimecmp_14__78 (.D(mtimecmp[18]), .CK(clk_c), .Q(mtimecmp[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_14__78.GSR = "DISABLED";
    FD1S3AX mtimecmp_13__79 (.D(mtimecmp[17]), .CK(clk_c), .Q(mtimecmp[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_13__79.GSR = "DISABLED";
    FD1S3AX mtimecmp_12__80 (.D(mtimecmp[16]), .CK(clk_c), .Q(mtimecmp[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_12__80.GSR = "DISABLED";
    FD1S3AX mtimecmp_11__81 (.D(mtimecmp[15]), .CK(clk_c), .Q(mtimecmp[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_11__81.GSR = "DISABLED";
    FD1S3AX mtimecmp_10__82 (.D(mtimecmp[14]), .CK(clk_c), .Q(mtimecmp[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_10__82.GSR = "DISABLED";
    FD1S3AX mtimecmp_9__83 (.D(mtimecmp[13]), .CK(clk_c), .Q(mtimecmp[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_9__83.GSR = "DISABLED";
    FD1S3AX mtimecmp_8__84 (.D(mtimecmp[12]), .CK(clk_c), .Q(mtimecmp[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_8__84.GSR = "DISABLED";
    FD1S3AX mtimecmp_7__85 (.D(mtimecmp[11]), .CK(clk_c), .Q(\mtimecmp[7] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_7__85.GSR = "DISABLED";
    FD1S3AX mtimecmp_6__86 (.D(mtimecmp[10]), .CK(clk_c), .Q(\mtimecmp[6] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_6__86.GSR = "DISABLED";
    FD1S3AX mtimecmp_5__87 (.D(mtimecmp[9]), .CK(clk_c), .Q(\mtimecmp[5] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_5__87.GSR = "DISABLED";
    FD1S3AX mtimecmp_4__88 (.D(mtimecmp[8]), .CK(clk_c), .Q(\mtimecmp[4] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_4__88.GSR = "DISABLED";
    FD1S3JX cy_93 (.D(comparison[4]), .CK(clk_c), .PD(clk_c_enable_276), 
            .Q(cy_c)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(74[12] 76[8])
    defparam cy_93.GSR = "DISABLED";
    FD1S3AX mtimecmp_31__61 (.D(mtimecmp[3]), .CK(clk_c), .Q(mtimecmp[31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_31__61.GSR = "DISABLED";
    LUT4 mtime_out_3__I_0_96_i4_3_lut (.A(mtime_out[3]), .B(\mtimecmp[7] ), 
         .C(\addr[2] ), .Z(timer_data[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i4_3_lut.init = 16'hcaca;
    LUT4 mtime_out_3__I_0_96_i3_3_lut (.A(mtime_out[2]), .B(\mtimecmp[6] ), 
         .C(\addr[2] ), .Z(timer_data[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i3_3_lut.init = 16'hcaca;
    LUT4 mtime_out_3__I_0_96_i1_3_lut (.A(\mtime_out[0] ), .B(\mtimecmp[4] ), 
         .C(\addr[2] ), .Z(timer_data[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i1_3_lut.init = 16'hcaca;
    FD1S3IX mtimecmp_3__89 (.D(mtimecmp_3__N_1935), .CK(clk_c), .CD(n27326), 
            .Q(mtimecmp[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_3__89.GSR = "DISABLED";
    FD1P3AX timer_interrupt_94 (.D(timer_interrupt_N_1954), .SP(clk_c_enable_276), 
            .CK(clk_c), .Q(timer_interrupt)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(78[12] 80[8])
    defparam timer_interrupt_94.GSR = "DISABLED";
    LUT4 mtime_out_3__I_0_96_i2_3_lut (.A(mtime_out[1]), .B(\mtimecmp[5] ), 
         .C(\addr[2] ), .Z(timer_data[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i2_3_lut.init = 16'hcaca;
    PFUMX i24337 (.BLUT(n27380), .ALUT(n27381), .C0(mtime_out[2]), .Z(timer_interrupt_N_1954));
    LUT4 i3974_3_lut (.A(mtime_out[3]), .B(\mtimecmp[7] ), .C(n6), .Z(comparison[4])) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i3974_3_lut.init = 16'hb2b2;
    LUT4 i3967_3_lut (.A(mtime_out[2]), .B(\mtimecmp[6] ), .C(n4), .Z(n6)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i3967_3_lut.init = 16'hb2b2;
    LUT4 i3960_3_lut (.A(mtime_out[1]), .B(\mtimecmp[5] ), .C(n2), .Z(n4)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i3960_3_lut.init = 16'hb2b2;
    LUT4 i3953_3_lut (.A(\mtime_out[0] ), .B(\mtimecmp[4] ), .C(cy_c), 
         .Z(n2)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i3953_3_lut.init = 16'hb2b2;
    LUT4 i12346_4_lut_then_4_lut (.A(mtime_out[3]), .B(n4), .C(\mtimecmp[6] ), 
         .D(\mtimecmp[7] ), .Z(n27381)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;
    defparam i12346_4_lut_then_4_lut.init = 16'h8241;
    LUT4 i12346_4_lut_else_4_lut (.A(mtime_out[3]), .B(n4), .C(\mtimecmp[6] ), 
         .D(\mtimecmp[7] ), .Z(n27380)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A (B (C+(D))+!B !(C (D))))) */ ;
    defparam i12346_4_lut_else_4_lut.init = 16'h1824;
    LUT4 time_pulse_I_0_2_lut_rep_632 (.A(n8869), .B(time_pulse_r), .Z(n27257)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(37[14:39])
    defparam time_pulse_I_0_2_lut_rep_632.init = 16'hdddd;
    tinyqv_counter i_mtime (.clk_c(clk_c), .n27326(n27326), .cy(cy), .mtime_out({mtime_out[3:1], 
            \mtime_out[0] }), .rst_reg_n(rst_reg_n), .n28575(n28575), 
            .\cycle_count_wide[3] (\cycle_count_wide[3] ), .n27180(n27180), 
            .clk_c_enable_276(clk_c_enable_276), .clk_c_enable_73(clk_c_enable_73), 
            .no_write_in_progress(no_write_in_progress), .is_store(is_store), 
            .n27300(n27300), .\reg_access[4][3] (\reg_access[4][3] ), .clk_c_enable_31(clk_c_enable_31), 
            .address_ready(address_ready), .n27226(n27226), .\instr_data[0] (\instr_data[0] ), 
            .\instr_data_0__15__N_638[0] (\instr_data_0__15__N_638[0] ), .clk_c_enable_272(clk_c_enable_272), 
            .\reg_access[3][2] (\reg_access[3][2] ), .clk_c_enable_60(clk_c_enable_60), 
            .n27309(n27309), .clk_c_enable_64(clk_c_enable_64), .n27306(n27306), 
            .clk_c_enable_67(clk_c_enable_67), .clk_c_enable_231(clk_c_enable_231), 
            .\instr_data[1] (\instr_data[1] ), .\instr_data_0__15__N_638[49] (\instr_data_0__15__N_638[49] ), 
            .\addr[2] (\addr[2] ), .n27358(n27358), .is_timer_addr(is_timer_addr), 
            .n27219(n27219), .n27236(n27236), .\data_out_slice[2] (\data_out_slice[2] ), 
            .n27220(n27220), .n27222(n27222), .\data_out_slice[0] (\data_out_slice[0] ), 
            .n27214(n27214)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(34[20] 42[6])
    
endmodule
//
// Verilog Description of module tinyqv_counter
//

module tinyqv_counter (clk_c, n27326, cy, mtime_out, rst_reg_n, n28575, 
            \cycle_count_wide[3] , n27180, clk_c_enable_276, clk_c_enable_73, 
            no_write_in_progress, is_store, n27300, \reg_access[4][3] , 
            clk_c_enable_31, address_ready, n27226, \instr_data[0] , 
            \instr_data_0__15__N_638[0] , clk_c_enable_272, \reg_access[3][2] , 
            clk_c_enable_60, n27309, clk_c_enable_64, n27306, clk_c_enable_67, 
            clk_c_enable_231, \instr_data[1] , \instr_data_0__15__N_638[49] , 
            \addr[2] , n27358, is_timer_addr, n27219, n27236, \data_out_slice[2] , 
            n27220, n27222, \data_out_slice[0] , n27214) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output n27326;
    output cy;
    output [3:0]mtime_out;
    input rst_reg_n;
    input n28575;
    input \cycle_count_wide[3] ;
    input n27180;
    input clk_c_enable_276;
    output clk_c_enable_73;
    input no_write_in_progress;
    input is_store;
    output n27300;
    input \reg_access[4][3] ;
    output clk_c_enable_31;
    input address_ready;
    output n27226;
    input \instr_data[0] ;
    output \instr_data_0__15__N_638[0] ;
    output clk_c_enable_272;
    input \reg_access[3][2] ;
    output clk_c_enable_60;
    input n27309;
    output clk_c_enable_64;
    input n27306;
    output clk_c_enable_67;
    output clk_c_enable_231;
    input \instr_data[1] ;
    output \instr_data_0__15__N_638[49] ;
    input \addr[2] ;
    input n27358;
    input is_timer_addr;
    input n27219;
    input n27236;
    input \data_out_slice[2] ;
    input n27220;
    input n27222;
    input \data_out_slice[0] ;
    input n27214;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    wire [4:0]increment_result;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[16:32])
    
    wire n8128;
    wire [4:0]increment_result_3__N_1925;
    
    wire n27193, n27161;
    
    FD1S3IX register_2__48 (.D(increment_result[2]), .CK(clk_c), .CD(n27326), 
            .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result[1]), .CK(clk_c), .CD(n27326), 
            .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(increment_result[0]), .CK(clk_c), .CD(n27326), 
            .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3IX cy_51 (.D(increment_result_3__N_1925[4]), .CK(clk_c), .CD(n8128), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(register[10])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(register[9])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(register[8])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(mtime_out[3])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(register[10]), .CK(clk_c), .Q(mtime_out[2])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(register[9]), .CK(clk_c), .Q(mtime_out[1])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(register[8]), .CK(clk_c), .Q(mtime_out[0])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result[3]), .CK(clk_c), .CD(n27326), 
            .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 rstn_I_0_1_lut_rep_701 (.A(rst_reg_n), .Z(n27326)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam rstn_I_0_1_lut_rep_701.init = 16'h5555;
    LUT4 i3350_4_lut_4_lut (.A(n28575), .B(\cycle_count_wide[3] ), .C(n27180), 
         .D(clk_c_enable_276), .Z(clk_c_enable_73)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3350_4_lut_4_lut.init = 16'hd555;
    LUT4 i3324_3_lut_rep_675_3_lut (.A(n28575), .B(no_write_in_progress), 
         .C(is_store), .Z(n27300)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3324_3_lut_rep_675_3_lut.init = 16'hd5d5;
    LUT4 i23495_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(\reg_access[4][3] ), 
         .C(no_write_in_progress), .D(is_store), .Z(clk_c_enable_31)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i23495_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i1_2_lut_rep_601_3_lut_3_lut (.A(n28575), .B(address_ready), .C(is_store), 
         .Z(n27226)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_rep_601_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i12171_2_lut_2_lut (.A(rst_reg_n), .B(\instr_data[0] ), .Z(\instr_data_0__15__N_638[0] )) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i12171_2_lut_2_lut.init = 16'hdddd;
    LUT4 i3321_2_lut_2_lut (.A(rst_reg_n), .B(address_ready), .Z(clk_c_enable_272)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3321_2_lut_2_lut.init = 16'hdddd;
    LUT4 i23432_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(\reg_access[3][2] ), 
         .C(no_write_in_progress), .D(is_store), .Z(clk_c_enable_60)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i23432_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i23556_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n27309), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_64)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i23556_2_lut_4_lut_4_lut.init = 16'h3111;
    LUT4 i23493_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n27306), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_67)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i23493_2_lut_4_lut_4_lut.init = 16'h3111;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(clk_c_enable_276), 
         .C(address_ready), .D(is_store), .Z(clk_c_enable_231)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hfddd;
    LUT4 i12437_2_lut_2_lut (.A(rst_reg_n), .B(\instr_data[1] ), .Z(\instr_data_0__15__N_638[49] )) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i12437_2_lut_2_lut.init = 16'hdddd;
    LUT4 i5810_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(\addr[2] ), .C(n27358), 
         .D(is_timer_addr), .Z(n8128)) /* synthesis lut_function=(!(A (B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i5810_2_lut_3_lut_4_lut_4_lut.init = 16'h5755;
    LUT4 i4177_2_lut_3_lut_4_lut (.A(mtime_out[1]), .B(n27219), .C(mtime_out[3]), 
         .D(mtime_out[2]), .Z(increment_result_3__N_1925[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4177_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4163_2_lut_rep_568_3_lut (.A(mtime_out[0]), .B(n27236), .C(mtime_out[1]), 
         .Z(n27193)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4163_2_lut_rep_568_3_lut.init = 16'h8080;
    LUT4 i4170_2_lut_rep_536_3_lut_4_lut (.A(mtime_out[0]), .B(n27236), 
         .C(mtime_out[2]), .D(mtime_out[1]), .Z(n27161)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4170_2_lut_rep_536_3_lut_4_lut.init = 16'h8000;
    LUT4 increment_result_3__I_168_i3_4_lut (.A(mtime_out[2]), .B(\data_out_slice[2] ), 
         .C(n27220), .D(n27193), .Z(increment_result[2])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i3_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_168_i2_4_lut (.A(mtime_out[1]), .B(n27222), 
         .C(n27220), .D(n27219), .Z(increment_result[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i2_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_168_i1_4_lut (.A(mtime_out[0]), .B(\data_out_slice[0] ), 
         .C(n27220), .D(n27236), .Z(increment_result[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i1_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_168_i4_4_lut (.A(mtime_out[3]), .B(n27214), 
         .C(n27220), .D(n27161), .Z(increment_result[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i4_4_lut.init = 16'hc5ca;
    
endmodule
//
// Verilog Description of module tinyqv_decoder
//

module tinyqv_decoder (n27197, \instr[31] , n27205, n4722, n28564, 
            n26779, n27212, n26206, n27209, n27179, n28563, n27211, 
            n26745, n23744, n8274, n26, n23750, n27189, n27185, 
            n23842, n23792, n23798, n7, n27172, n27200, is_auipc_de, 
            n28575, n23820, n2328, \instr[17] , n4634, n2163, n23804, 
            n23810, n27186, n26803, \mem_op_de[2] , n6, n27174, 
            \instr[26] , n27173, n27192, n27203, n27178, n27177, 
            n27204, n27202, n9124, n27158, n26804, n27152, n27199, 
            n27201, n27166, n27198, is_alu_imm_de, n27142, n23588, 
            n19, n23594, n2898, n27131, n27130, n27157, n27206, 
            n27207, n27132, n27138, n28562, n27, n24030, \instr[25] , 
            n3259, n27101, n4057, n27099, n27260, n4075, n24988, 
            \instr[27] , n3257, n24516, n28143, n27_adj_7, n27135, 
            n23650, \instr[30] , n3, n27145, n23658, n27184, n1741, 
            n24640, n23868, \instr[16] , n2141, n4707, n27151, \instr[20] , 
            n22909, mem_op_increment_reg_de, \alu_op_3__N_1337[2] , n10, 
            n24, n23712, n23718, n23756, n23762, n27148, n14587, 
            n27121, n27175, is_ret_de, n27176, clk_c_enable_34, \additional_mem_ops[2] , 
            n4117, n30, n30_adj_8, n7711, n27156, n6985, n26867, 
            is_system_de, n2897, n22100, n22101, n15, n23768, n23774, 
            n27128, alu_op_de, n25707, n26874, n4718, \instr[24] , 
            n4710, \instr[29] , n4705, n4709, n26289, n26290, n4719, 
            n24641, n1745, n24635, n15_adj_9, n25708, n4720, \instr[19] , 
            n26296, n27123, n26277, n26278, \instr[28] , n4706, 
            is_alu_reg_de, n1744, n24633, n1746, n24627, n8123, 
            n1747, n24625, is_jalr_de, is_lui_N_1365, is_lui_de, n4721, 
            is_store_de, n8, n25126, is_load_de, n23544, n27167, 
            is_branch_de, n22164, n15_adj_10, n30_adj_11, n23598, 
            n27109, n3166, is_jal_de, n27170, n12, n4729, n4727, 
            n4734, n4730, \mem_op_de[1] , n2890, n23682, n27114, 
            n27108, n10_adj_12, n27169, n23698, n23704, n27129) /* synthesis syn_module_defined=1 */ ;
    input n27197;
    input \instr[31] ;
    input n27205;
    output n4722;
    input n28564;
    input n26779;
    input n27212;
    input n26206;
    input n27209;
    input n27179;
    input n28563;
    input n27211;
    input n26745;
    input n23744;
    input n8274;
    input n26;
    output n23750;
    input n27189;
    input n27185;
    output n23842;
    input n23792;
    output n23798;
    input n7;
    input n27172;
    input n27200;
    output is_auipc_de;
    input n28575;
    output n23820;
    input n2328;
    input \instr[17] ;
    input n4634;
    output n2163;
    input n23804;
    output n23810;
    input n27186;
    output n26803;
    output \mem_op_de[2] ;
    output n6;
    input n27174;
    input \instr[26] ;
    input n27173;
    input n27192;
    input n27203;
    input n27178;
    input n27177;
    input n27204;
    input n27202;
    output n9124;
    output n27158;
    output n26804;
    input n27152;
    input n27199;
    input n27201;
    output n27166;
    input n27198;
    output is_alu_imm_de;
    output n27142;
    input n23588;
    input n19;
    output n23594;
    output n2898;
    output n27131;
    output n27130;
    output n27157;
    input n27206;
    input n27207;
    output n27132;
    output n27138;
    output n28562;
    input n27;
    output n24030;
    input \instr[25] ;
    output n3259;
    input n27101;
    output n4057;
    output n27099;
    input n27260;
    input n4075;
    output n24988;
    input \instr[27] ;
    output n3257;
    output n24516;
    input n28143;
    output n27_adj_7;
    output n27135;
    output n23650;
    input \instr[30] ;
    input n3;
    output n27145;
    output n23658;
    input n27184;
    input n1741;
    output n24640;
    output n23868;
    input \instr[16] ;
    output n2141;
    output n4707;
    output n27151;
    input \instr[20] ;
    output n22909;
    output mem_op_increment_reg_de;
    output \alu_op_3__N_1337[2] ;
    output n10;
    output n24;
    input n23712;
    output n23718;
    input n23756;
    output n23762;
    output n27148;
    output n14587;
    output n27121;
    input n27175;
    output is_ret_de;
    input n27176;
    input clk_c_enable_34;
    input \additional_mem_ops[2] ;
    output n4117;
    input n30;
    input n30_adj_8;
    output n7711;
    input n27156;
    output n6985;
    output n26867;
    output is_system_de;
    output n2897;
    input n22100;
    output n22101;
    output n15;
    input n23768;
    output n23774;
    input n27128;
    output [3:0]alu_op_de;
    input n25707;
    output n26874;
    output n4718;
    input \instr[24] ;
    output n4710;
    input \instr[29] ;
    output n4705;
    output n4709;
    input n26289;
    output n26290;
    output n4719;
    output n24641;
    input n1745;
    output n24635;
    input n15_adj_9;
    input n25708;
    output n4720;
    input \instr[19] ;
    output n26296;
    output n27123;
    input n26277;
    output n26278;
    input \instr[28] ;
    output n4706;
    output is_alu_reg_de;
    input n1744;
    output n24633;
    input n1746;
    output n24627;
    output n8123;
    input n1747;
    output n24625;
    output is_jalr_de;
    input is_lui_N_1365;
    output is_lui_de;
    output n4721;
    output is_store_de;
    input n8;
    input n25126;
    output is_load_de;
    output n23544;
    input n27167;
    output is_branch_de;
    input n22164;
    input n15_adj_10;
    input n30_adj_11;
    input n23598;
    input n27109;
    output n3166;
    output is_jal_de;
    input n27170;
    output n12;
    output n4729;
    output n4727;
    output n4734;
    output n4730;
    output \mem_op_de[1] ;
    output n2890;
    input n23682;
    input n27114;
    input n27108;
    output n10_adj_12;
    input n27169;
    input n23698;
    output n23704;
    output n27129;
    
    
    wire n26877, n26876, n7601, n27143, n26782, n26781, n26783, 
        n26778, n26780, n26207, n26208, n28567, n28566, n26744, 
        n27137, n26746, n27149, n151, n7_adj_2624, n19_c, n27133, 
        n15222;
    wire [3:0]alu_op_3__N_1170;
    
    wire n23030, alu_op_3__N_1181, n28568, n27834, n27139, alu_op_3__N_1180, 
        is_jal_N_1374, n26785, n3_c, n23046, n27141, imm_31__N_1169, 
        n27144;
    wire [3:0]n155;
    
    wire n24128, n27146, n22000, n22946, mem_op_2__N_1384, n27182, 
        n27829;
    wire [3:0]n328;
    
    wire n27153, n15_c, n15_adj_2628, n15_adj_2629, n14503, n23962, 
        n23956, n24579, n23944;
    wire [2:0]additional_mem_ops_2__N_1129;
    
    wire n7709, n7705, n6983, is_jalr_N_1370, n22965, n15143, n24050;
    
    PFUMX i24217 (.BLUT(n26877), .ALUT(n26876), .C0(n27197), .Z(n7601));
    LUT4 mux_2842_i13_3_lut_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n27205), .Z(n4722)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_2842_i13_3_lut_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i24154 (.BLUT(n26782), .ALUT(n26781), .C0(n28564), .Z(n26783));
    PFUMX i24151 (.BLUT(n26779), .ALUT(n26778), .C0(n27212), .Z(n26780));
    PFUMX i23817 (.BLUT(n26207), .ALUT(n26206), .C0(n27209), .Z(n26208));
    LUT4 i24561_then_4_lut (.A(n27179), .B(n27209), .C(n28563), .D(n27211), 
         .Z(n28567)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam i24561_then_4_lut.init = 16'h4470;
    LUT4 i24561_else_4_lut (.A(n27179), .B(n27209), .C(n28563), .D(n27211), 
         .Z(n28566)) /* synthesis lut_function=(!(A (B+(D))+!A !(B (C+(D))+!B !(D)))) */ ;
    defparam i24561_else_4_lut.init = 16'h4473;
    PFUMX i24132 (.BLUT(n26745), .ALUT(n26744), .C0(n27137), .Z(n26746));
    LUT4 i1_4_lut_4_lut (.A(n27179), .B(n23744), .C(n8274), .D(n26), 
         .Z(n23750)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h0400;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n27179), .B(n27189), .C(n27185), .D(n27212), 
         .Z(n23842)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h1000;
    LUT4 i1_4_lut_4_lut_adj_292 (.A(n27179), .B(n23792), .C(n8274), .D(n26), 
         .Z(n23798)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_292.init = 16'h0400;
    LUT4 i23461_3_lut_4_lut_4_lut (.A(n27179), .B(n7), .C(n27172), .D(n27200), 
         .Z(is_auipc_de)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i23461_3_lut_4_lut_4_lut.init = 16'h0200;
    LUT4 i1_4_lut_4_lut_adj_293 (.A(n27179), .B(n28575), .C(n27205), .D(n8274), 
         .Z(n23820)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_293.init = 16'h0040;
    LUT4 mux_1383_i3_4_lut_4_lut (.A(n27179), .B(n2328), .C(\instr[17] ), 
         .D(n4634), .Z(n2163)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;
    defparam mux_1383_i3_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i1_4_lut_4_lut_adj_294 (.A(n27179), .B(n23804), .C(n8274), .D(n26), 
         .Z(n23810)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_294.init = 16'h0400;
    LUT4 is_alu_imm_N_1367_bdd_3_lut_24162_4_lut (.A(n27205), .B(n27186), 
         .C(n27211), .D(n28563), .Z(n26803)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam is_alu_imm_N_1367_bdd_3_lut_24162_4_lut.init = 16'h0002;
    LUT4 i1_3_lut_4_lut (.A(n27185), .B(n27189), .C(n26746), .D(n27149), 
         .Z(\mem_op_de[2] )) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0010;
    LUT4 i23665_2_lut_3_lut_3_lut_4_lut (.A(n27185), .B(n27189), .C(n27211), 
         .D(n27179), .Z(n6)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;
    defparam i23665_2_lut_3_lut_3_lut_4_lut.init = 16'h1101;
    LUT4 i5281_2_lut_3_lut_4_lut (.A(n27200), .B(n27174), .C(\instr[26] ), 
         .D(n27173), .Z(n151)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam i5281_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 instr_1__I_0_139_i7_4_lut (.A(n27192), .B(n27203), .C(n27212), 
         .D(n27178), .Z(n7_adj_2624)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam instr_1__I_0_139_i7_4_lut.init = 16'h0a3a;
    LUT4 i6784_3_lut_4_lut (.A(n27177), .B(n27204), .C(n27202), .D(n28563), 
         .Z(n9124)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(282[33:52])
    defparam i6784_3_lut_4_lut.init = 16'h10f0;
    LUT4 is_alu_imm_N_1367_bdd_3_lut_4_lut (.A(n27202), .B(n27158), .C(n27211), 
         .D(n28563), .Z(n26804)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(282[33:52])
    defparam is_alu_imm_N_1367_bdd_3_lut_4_lut.init = 16'h2000;
    LUT4 i12907_4_lut (.A(n19_c), .B(n27133), .C(n28564), .D(n27152), 
         .Z(n15222)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i12907_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut (.A(n7601), .B(alu_op_3__N_1170[2]), .C(n28564), .Z(n23030)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 instr_6__I_0_142_i10_2_lut_3_lut (.A(n27199), .B(n27201), .C(n27166), 
         .Z(alu_op_3__N_1181)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam instr_6__I_0_142_i10_2_lut_3_lut.init = 16'h0808;
    LUT4 i1_3_lut_rep_541 (.A(n27197), .B(n27198), .C(n27200), .Z(n27166)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_rep_541.init = 16'hf7f7;
    LUT4 n27833_bdd_3_lut_4_lut (.A(n28563), .B(n27179), .C(n27212), .D(n28568), 
         .Z(n27834)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam n27833_bdd_3_lut_4_lut.init = 16'h2f20;
    LUT4 instr_6__I_0_157_i9_2_lut_rep_514_4_lut (.A(n27197), .B(n27198), 
         .C(n27200), .D(n27174), .Z(n27139)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam instr_6__I_0_157_i9_2_lut_rep_514_4_lut.init = 16'hfff7;
    LUT4 instr_6__I_0_130_i10_2_lut_4_lut (.A(n27197), .B(n27198), .C(n27200), 
         .D(n27172), .Z(alu_op_3__N_1180)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam instr_6__I_0_130_i10_2_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n27209), .B(n28564), .C(n27211), 
         .D(n28563), .Z(is_jal_N_1374)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 n26785_bdd_3_lut_4_lut (.A(n27209), .B(n28564), .C(n26780), .D(n26785), 
         .Z(is_alu_imm_de)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam n26785_bdd_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut (.A(n27149), .B(n3_c), .C(n27204), .D(n27137), .Z(n23046)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i1_4_lut.init = 16'h5044;
    LUT4 i1_3_lut_rep_516_4_lut (.A(n27198), .B(n27197), .C(n27200), .D(n27209), 
         .Z(n27141)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(218[25] 223[32])
    defparam i1_3_lut_rep_516_4_lut.init = 16'h8000;
    LUT4 i1_3_lut_rep_517_4_lut (.A(n27201), .B(n27200), .C(n27199), .D(n7), 
         .Z(n27142)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam i1_3_lut_rep_517_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_518_3_lut (.A(n27199), .B(n27201), .C(n27200), .Z(n27143)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam i1_2_lut_rep_518_3_lut.init = 16'hbfbf;
    LUT4 i1_4_lut_4_lut_adj_295 (.A(n27179), .B(n23588), .C(n8274), .D(n19), 
         .Z(n23594)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_295.init = 16'h0400;
    LUT4 mux_1900_i9_3_lut_4_lut_4_lut_4_lut (.A(n27199), .B(n27201), .C(n27212), 
         .D(n27200), .Z(n2898)) /* synthesis lut_function=(A (C+(D))+!A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_1900_i9_3_lut_4_lut_4_lut_4_lut.init = 16'hefa0;
    LUT4 instr_6__I_0_127_i10_2_lut_3_lut_4_lut (.A(n27199), .B(n27201), 
         .C(n27173), .D(n27200), .Z(imm_31__N_1169)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam instr_6__I_0_127_i10_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i4686_4_lut (.A(n27205), .B(n27211), .C(n151), .D(n27139), 
         .Z(alu_op_3__N_1170[0])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[18] 85[91])
    defparam i4686_4_lut.init = 16'hcacc;
    LUT4 i12282_2_lut_rep_506_3_lut_4_lut (.A(n27199), .B(n27201), .C(n27197), 
         .D(n27200), .Z(n27131)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam i12282_2_lut_rep_506_3_lut_4_lut.init = 16'hfbff;
    LUT4 i23554_2_lut_rep_508_3_lut_4_lut (.A(n27198), .B(n27197), .C(n27174), 
         .D(n27200), .Z(n27133)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(66[27:51])
    defparam i23554_2_lut_rep_508_3_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_519_3_lut (.A(n27198), .B(n27197), .C(n27200), .Z(n27144)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(66[27:51])
    defparam i1_2_lut_rep_519_3_lut.init = 16'hfdfd;
    LUT4 mux_29_i2_4_lut (.A(n28563), .B(n151), .C(n27139), .D(n27211), 
         .Z(alu_op_3__N_1170[1])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[18] 85[91])
    defparam mux_29_i2_4_lut.init = 16'hfaca;
    LUT4 i1_2_lut_rep_505_3_lut_4_lut (.A(n27198), .B(n27197), .C(n27174), 
         .D(n27200), .Z(n27130)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(66[27:51])
    defparam i1_2_lut_rep_505_3_lut_4_lut.init = 16'hfffd;
    LUT4 mux_28_i3_3_lut_4_lut_3_lut_4_lut (.A(n27201), .B(n27199), .C(n27166), 
         .D(n28563), .Z(n155[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam mux_28_i3_3_lut_4_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 n22212_bdd_2_lut_24153_3_lut_4_lut (.A(n27201), .B(n27199), .C(n7), 
         .D(n27200), .Z(n26781)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam n22212_bdd_2_lut_24153_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n27201), .B(n27199), .C(n7601), .D(n27166), 
         .Z(n24128)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_rep_532_3_lut_4_lut (.A(n27212), .B(n28564), .C(n27211), 
         .D(n28563), .Z(n27157)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i1_2_lut_rep_532_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_rep_521_4_lut (.A(n27206), .B(n27207), .C(n27203), .D(n27204), 
         .Z(n27146)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(282[33:52])
    defparam i1_3_lut_rep_521_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_533_3_lut (.A(n27206), .B(n27207), .C(n27204), .Z(n27158)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(282[33:52])
    defparam i1_2_lut_rep_533_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_507_3_lut_4_lut (.A(n27206), .B(n27207), .C(n27202), 
         .D(n27204), .Z(n27132)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(282[33:52])
    defparam i1_2_lut_rep_507_3_lut_4_lut.init = 16'hffef;
    LUT4 i23421_2_lut_rep_513_3_lut_4_lut (.A(n28563), .B(n27211), .C(n27212), 
         .D(n28564), .Z(n27138)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i23421_2_lut_rep_513_3_lut_4_lut.init = 16'h0001;
    LUT4 n22212_bdd_2_lut_24156_3_lut (.A(n28563), .B(n27211), .C(n27212), 
         .Z(n26782)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam n22212_bdd_2_lut_24156_3_lut.init = 16'h0101;
    LUT4 i23505_2_lut_3_lut (.A(n28563), .B(n27211), .C(n27212), .Z(n22000)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i23505_2_lut_3_lut.init = 16'h0101;
    LUT4 i169_2_lut_rep_758 (.A(n27209), .B(n28564), .C(n27211), .Z(n28562)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i169_2_lut_rep_758.init = 16'h7070;
    LUT4 is_alu_imm_N_1367_bdd_2_lut_3_lut_4_lut (.A(n28563), .B(n27211), 
         .C(n27186), .D(n27205), .Z(n26778)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam is_alu_imm_N_1367_bdd_2_lut_3_lut_4_lut.init = 16'h1110;
    LUT4 i1_3_lut_4_lut_adj_296 (.A(n27209), .B(n28564), .C(n27), .D(n27212), 
         .Z(n24030)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !((D)+!C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_3_lut_4_lut_adj_296.init = 16'h88f8;
    LUT4 i5497_3_lut_4_lut (.A(n27209), .B(n28564), .C(\instr[25] ), .D(n27205), 
         .Z(n3259)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5497_3_lut_4_lut.init = 16'hf780;
    LUT4 i5494_rep_474_4_lut (.A(n27209), .B(n28564), .C(n27101), .D(n4057), 
         .Z(n27099)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5494_rep_474_4_lut.init = 16'h08f8;
    LUT4 i23697_3_lut_4_lut (.A(n27209), .B(n28564), .C(n27260), .D(n4075), 
         .Z(n24988)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i23697_3_lut_4_lut.init = 16'hff08;
    LUT4 i5501_3_lut_4_lut (.A(n27209), .B(n28564), .C(\instr[27] ), .D(n27202), 
         .Z(n3257)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5501_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_29_i3_4_lut (.A(\instr[27] ), .B(n155[2]), .C(n27139), .D(n151), 
         .Z(alu_op_3__N_1170[2])) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[18] 85[91])
    defparam mux_29_i3_4_lut.init = 16'haccc;
    LUT4 i22239_2_lut_3_lut (.A(n27209), .B(n28564), .C(n28563), .Z(n24516)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i22239_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut (.A(n27209), .B(n28564), .C(n28143), .Z(n27_adj_7)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i168_2_lut_rep_510_2_lut_3_lut (.A(n27209), .B(n28564), .C(n28563), 
         .Z(n27135)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i168_2_lut_rep_510_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_adj_297 (.A(n27209), .B(n28564), .C(n27202), 
         .D(n27146), .Z(n23650)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_2_lut_3_lut_3_lut_4_lut_adj_297.init = 16'h7770;
    LUT4 i12509_4_lut (.A(\instr[30] ), .B(n151), .C(n27198), .D(n3), 
         .Z(n155[3])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(85[18:91])
    defparam i12509_4_lut.init = 16'hecee;
    LUT4 i12699_2_lut_rep_520_3_lut (.A(n27209), .B(n28564), .C(\instr[31] ), 
         .Z(n27145)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i12699_2_lut_rep_520_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_298 (.A(n27209), .B(n28564), .C(n28575), .Z(n23658)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_2_lut_3_lut_adj_298.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_adj_299 (.A(n27209), .B(n28564), .C(n27211), 
         .D(n27184), .Z(n22946)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_2_lut_3_lut_3_lut_4_lut_adj_299.init = 16'h7000;
    LUT4 mux_1083_i11_rep_97_3_lut_3_lut_4_lut (.A(n27209), .B(n28564), 
         .C(n1741), .D(n27206), .Z(n24640)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam mux_1083_i11_rep_97_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_300 (.A(n27209), .B(n28564), .C(n8274), 
         .D(n28575), .Z(n23868)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_2_lut_3_lut_4_lut_adj_300.init = 16'h0700;
    LUT4 i12518_2_lut_3_lut (.A(n27209), .B(n28564), .C(\instr[16] ), 
         .Z(n2141)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i12518_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_2842_i28_3_lut_3_lut_4_lut (.A(n27209), .B(n28564), .C(n4075), 
         .D(\instr[31] ), .Z(n4707)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam mux_2842_i28_3_lut_3_lut_4_lut.init = 16'hf800;
    LUT4 i167_2_lut_rep_512_2_lut_3_lut (.A(n27209), .B(n28564), .C(n27212), 
         .Z(n27137)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i167_2_lut_rep_512_2_lut_3_lut.init = 16'h7070;
    LUT4 i4848_2_lut_rep_524_3_lut_4_lut (.A(n27209), .B(n28564), .C(n27211), 
         .D(n28563), .Z(n27149)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i4848_2_lut_rep_524_3_lut_4_lut.init = 16'h7770;
    LUT4 i23691_2_lut_rep_526_3_lut (.A(n27209), .B(n28564), .C(n28575), 
         .Z(n27151)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i23691_2_lut_rep_526_3_lut.init = 16'h8f8f;
    LUT4 i1_3_lut_3_lut_4_lut (.A(n27209), .B(n28564), .C(\instr[20] ), 
         .D(n27101), .Z(n22909)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i12217_2_lut_2_lut_3_lut (.A(n27209), .B(n28564), .C(mem_op_2__N_1384), 
         .Z(mem_op_increment_reg_de)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i12217_2_lut_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_3_lut_rep_557 (.A(n27197), .B(n27205), .C(n27198), .Z(n27182)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam i1_3_lut_rep_557.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut (.A(n27197), .B(n27205), .C(n27198), .D(n27186), 
         .Z(\alu_op_3__N_1337[2] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    LUT4 is_jalr_N_1372_bdd_2_lut_24167_3_lut (.A(n28563), .B(n27212), .C(n27211), 
         .Z(n26207)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam is_jalr_N_1372_bdd_2_lut_24167_3_lut.init = 16'h7070;
    LUT4 i2_2_lut_3_lut (.A(n28563), .B(n27212), .C(n27211), .Z(n10)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i2_2_lut_3_lut.init = 16'h8080;
    LUT4 i37_3_lut_3_lut (.A(n28563), .B(n27212), .C(n27211), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i37_3_lut_3_lut.init = 16'h7a7a;
    LUT4 i1_4_lut_4_lut_adj_301 (.A(n27179), .B(n23712), .C(n8274), .D(n26), 
         .Z(n23718)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_301.init = 16'h0400;
    LUT4 n27208_bdd_4_lut_24591_4_lut (.A(n27209), .B(n28564), .C(n27211), 
         .D(mem_op_2__N_1384), .Z(n27829)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam n27208_bdd_4_lut_24591_4_lut.init = 16'h808a;
    LUT4 i12716_4_lut_4_lut_4_lut (.A(n27204), .B(n27203), .C(n328[1]), 
         .D(n27153), .Z(n15_c)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!B))) */ ;
    defparam i12716_4_lut_4_lut_4_lut.init = 16'h00c4;
    LUT4 i1_4_lut_4_lut_adj_302 (.A(n27179), .B(n23756), .C(n8274), .D(n26), 
         .Z(n23762)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_302.init = 16'h0400;
    LUT4 i12531_3_lut_3_lut_4_lut (.A(n27204), .B(n27203), .C(n328[0]), 
         .D(n27153), .Z(n15_adj_2628)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;
    defparam i12531_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 i563_2_lut_rep_523_3_lut (.A(n27204), .B(n27203), .C(n27205), 
         .Z(n27148)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i563_2_lut_rep_523_3_lut.init = 16'h8080;
    LUT4 i12285_2_lut_3_lut_4_lut (.A(n27204), .B(n27203), .C(n28564), 
         .D(n27205), .Z(n14587)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12285_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i12787_2_lut_3_lut_4_lut (.A(n27204), .B(n27203), .C(n27153), 
         .D(n27205), .Z(n15_adj_2629)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i12787_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i559_4_lut_rep_496 (.A(n27211), .B(mem_op_2__N_1384), .C(n14503), 
         .D(n27205), .Z(n27121)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(93[13] 98[16])
    defparam i559_4_lut_rep_496.init = 16'h3b33;
    LUT4 i1_2_lut_4_lut_adj_303 (.A(n27211), .B(mem_op_2__N_1384), .C(n14503), 
         .D(n27205), .Z(n3_c)) /* synthesis lut_function=(A (B (C (D)))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(93[13] 98[16])
    defparam i1_2_lut_4_lut_adj_303.init = 16'hc400;
    LUT4 i1_4_lut_adj_304 (.A(n27175), .B(n23962), .C(n23956), .D(n24579), 
         .Z(is_ret_de)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_4_lut_adj_304.init = 16'h0080;
    LUT4 i1_4_lut_adj_305 (.A(n7), .B(n23944), .C(n27176), .D(n27201), 
         .Z(n23962)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_305.init = 16'h0004;
    LUT4 i1_3_lut_adj_306 (.A(n28563), .B(n27205), .C(n27146), .Z(n23956)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_adj_306.init = 16'h1010;
    LUT4 i22300_3_lut (.A(n27211), .B(n27204), .C(n27202), .Z(n24579)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i22300_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_adj_307 (.A(n27207), .B(n27209), .C(n27206), .Z(n23944)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_307.init = 16'h4040;
    LUT4 mux_55_i3_4_lut_4_lut (.A(n27179), .B(clk_c_enable_34), .C(additional_mem_ops_2__N_1129[2]), 
         .D(\additional_mem_ops[2] ), .Z(n4117)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;
    defparam mux_55_i3_4_lut_4_lut.init = 16'h7340;
    LUT4 i1_3_lut_rep_528_4_lut_4_lut (.A(n28564), .B(n27212), .C(n27211), 
         .D(n28563), .Z(n27153)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_3_lut_rep_528_4_lut_4_lut.init = 16'hfff7;
    LUT4 i5391_4_lut_4_lut (.A(n28564), .B(n155[3]), .C(n30), .D(n24128), 
         .Z(n7709)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5391_4_lut_4_lut.init = 16'hd850;
    LUT4 i23304_3_lut_4_lut_4_lut (.A(n28564), .B(n30_adj_8), .C(n27121), 
         .D(n28563), .Z(n7711)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i23304_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 i5387_4_lut_4_lut (.A(n28564), .B(n7601), .C(n30), .D(alu_op_3__N_1170[1]), 
         .Z(n7705)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5387_4_lut_4_lut.init = 16'hd850;
    LUT4 i4691_4_lut_4_lut (.A(n28564), .B(n7601), .C(n22000), .D(alu_op_3__N_1170[0]), 
         .Z(n6983)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i4691_4_lut_4_lut.init = 16'hd850;
    LUT4 i4693_4_lut_4_lut (.A(n28564), .B(n27156), .C(n27206), .D(n27121), 
         .Z(n6985)) /* synthesis lut_function=(A (D)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i4693_4_lut_4_lut.init = 16'hea40;
    LUT4 n1_bdd_3_lut_3_lut (.A(n28564), .B(n27212), .C(n28563), .Z(n26867)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam n1_bdd_3_lut_3_lut.init = 16'h1414;
    LUT4 n26208_bdd_3_lut_4_lut (.A(n27141), .B(n27174), .C(n28564), .D(n26208), 
         .Z(is_system_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam n26208_bdd_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_1900_i11_rep_80_3_lut_4_lut (.A(n27199), .B(n27143), .C(n27212), 
         .D(n27205), .Z(n2897)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(205[25] 214[32])
    defparam mux_1900_i11_rep_80_3_lut_4_lut.init = 16'hbfb0;
    LUT4 i1_2_lut_3_lut_adj_308 (.A(n27202), .B(n27146), .C(n22100), .Z(n22101)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_3_lut_adj_308.init = 16'he0e0;
    PFUMX instr_1__I_0_133_Mux_0_i15 (.BLUT(n23046), .ALUT(n22946), .C0(n27189), 
          .Z(n15)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 i1_4_lut_4_lut_adj_309 (.A(n27179), .B(n23768), .C(n8274), .D(n26), 
         .Z(n23774)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_309.init = 16'h0400;
    LUT4 i12421_2_lut_3_lut_4_lut (.A(n27202), .B(n27146), .C(n27128), 
         .D(n27185), .Z(is_jalr_N_1370)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i12421_2_lut_3_lut_4_lut.init = 16'he000;
    PFUMX i4692 (.BLUT(n15_adj_2628), .ALUT(n6983), .C0(n27209), .Z(alu_op_de[0]));
    PFUMX i5388 (.BLUT(n15_c), .ALUT(n7705), .C0(n25707), .Z(alu_op_de[1]));
    LUT4 n26873_bdd_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(\instr[30] ), .Z(n26874)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam n26873_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_2842_i17_3_lut_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(\instr[16] ), .Z(n4718)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_2842_i17_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_2842_i25_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[24] ), 
         .D(\instr[31] ), .Z(n4710)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_2842_i25_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_2842_i30_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[29] ), 
         .D(\instr[31] ), .Z(n4705)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_2842_i30_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_2842_i26_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[25] ), 
         .D(\instr[31] ), .Z(n4709)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_2842_i26_3_lut_4_lut.init = 16'hfe10;
    LUT4 n26289_bdd_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n26289), .Z(n26290)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam n26289_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_2842_i16_3_lut_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n27212), .Z(n4719)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_2842_i16_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1083_i11_rep_98_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n1741), .Z(n24641)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1083_i11_rep_98_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1083_i7_rep_92_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n1745), .Z(n24635)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1083_i7_rep_92_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i5390 (.BLUT(n15_adj_9), .ALUT(n23030), .C0(n25708), .Z(alu_op_de[2]));
    PFUMX i5392 (.BLUT(n22965), .ALUT(n7709), .C0(n25708), .Z(alu_op_de[3]));
    LUT4 mux_2842_i15_3_lut_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n28563), .Z(n4720)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_2842_i15_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n4069_bdd_3_lut_23868_4_lut (.A(n27143), .B(n27197), .C(\instr[19] ), 
         .D(\instr[31] ), .Z(n26296)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam n4069_bdd_3_lut_23868_4_lut.init = 16'hfe10;
    LUT4 i12444_2_lut_rep_498_3_lut_4_lut (.A(n27143), .B(n27197), .C(n27144), 
         .D(n27174), .Z(n27123)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;
    defparam i12444_2_lut_rep_498_3_lut_4_lut.init = 16'heee0;
    LUT4 n26277_bdd_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n26277), .Z(n26278)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam n26277_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_2842_i29_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[28] ), 
         .D(\instr[31] ), .Z(n4706)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_2842_i29_3_lut_4_lut.init = 16'hfe10;
    PFUMX i12908 (.BLUT(n15_adj_2629), .ALUT(n15222), .C0(n25708), .Z(is_alu_reg_de));
    LUT4 mux_1083_i8_rep_90_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n1744), .Z(n24633)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1083_i8_rep_90_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1083_i6_rep_84_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n1746), .Z(n24627)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1083_i6_rep_84_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5805_3_lut_4_lut (.A(n27143), .B(n27197), .C(n4075), .D(n27179), 
         .Z(n8123)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i5805_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_1083_i5_rep_82_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n1747), .Z(n24625)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1083_i5_rep_82_3_lut_4_lut.init = 16'hf1e0;
    PFUMX is_jalr_I_0 (.BLUT(is_jalr_N_1370), .ALUT(alu_op_3__N_1180), .C0(n27179), 
          .Z(is_jalr_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    PFUMX is_lui_I_0 (.BLUT(is_lui_N_1365), .ALUT(imm_31__N_1169), .C0(n27179), 
          .Z(is_lui_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 mux_2842_i14_3_lut_3_lut_4_lut (.A(n27143), .B(n27197), .C(\instr[31] ), 
         .D(n27211), .Z(n4721)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_2842_i14_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 is_store_I_0_4_lut (.A(n15143), .B(n27130), .C(n27179), .D(n27175), 
         .Z(is_store_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam is_store_I_0_4_lut.init = 16'h3a30;
    LUT4 i12833_4_lut (.A(n27209), .B(n28563), .C(n27211), .D(n27203), 
         .Z(n15143)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i12833_4_lut.init = 16'hcdcc;
    PFUMX i21 (.BLUT(n7_adj_2624), .ALUT(n8), .C0(n25126), .Z(is_load_de));
    LUT4 i1_4_lut_4_lut_adj_310 (.A(n27153), .B(n27182), .C(n27204), .D(n27203), 
         .Z(n22965)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i1_4_lut_4_lut_adj_310.init = 16'h1050;
    LUT4 i1_3_lut_4_lut_4_lut_adj_311 (.A(n27179), .B(n27185), .C(n28575), 
         .D(n27212), .Z(n23544)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_311.init = 16'h1000;
    LUT4 is_branch_I_0_4_lut (.A(n27184), .B(n27139), .C(n27179), .D(n27167), 
         .Z(is_branch_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam is_branch_I_0_4_lut.init = 16'h3a30;
    LUT4 additional_mem_ops_2__N_1132_0__bdd_3_lut (.A(n27203), .B(n27204), 
         .C(n27197), .Z(n26744)) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam additional_mem_ops_2__N_1132_0__bdd_3_lut.init = 16'h1515;
    LUT4 i1_4_lut_adj_312 (.A(n27199), .B(n22164), .C(n27201), .D(n27197), 
         .Z(n4057)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_312.init = 16'h0400;
    PFUMX instr_1__I_0_138_Mux_2_i31 (.BLUT(n15_adj_10), .ALUT(n30_adj_11), 
          .C0(n25707), .Z(additional_mem_ops_2__N_1129[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 i4942_4_lut_4_lut_4_lut (.A(n27143), .B(n27205), .C(n23598), 
         .D(n27109), .Z(n3166)) /* synthesis lut_function=(A (B ((D)+!C))+!A (B+!((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam i4942_4_lut_4_lut_4_lut.init = 16'hcc5c;
    PFUMX i24961 (.BLUT(n28566), .ALUT(n28567), .C0(mem_op_2__N_1384), 
          .Z(n28568));
    PFUMX is_jal_I_0 (.BLUT(is_jal_N_1374), .ALUT(alu_op_3__N_1181), .C0(n27179), 
          .Z(is_jal_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 n26784_bdd_3_lut_4_lut (.A(n27178), .B(n27212), .C(n27209), .D(n26783), 
         .Z(n26785)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam n26784_bdd_3_lut_4_lut.init = 16'hf101;
    LUT4 i12540_2_lut_4_lut (.A(n27170), .B(n7), .C(n27199), .D(n27211), 
         .Z(n19_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam i12540_2_lut_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_4_lut (.A(n27170), .B(n7), .C(n27199), .D(n27149), 
         .Z(n12)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam i2_2_lut_4_lut.init = 16'hfffe;
    LUT4 i12663_2_lut_3_lut_4_lut (.A(n27200), .B(n27172), .C(\instr[25] ), 
         .D(n27197), .Z(n4729)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam i12663_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i12665_2_lut_3_lut_4_lut (.A(n27200), .B(n27172), .C(\instr[27] ), 
         .D(n27197), .Z(n4727)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam i12665_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i12338_2_lut_3_lut_4_lut (.A(n27200), .B(n27172), .C(n27206), 
         .D(n27197), .Z(n4734)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam i12338_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i12662_2_lut_3_lut_4_lut (.A(n27200), .B(n27172), .C(n27203), 
         .D(n27197), .Z(n4730)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam i12662_2_lut_3_lut_4_lut.init = 16'hf0d0;
    PFUMX i24563 (.BLUT(n27834), .ALUT(n27829), .C0(n28564), .Z(\mem_op_de[1] ));
    LUT4 mux_1900_i17_3_lut_4_lut (.A(n27200), .B(n27172), .C(n27212), 
         .D(n27205), .Z(n2890)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_1900_i17_3_lut_4_lut.init = 16'h2f20;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n27179), .B(n23682), .C(n27114), 
         .D(n27108), .Z(n10_adj_12)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 mux_61_i1_3_lut_4_lut (.A(n27200), .B(n27172), .C(n27205), .D(n27169), 
         .Z(n328[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_61_i1_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_61_i2_3_lut_4_lut (.A(n27200), .B(n27172), .C(n27205), .D(n27197), 
         .Z(n328[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_61_i2_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i1_4_lut_4_lut_adj_313 (.A(n27179), .B(n23698), .C(n8274), .D(n26), 
         .Z(n23704)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_313.init = 16'h0400;
    LUT4 i12202_2_lut_3_lut_4_lut (.A(n27200), .B(n27173), .C(n27142), 
         .D(n27174), .Z(n14503)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i12202_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 instr_3__bdd_3_lut (.A(n27201), .B(n27198), .C(n27200), .Z(n26876)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam instr_3__bdd_3_lut.init = 16'hf7f7;
    LUT4 instr_3__bdd_4_lut (.A(n27199), .B(n27201), .C(n27198), .D(n27200), 
         .Z(n26877)) /* synthesis lut_function=(A+(B (C+!(D))+!B (D))) */ ;
    defparam instr_3__bdd_4_lut.init = 16'hfbee;
    LUT4 i1_4_lut_adj_314 (.A(n27211), .B(n27144), .C(n28563), .D(n24050), 
         .Z(mem_op_2__N_1384)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_314.init = 16'hffdf;
    LUT4 i1_3_lut_adj_315 (.A(n27199), .B(n27205), .C(n27201), .Z(n24050)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_315.init = 16'hfefe;
    LUT4 i1_2_lut_rep_504_4_lut (.A(n27204), .B(n27177), .C(n27203), .D(n27202), 
         .Z(n27129)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(282[33:52])
    defparam i1_2_lut_rep_504_4_lut.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module tinyqv_core
//

module tinyqv_core (n26927, \imm[0] , mstatus_mpie, clk_c, clk_c_enable_424, 
            n9675, n27218, time_hi, n27326, \debug_branch_N_446[31] , 
            tmp_data, load_done, clk_c_enable_71, n6982, instr_retired, 
            n14783, instr_complete_N_1647, n27367, n27369, n24404, 
            n27287, n27348, n15, cycle, \shift_amt[0] , n92, n5434, 
            n27279, clk_c_enable_73, \mie[14] , n926, \mie[13] , \mie[10] , 
            n893, \mie[9] , \mie[6] , n860, \mie[5] , \mie[2] , 
            n793, \mie[1] , cmp, \mepc[0] , \next_fsm_state_3__N_2499[3] , 
            cy, mstatus_mte, n26930, \imm[10] , n27374, n27305, 
            n27238, \addr_out[0] , \addr_out[1] , \next_pc_for_core[7] , 
            \next_pc_for_core[3] , counter_hi, \addr_out[23] , \addr_out[22] , 
            \addr_out[21] , \tmp_data[31] , alu_op, \tmp_data[30] , 
            \addr_out[20] , \addr_out[19] , \addr_out[18] , \addr_out[17] , 
            \next_pc_for_core[15] , \next_pc_for_core[11] , \addr_out[16] , 
            n27309, \imm[6] , \imm[2] , \addr_out[15] , \next_pc_for_core[23] , 
            \next_pc_for_core[19] , \addr_out[14] , \addr_out[13] , \addr_out[12] , 
            \addr_out[11] , \addr_out[10] , \addr_out[9] , \addr_out[8] , 
            \addr_out[7] , n27196, mstatus_mie, \addr_out[6] , \addr_out[5] , 
            \addr_out[4] , \addr_out[3] , n22121, \imm[1] , n27332, 
            interrupt_core, n27306, \csr_read_3__N_1443[0] , \csr_read_3__N_1451[0] , 
            n27292, \cycle_count_wide[0] , \instrret_count[0] , \debug_rd_3__N_405[28] , 
            \debug_rd_3__N_405[30] , \debug_rd_3__N_405[29] , \debug_rd_3__N_405[31] , 
            \next_pc_for_core[14] , \next_pc_for_core[10] , \time_count[2] , 
            mip_reg, clk_c_enable_350, n24216, n8162, \next_pc_for_core[22] , 
            \next_pc_for_core[18] , clk_c_enable_367, n26855, n27112, 
            n27106, n23738, n27109, n2123, n23798, n22721, n23750, 
            n22745, n23718, n22551, n24822, \debug_branch_N_442[28] , 
            n157, n23704, n22559, n23774, n22733, n23450, n22700, 
            n8, n23820, n26, n26345, n23690, n2322, n23810, n22715, 
            debug_rd_3__N_1575, load_top_bit_next_N_1731, mem_op, n24516, 
            n8274, n24, n23838, n23824, n3295, n23762, n22739, 
            \imm[4] , n27329, n24360, n23842, n12, n23848, n24601, 
            n24505, \a_for_shift_right[31] , data_rs1, n23894, n22784, 
            n23650, n27122, n23656, n27391, n23498, n23594, n27114, 
            n27108, n23598, n27110, rst_reg_n, n27342, load_top_bit, 
            data_out_3__N_1385, alu_a_in_3__N_1552, \debug_branch_N_442[29] , 
            \alu_a_in[1] , \debug_branch_N_840[29] , \timer_data[1] , 
            is_timer_addr, n27347, \mul_out[2] , \mul_out[3] , \mul_out[1] , 
            n27290, \ui_in_sync[1] , n1167, n27276, n27249, n27248, 
            n26686, n27302, n25069, n26049, clk_c_enable_276, debug_rd, 
            \shift_amt[1] , stall_core, n27263, is_load, n856, n22226, 
            clk_c_enable_423, n22898, any_additional_mem_ops, clk_c_enable_275, 
            accum, d_3__N_1868, \shift_out[1] , n27368, n27366, \imm[7] , 
            n7717, n26733, \debug_branch_N_450[0] , debug_instr_valid, 
            n27376, n27256, data_rs2, alu_b_in, is_auipc, is_jal, 
            n5160, n5171, n22499, n4575, n1766, \instr_write_offset_3__N_934[1] , 
            n1767, \instr_write_offset_3__N_934[0] , n27111, n27288, 
            n1768, pc_2__N_932, \mcause[1] , n616, \mcause[2] , \mcause[5] , 
            is_branch, is_jalr, is_system, is_alu_imm, is_alu_reg, 
            clk_c_enable_422, n15206, \debug_branch_N_450[3] , is_lui, 
            n27350, \debug_branch_N_442[31] , n27293, n27322, interrupt_pending_N_1671, 
            no_write_in_progress, n5168, \imm[3] , \imm[5] , n22178, 
            n26802, \imm[8] , \imm[9] , \debug_branch_N_442[30] , n26318, 
            n27338, n28573, n28571, n18, n27343, timer_interrupt, 
            n27349, n27362, n25142, n27231, n20, n14, n24838, 
            debug_rd_3__N_413, \tmp_data_in_3__N_1514[3] , n27274, \debug_rd_3__N_1567[0] , 
            debug_reg_wen_N_1692, \shift_out[0] , n25132, \pc[21] , 
            \pc[17] , n26200, \next_pc_for_core[20] , \next_pc_for_core[16] , 
            n225, \pc[23] , \pc[19] , n26175, \pc[20] , \pc[16] , 
            n225_adj_4, \next_pc_for_core[21] , \next_pc_for_core[17] , 
            n226, \pc[22] , \pc[18] , n26195, n26685, \data_out_slice[2] , 
            n27214, n27223, \mtimecmp[7] , mtimecmp_3__N_1935, n24772, 
            \debug_branch_N_446[29] , n27222, \mtimecmp[5] , mtimecmp_1__N_1941, 
            n27247, n27296, n27321, address_ready, n28575, n24775, 
            \debug_branch_N_446[30] , n26336, n26335, \addr_offset[2] , 
            n701, is_store, n24611, n26717, \debug_branch_N_450[2] , 
            n24774, \csr_read_3__N_1459[0] , n24616, \debug_branch_N_840[31] , 
            \data_out_slice[0] , \csr_read_3__N_1459[3] , n27023, \csr_read_3__N_1459[1] , 
            \cycle_count_wide[1] , \csr_read_3__N_1439[3] , n22090, \imm[11] , 
            n26976, instr_complete_N_1651, \time_count[3] , n5115, n26932, 
            \next_accum[5] , \next_accum[6] , \next_accum[7] , GND_net, 
            VCC_net, \next_accum[8] , \next_accum[9] , \next_accum[10] , 
            \next_accum[11] , \next_accum[12] , \next_accum[13] , \next_accum[14] , 
            \next_accum[15] , \next_accum[16] , \next_accum[17] , \next_accum[18] , 
            \next_accum[19] , \next_accum[4] , n62, n27377, n8157, 
            n8153, n7278, n25292, n63, \shift_amt[5] , rs1, rd, 
            rs2, return_addr, \reg_access[4][3] , n24605, \reg_access[3][2] , 
            n27205, n27113, n2356, cy_adj_5, \increment_result_3__N_1925[0] , 
            \instrret_count[3] , n27229, n27246, cy_adj_6, \increment_result_3__N_1911[1] , 
            \increment_result_3__N_1911[0] , \cycle_count_wide[6] , \cycle_count_wide[5] , 
            \cycle_count_wide[4] , \cycle_count_wide[3] , n27228, n27245, 
            n27180, n27187, n24124, n27188, n27252, n27215, n27154, 
            n27181, n23342, n27267, n27266, n27270) /* synthesis syn_module_defined=1 */ ;
    input n26927;
    input \imm[0] ;
    output mstatus_mpie;
    input clk_c;
    input clk_c_enable_424;
    input n9675;
    output n27218;
    output [2:0]time_hi;
    input n27326;
    input \debug_branch_N_446[31] ;
    output [31:0]tmp_data;
    output load_done;
    input clk_c_enable_71;
    input n6982;
    output instr_retired;
    input n14783;
    output instr_complete_N_1647;
    input n27367;
    input n27369;
    input n24404;
    output n27287;
    input n27348;
    output n15;
    output [1:0]cycle;
    output \shift_amt[0] ;
    input [3:0]n92;
    input n5434;
    output n27279;
    input clk_c_enable_73;
    output \mie[14] ;
    input n926;
    output \mie[13] ;
    output \mie[10] ;
    input n893;
    output \mie[9] ;
    output \mie[6] ;
    input n860;
    output \mie[5] ;
    output \mie[2] ;
    input n793;
    output \mie[1] ;
    output cmp;
    output \mepc[0] ;
    input \next_fsm_state_3__N_2499[3] ;
    output cy;
    output mstatus_mte;
    input n26930;
    input \imm[10] ;
    input n27374;
    input n27305;
    output n27238;
    output \addr_out[0] ;
    output \addr_out[1] ;
    input \next_pc_for_core[7] ;
    input \next_pc_for_core[3] ;
    input [4:2]counter_hi;
    output \addr_out[23] ;
    output \addr_out[22] ;
    output \addr_out[21] ;
    output \tmp_data[31] ;
    input [3:0]alu_op;
    output \tmp_data[30] ;
    output \addr_out[20] ;
    output \addr_out[19] ;
    output \addr_out[18] ;
    output \addr_out[17] ;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[11] ;
    output \addr_out[16] ;
    input n27309;
    input \imm[6] ;
    input \imm[2] ;
    output \addr_out[15] ;
    input \next_pc_for_core[23] ;
    input \next_pc_for_core[19] ;
    output \addr_out[14] ;
    output \addr_out[13] ;
    output \addr_out[12] ;
    output \addr_out[11] ;
    output \addr_out[10] ;
    output \addr_out[9] ;
    output \addr_out[8] ;
    output \addr_out[7] ;
    input n27196;
    output mstatus_mie;
    output \addr_out[6] ;
    output \addr_out[5] ;
    output \addr_out[4] ;
    output \addr_out[3] ;
    input n22121;
    input \imm[1] ;
    output n27332;
    input interrupt_core;
    input n27306;
    input \csr_read_3__N_1443[0] ;
    input \csr_read_3__N_1451[0] ;
    input n27292;
    output \cycle_count_wide[0] ;
    output \instrret_count[0] ;
    input \debug_rd_3__N_405[28] ;
    input \debug_rd_3__N_405[30] ;
    input \debug_rd_3__N_405[29] ;
    input \debug_rd_3__N_405[31] ;
    input \next_pc_for_core[14] ;
    input \next_pc_for_core[10] ;
    input \time_count[2] ;
    output [17:16]mip_reg;
    input clk_c_enable_350;
    input n24216;
    input n8162;
    input \next_pc_for_core[22] ;
    input \next_pc_for_core[18] ;
    input clk_c_enable_367;
    input n26855;
    output n27112;
    output n27106;
    input n23738;
    output n27109;
    output n2123;
    input n23798;
    output n22721;
    input n23750;
    output n22745;
    input n23718;
    output n22551;
    input n24822;
    input \debug_branch_N_442[28] ;
    input n157;
    input n23704;
    output n22559;
    input n23774;
    output n22733;
    input n23450;
    output n22700;
    input n8;
    input n23820;
    input n26;
    output n26345;
    input n23690;
    output n2322;
    input n23810;
    output n22715;
    input debug_rd_3__N_1575;
    output load_top_bit_next_N_1731;
    input [2:0]mem_op;
    input n24516;
    input n8274;
    input n24;
    output n23838;
    input n23824;
    output n3295;
    input n23762;
    output n22739;
    input \imm[4] ;
    output n27329;
    input n24360;
    input n23842;
    input n12;
    output n23848;
    input n24601;
    output n24505;
    output \a_for_shift_right[31] ;
    output [3:0]data_rs1;
    input n23894;
    output n22784;
    input n23650;
    input n27122;
    output n23656;
    input n27391;
    output n23498;
    input n23594;
    input n27114;
    output n27108;
    output n23598;
    input n27110;
    input rst_reg_n;
    input n27342;
    output load_top_bit;
    output data_out_3__N_1385;
    output alu_a_in_3__N_1552;
    input \debug_branch_N_442[29] ;
    output \alu_a_in[1] ;
    input \debug_branch_N_840[29] ;
    input \timer_data[1] ;
    input is_timer_addr;
    input n27347;
    input \mul_out[2] ;
    input \mul_out[3] ;
    input \mul_out[1] ;
    input n27290;
    input \ui_in_sync[1] ;
    output n1167;
    input n27276;
    input n27249;
    input n27248;
    input n26686;
    input n27302;
    input n25069;
    input n26049;
    input clk_c_enable_276;
    output [3:0]debug_rd;
    output \shift_amt[1] ;
    input stall_core;
    input n27263;
    input is_load;
    output n856;
    input n22226;
    output clk_c_enable_423;
    output n22898;
    input any_additional_mem_ops;
    output clk_c_enable_275;
    output [15:0]accum;
    output [19:0]d_3__N_1868;
    input \shift_out[1] ;
    input n27368;
    input n27366;
    input \imm[7] ;
    output n7717;
    input n26733;
    input \debug_branch_N_450[0] ;
    input debug_instr_valid;
    input n27376;
    input n27256;
    output [3:0]data_rs2;
    output [3:0]alu_b_in;
    input is_auipc;
    input is_jal;
    input n5160;
    output n5171;
    output n22499;
    input [1:0]n4575;
    input n1766;
    output \instr_write_offset_3__N_934[1] ;
    input n1767;
    output \instr_write_offset_3__N_934[0] ;
    output n27111;
    input n27288;
    input [1:0]n1768;
    output [1:0]pc_2__N_932;
    output \mcause[1] ;
    input n616;
    output \mcause[2] ;
    output \mcause[5] ;
    input is_branch;
    input is_jalr;
    input is_system;
    input is_alu_imm;
    input is_alu_reg;
    input clk_c_enable_422;
    input n15206;
    input \debug_branch_N_450[3] ;
    input is_lui;
    input n27350;
    input \debug_branch_N_442[31] ;
    output n27293;
    output n27322;
    output interrupt_pending_N_1671;
    input no_write_in_progress;
    output n5168;
    input \imm[3] ;
    input \imm[5] ;
    output n22178;
    input n26802;
    input \imm[8] ;
    input \imm[9] ;
    input \debug_branch_N_442[30] ;
    input n26318;
    output n27338;
    input n28573;
    input n28571;
    output n18;
    output n27343;
    input timer_interrupt;
    output n27349;
    input n27362;
    output n25142;
    input n27231;
    input n20;
    input n14;
    input n24838;
    input debug_rd_3__N_413;
    input \tmp_data_in_3__N_1514[3] ;
    input n27274;
    input \debug_rd_3__N_1567[0] ;
    input debug_reg_wen_N_1692;
    input \shift_out[0] ;
    input n25132;
    input \pc[21] ;
    input \pc[17] ;
    output n26200;
    input \next_pc_for_core[20] ;
    input \next_pc_for_core[16] ;
    output n225;
    input \pc[23] ;
    input \pc[19] ;
    output n26175;
    input \pc[20] ;
    input \pc[16] ;
    output n225_adj_4;
    input \next_pc_for_core[21] ;
    input \next_pc_for_core[17] ;
    output n226;
    input \pc[22] ;
    input \pc[18] ;
    output n26195;
    output n26685;
    output \data_out_slice[2] ;
    output n27214;
    input n27223;
    input \mtimecmp[7] ;
    output mtimecmp_3__N_1935;
    input n24772;
    input \debug_branch_N_446[29] ;
    output n27222;
    input \mtimecmp[5] ;
    output mtimecmp_1__N_1941;
    input n27247;
    input n27296;
    input n27321;
    output address_ready;
    input n28575;
    input n24775;
    input \debug_branch_N_446[30] ;
    input n26336;
    input n26335;
    input \addr_offset[2] ;
    output n701;
    input is_store;
    input n24611;
    input n26717;
    input \debug_branch_N_450[2] ;
    input n24774;
    input \csr_read_3__N_1459[0] ;
    input n24616;
    input \debug_branch_N_840[31] ;
    output \data_out_slice[0] ;
    input \csr_read_3__N_1459[3] ;
    output n27023;
    input \csr_read_3__N_1459[1] ;
    output \cycle_count_wide[1] ;
    input \csr_read_3__N_1439[3] ;
    input n22090;
    input \imm[11] ;
    input n26976;
    input instr_complete_N_1651;
    input \time_count[3] ;
    input n5115;
    output n26932;
    input \next_accum[5] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input GND_net;
    input VCC_net;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[4] ;
    output n62;
    input n27377;
    output n8157;
    output n8153;
    output n7278;
    input n25292;
    input n63;
    output \shift_amt[5] ;
    input [3:0]rs1;
    input [3:0]rd;
    input [3:0]rs2;
    output [23:1]return_addr;
    output \reg_access[4][3] ;
    input n24605;
    output \reg_access[3][2] ;
    input n27205;
    input n27113;
    output n2356;
    output cy_adj_5;
    input \increment_result_3__N_1925[0] ;
    output \instrret_count[3] ;
    input n27229;
    input n27246;
    output cy_adj_6;
    input \increment_result_3__N_1911[1] ;
    input \increment_result_3__N_1911[0] ;
    output \cycle_count_wide[6] ;
    output \cycle_count_wide[5] ;
    output \cycle_count_wide[4] ;
    output \cycle_count_wide[3] ;
    input n27228;
    input n27245;
    output n27180;
    input n27187;
    input n24124;
    input n27188;
    input n27252;
    input n27215;
    input n27154;
    input n27181;
    input n23342;
    input n27267;
    input n27266;
    input n27270;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n26928, n26929, clk_c_enable_3, n5545;
    wire [23:0]mepc;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(68[16:20])
    wire [3:0]n658;
    wire [16:0]mie;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(323[16:19])
    
    wire clk_c_enable_91, n26533;
    wire [2:0]n1;
    
    wire n27474, n25072, n27475, clk_c_enable_321, n9673;
    wire [3:0]tmp_data_in_3__N_1514;
    
    wire n652;
    wire [3:0]debug_rd_3__N_1563;
    wire [3:0]n196;
    
    wire n26059, clk_c_enable_68, n20944, clk_c_enable_289, is_double_fault_r;
    wire [2:0]n498;
    
    wire clk_c_enable_74, n21486, clk_c_enable_78, n21490, n21454, 
        n928, clk_c_enable_83, n21488, n21452, n895, clk_c_enable_87, 
        n21484, n21450, n862, n21482, n26328, cmp_out;
    wire [31:0]tmp_data_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(88[16:24])
    wire [1:0]last_interrupt_req;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(417[15:33])
    
    wire clk_c_enable_345, cy_out, clk_c_enable_101, mstatus_mte_N_1703, 
        n26931;
    wire [31:0]a_for_shift_right;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[17:34])
    
    wire n27230, n27472, n27280, n24607, n27471, n27408, n27407, 
        n27235;
    wire [3:0]n5123;
    wire [3:0]n5155;
    wire [5:0]mcause;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(325[15:21])
    
    wire n27414, n27413, n5215, n25081;
    wire [6:0]cycle_count_wide;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(279[16:32])
    wire [3:0]instrret_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(301[16:30])
    
    wire n26968, n24800, n22788, instr_complete_N_1652, n26977, n8786, 
        n23213, n27489, n27415, n26978, n26979, n27021;
    wire [3:0]n191;
    wire [3:0]debug_rd_3__N_1559;
    wire [1:0]n979;
    wire [3:0]csr_read_3__N_1455;
    
    wire n27022, n27019, n27409, n27020, n27488;
    wire [5:0]n611;
    
    wire n4521;
    wire [3:0]alu_a_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[16:24])
    
    wire n24242, n27195, clk_c_enable_421, n19988, n24034;
    wire [3:0]n653;
    
    wire n14470, n26060, n26061, n27346;
    wire [3:0]alu_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(110[16:23])
    
    wire n26684;
    wire [1:0]n948;
    
    wire n5;
    wire [1:0]n822;
    
    wire n27490;
    wire [1:0]n809;
    
    wire n26327, n26343, n26687, n26341, n26342, n27473, n28360, 
        n28358, n26360, n26062, debug_rd_3__N_1400;
    wire [4:0]shift_amt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(124[15:24])
    
    wire clk_c_enable_290, n23326, n26359;
    wire [3:0]tmp_data_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(242[15:26])
    
    wire n46, n25053;
    wire [3:0]debug_rd_3__N_1571;
    
    wire n7590, debug_reg_wen_N_1689;
    wire [3:0]csr_read_3__N_1447;
    
    wire n24410, n27242, n27278, alu_b_in_3__N_1504, instr_complete_N_1656, 
        instr_complete_N_1654, n24801, instr_complete_N_1648, n23264, 
        n27308, n24018, n24014, mstatus_mie_N_1707, debug_rd_3__N_1401, 
        n26532, n23318, n24789;
    wire [3:0]tmp_data_in_3__N_1582;
    wire [16:0]interrupt_pending_N_1672;
    wire [2:0]n4674;
    
    wire n28580, n23101;
    wire [3:0]n234;
    
    wire n27491, n5_adj_2620, mstatus_mie_N_1709;
    wire [3:0]debug_rd_3__N_1396;
    wire [3:0]debug_rd_3__N_1392;
    
    wire instr_complete_N_1650, instr_complete_N_1649, debug_reg_wen, 
        n25119;
    wire [65:0]dr_3__N_1864;
    
    wire n28361, n28359, n27234;
    wire [3:0]debug_rd_3__N_1567;
    
    wire n28581, n8197, n24290, n24787, n24788, n24799;
    wire [3:0]mul_out_3__N_1510;
    
    wire n26482, n26484;
    wire [3:0]n4528;
    
    PFUMX i24240 (.BLUT(n26928), .ALUT(n26927), .C0(\imm[0] ), .Z(n26929));
    FD1P3AX mstatus_mpie_525 (.D(n5545), .SP(clk_c_enable_3), .CK(clk_c), 
            .Q(mstatus_mpie)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam mstatus_mpie_525.GSR = "DISABLED";
    FD1P3IX mepc_i0_i21 (.D(n658[1]), .SP(clk_c_enable_424), .CD(n9675), 
            .CK(clk_c), .Q(mepc[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i21.GSR = "DISABLED";
    FD1P3IX mie__i0 (.D(n26533), .SP(clk_c_enable_91), .CD(n27218), .CK(clk_c), 
            .Q(mie[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i0.GSR = "DISABLED";
    FD1P3IX mepc_i0_i20 (.D(n658[0]), .SP(clk_c_enable_424), .CD(n9675), 
            .CK(clk_c), .Q(mepc[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i20.GSR = "DISABLED";
    FD1S3IX time_hi__i0 (.D(n1[0]), .CK(clk_c), .CD(n27326), .Q(time_hi[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i0.GSR = "DISABLED";
    PFUMX i24383 (.BLUT(n27474), .ALUT(\debug_branch_N_446[31] ), .C0(n25072), 
          .Z(n27475));
    FD1P3IX tmp_data_i0_i29 (.D(tmp_data_in_3__N_1514[1]), .SP(clk_c_enable_321), 
            .CD(n9673), .CK(clk_c), .Q(tmp_data[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i29.GSR = "DISABLED";
    FD1P3AX load_done_515 (.D(n6982), .SP(clk_c_enable_71), .CK(clk_c), 
            .Q(load_done)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(232[12] 235[8])
    defparam load_done_515.GSR = "DISABLED";
    FD1S3IX instr_retired_518 (.D(instr_complete_N_1647), .CK(clk_c), .CD(n14783), 
            .Q(instr_retired)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(303[12] 305[8])
    defparam instr_retired_518.GSR = "DISABLED";
    FD1P3IX tmp_data_i0_i28 (.D(tmp_data_in_3__N_1514[0]), .SP(clk_c_enable_321), 
            .CD(n9673), .CK(clk_c), .Q(tmp_data[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i28.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n27367), .B(n27369), .C(n24404), .D(n27287), 
         .Z(n652)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[25:55])
    defparam i1_3_lut_4_lut.init = 16'h0080;
    LUT4 debug_rd_3__N_1567_1__bdd_4_lut_24171_4_lut (.A(n27348), .B(n15), 
         .C(debug_rd_3__N_1563[1]), .D(n196[1]), .Z(n26059)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam debug_rd_3__N_1567_1__bdd_4_lut_24171_4_lut.init = 16'he4a0;
    FD1P3IX cycle__i1 (.D(n20944), .SP(clk_c_enable_68), .CD(n27326), 
            .CK(clk_c), .Q(cycle[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam cycle__i1.GSR = "DISABLED";
    FD1P3AX shift_amt__i1 (.D(n92[0]), .SP(clk_c_enable_289), .CK(clk_c), 
            .Q(\shift_amt[0] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i1.GSR = "DISABLED";
    FD1P3IX is_double_fault_r_520 (.D(n27279), .SP(clk_c_enable_71), .CD(n5434), 
            .CK(clk_c), .Q(is_double_fault_r)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(361[12] 364[8])
    defparam is_double_fault_r_520.GSR = "DISABLED";
    FD1P3IX time_hi__i2 (.D(n498[2]), .SP(clk_c_enable_73), .CD(n27326), 
            .CK(clk_c), .Q(time_hi[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i2.GSR = "DISABLED";
    FD1P3IX time_hi__i1 (.D(n498[1]), .SP(clk_c_enable_73), .CD(n27326), 
            .CK(clk_c), .Q(time_hi[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i1.GSR = "DISABLED";
    FD1P3IX mie__i16 (.D(n21486), .SP(clk_c_enable_74), .CD(n27218), .CK(clk_c), 
            .Q(mie[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i16.GSR = "DISABLED";
    FD1P3IX mie__i15 (.D(n21490), .SP(clk_c_enable_78), .CD(n27218), .CK(clk_c), 
            .Q(mie[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i15.GSR = "DISABLED";
    FD1P3IX mie__i14 (.D(n926), .SP(clk_c_enable_78), .CD(n27218), .CK(clk_c), 
            .Q(\mie[14] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i14.GSR = "DISABLED";
    FD1P3IX mie__i13 (.D(n21454), .SP(clk_c_enable_78), .CD(n27218), .CK(clk_c), 
            .Q(\mie[13] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i13.GSR = "DISABLED";
    FD1P3IX mie__i12 (.D(n928), .SP(clk_c_enable_78), .CD(n27218), .CK(clk_c), 
            .Q(mie[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i12.GSR = "DISABLED";
    FD1P3IX mie__i11 (.D(n21488), .SP(clk_c_enable_83), .CD(n27218), .CK(clk_c), 
            .Q(mie[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i11.GSR = "DISABLED";
    FD1P3IX mie__i10 (.D(n893), .SP(clk_c_enable_83), .CD(n27218), .CK(clk_c), 
            .Q(\mie[10] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i10.GSR = "DISABLED";
    FD1P3IX mie__i9 (.D(n21452), .SP(clk_c_enable_83), .CD(n27218), .CK(clk_c), 
            .Q(\mie[9] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i9.GSR = "DISABLED";
    FD1P3IX mie__i8 (.D(n895), .SP(clk_c_enable_83), .CD(n27218), .CK(clk_c), 
            .Q(mie[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i8.GSR = "DISABLED";
    FD1P3IX mie__i7 (.D(n21484), .SP(clk_c_enable_87), .CD(n27218), .CK(clk_c), 
            .Q(mie[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i7.GSR = "DISABLED";
    FD1P3IX mie__i6 (.D(n860), .SP(clk_c_enable_87), .CD(n27218), .CK(clk_c), 
            .Q(\mie[6] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i6.GSR = "DISABLED";
    FD1P3IX mie__i5 (.D(n21450), .SP(clk_c_enable_87), .CD(n27218), .CK(clk_c), 
            .Q(\mie[5] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i5.GSR = "DISABLED";
    FD1P3IX mie__i4 (.D(n862), .SP(clk_c_enable_87), .CD(n27218), .CK(clk_c), 
            .Q(mie[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i4.GSR = "DISABLED";
    FD1P3IX mie__i3 (.D(n21482), .SP(clk_c_enable_91), .CD(n27218), .CK(clk_c), 
            .Q(mie[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i3.GSR = "DISABLED";
    FD1P3IX mie__i2 (.D(n793), .SP(clk_c_enable_91), .CD(n27218), .CK(clk_c), 
            .Q(\mie[2] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i2.GSR = "DISABLED";
    FD1P3IX mie__i1 (.D(n26328), .SP(clk_c_enable_91), .CD(n27218), .CK(clk_c), 
            .Q(\mie[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i1.GSR = "DISABLED";
    FD1S3AX cmp_511 (.D(cmp_out), .CK(clk_c), .Q(cmp)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(117[12] 120[8])
    defparam cmp_511.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i0 (.D(tmp_data_c[4]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i0.GSR = "DISABLED";
    FD1P3AX mepc_i0_i0 (.D(mepc[4]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(\mepc[0] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i0.GSR = "DISABLED";
    FD1P3AX last_interrupt_req_i0_i0 (.D(\next_fsm_state_3__N_2499[3] ), .SP(clk_c_enable_345), 
            .CK(clk_c), .Q(last_interrupt_req[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam last_interrupt_req_i0_i0.GSR = "DISABLED";
    FD1S3AX cy_510 (.D(cy_out), .CK(clk_c), .Q(cy)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(117[12] 120[8])
    defparam cy_510.GSR = "DISABLED";
    FD1P3BX mstatus_mte_523 (.D(mstatus_mte_N_1703), .SP(clk_c_enable_101), 
            .CK(clk_c), .PD(n27326), .Q(mstatus_mte)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(384[18] 390[12])
    defparam mstatus_mte_523.GSR = "DISABLED";
    LUT4 n26930_bdd_3_lut (.A(n26930), .B(n26929), .C(\imm[10] ), .Z(n26931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26930_bdd_3_lut.init = 16'hcaca;
    LUT4 tmp_data_31__I_0_542_i3_3_lut_rep_613_4_lut (.A(n27374), .B(n27305), 
         .C(mepc[2]), .D(tmp_data_c[6]), .Z(n27238)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i3_3_lut_rep_613_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i1_3_lut_4_lut (.A(n27374), .B(n27305), .C(\mepc[0] ), 
         .D(tmp_data_c[4]), .Z(\addr_out[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i2_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[1]), 
         .D(tmp_data_c[5]), .Z(\addr_out[1] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 debug_branch_N_446_31__bdd_3_lut (.A(\next_pc_for_core[7] ), .B(\next_pc_for_core[3] ), 
         .C(counter_hi[2]), .Z(n27474)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam debug_branch_N_446_31__bdd_3_lut.init = 16'hacac;
    LUT4 tmp_data_31__I_0_542_i24_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[23]), 
         .D(tmp_data_c[27]), .Z(\addr_out[23] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i23_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[22]), 
         .D(tmp_data_c[26]), .Z(\addr_out[22] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i22_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[21]), 
         .D(tmp_data_c[25]), .Z(\addr_out[21] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 i10330_3_lut (.A(\tmp_data[31] ), .B(tmp_data_c[0]), .C(alu_op[2]), 
         .Z(a_for_shift_right[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    defparam i10330_3_lut.init = 16'hcaca;
    LUT4 i10339_3_lut (.A(\tmp_data[30] ), .B(tmp_data_c[1]), .C(alu_op[2]), 
         .Z(a_for_shift_right[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    defparam i10339_3_lut.init = 16'hcaca;
    LUT4 tmp_data_31__I_0_542_i21_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[20]), 
         .D(tmp_data_c[24]), .Z(\addr_out[20] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 n27230_bdd_4_lut_24353 (.A(n27230), .B(counter_hi[4]), .C(counter_hi[2]), 
         .D(counter_hi[3]), .Z(clk_c_enable_78)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam n27230_bdd_4_lut_24353.init = 16'h4000;
    LUT4 tmp_data_31__I_0_542_i20_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[19]), 
         .D(tmp_data_c[23]), .Z(\addr_out[19] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i19_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[18]), 
         .D(tmp_data_c[22]), .Z(\addr_out[18] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i18_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[17]), 
         .D(tmp_data_c[21]), .Z(\addr_out[17] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 next_pc_for_core_23__bdd_3_lut (.A(\next_pc_for_core[15] ), .B(\next_pc_for_core[11] ), 
         .C(counter_hi[2]), .Z(n27472)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam next_pc_for_core_23__bdd_3_lut.init = 16'hacac;
    LUT4 tmp_data_31__I_0_542_i17_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[16]), 
         .D(tmp_data_c[20]), .Z(\addr_out[16] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 i22326_4_lut (.A(n27309), .B(n27280), .C(\imm[6] ), .D(\imm[2] ), 
         .Z(n24607)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22326_4_lut.init = 16'hfffe;
    LUT4 tmp_data_31__I_0_542_i16_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[15]), 
         .D(tmp_data_c[19]), .Z(\addr_out[15] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 next_pc_for_core_23__bdd_4_lut (.A(\next_pc_for_core[23] ), .B(\next_pc_for_core[19] ), 
         .C(counter_hi[3]), .D(counter_hi[2]), .Z(n27471)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam next_pc_for_core_23__bdd_4_lut.init = 16'h0a0c;
    LUT4 tmp_data_31__I_0_542_i15_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[14]), 
         .D(tmp_data_c[18]), .Z(\addr_out[14] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 n27230_bdd_4_lut (.A(n27230), .B(counter_hi[3]), .C(counter_hi[4]), 
         .D(counter_hi[2]), .Z(clk_c_enable_83)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam n27230_bdd_4_lut.init = 16'h0040;
    LUT4 mux_3193_i3_4_lut_then_4_lut (.A(mepc[2]), .B(\imm[6] ), .C(counter_hi[2]), 
         .D(counter_hi[4]), .Z(n27408)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3193_i3_4_lut_then_4_lut.init = 16'h3088;
    LUT4 mux_3193_i3_4_lut_else_4_lut (.A(mepc[2]), .B(\imm[6] ), .C(counter_hi[2]), 
         .D(counter_hi[4]), .Z(n27407)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3193_i3_4_lut_else_4_lut.init = 16'h888b;
    LUT4 tmp_data_31__I_0_542_i14_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[13]), 
         .D(tmp_data_c[17]), .Z(\addr_out[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i13_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[12]), 
         .D(tmp_data_c[16]), .Z(\addr_out[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i12_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[11]), 
         .D(tmp_data_c[15]), .Z(\addr_out[11] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i11_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[10]), 
         .D(tmp_data_c[14]), .Z(\addr_out[10] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i10_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[9]), 
         .D(tmp_data_c[13]), .Z(\addr_out[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i9_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[8]), 
         .D(tmp_data_c[12]), .Z(\addr_out[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i8_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[7]), 
         .D(tmp_data_c[11]), .Z(\addr_out[7] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 i12146_4_lut (.A(n27196), .B(n27218), .C(mstatus_mie), .D(n27235), 
         .Z(n5545)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam i12146_4_lut.init = 16'h3022;
    LUT4 tmp_data_31__I_0_542_i7_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[6]), 
         .D(tmp_data_c[10]), .Z(\addr_out[6] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i6_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[5]), 
         .D(tmp_data_c[9]), .Z(\addr_out[5] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i5_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[4]), 
         .D(tmp_data_c[8]), .Z(\addr_out[4] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i4_3_lut_4_lut (.A(n27374), .B(n27305), .C(mepc[3]), 
         .D(tmp_data_c[7]), .Z(\addr_out[3] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_3203_i2_4_lut (.A(n5123[1]), .B(mepc[1]), .C(\imm[0] ), .D(n22121), 
         .Z(n5155[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3203_i2_4_lut.init = 16'hca0a;
    LUT4 i12446_4_lut_then_4_lut (.A(\imm[1] ), .B(mcause[4]), .C(counter_hi[4]), 
         .D(counter_hi[3]), .Z(n27414)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i12446_4_lut_then_4_lut.init = 16'h0008;
    LUT4 i12446_4_lut_else_4_lut (.A(mcause[0]), .B(\imm[1] ), .C(counter_hi[4]), 
         .D(counter_hi[3]), .Z(n27413)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i12446_4_lut_else_4_lut.init = 16'h0008;
    LUT4 i23653_2_lut_3_lut_4_lut (.A(n27332), .B(n27305), .C(n5215), 
         .D(interrupt_core), .Z(n25081)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i23653_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 time_count_2__bdd_3_lut (.A(cycle_count_wide[2]), .B(\imm[1] ), 
         .C(instrret_count[2]), .Z(n26968)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam time_count_2__bdd_3_lut.init = 16'he2e2;
    LUT4 tmp_data_in_3__N_1581_I_0_588_2_lut_rep_610_3_lut_4_lut (.A(n27332), 
         .B(n27305), .C(n27306), .D(interrupt_core), .Z(n27235)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C)+!B (C+!(D))))) */ ;
    defparam tmp_data_in_3__N_1581_I_0_588_2_lut_rep_610_3_lut_4_lut.init = 16'h0f04;
    LUT4 i7326_2_lut_3_lut_4_lut (.A(n27332), .B(n27305), .C(clk_c_enable_321), 
         .D(interrupt_core), .Z(n9673)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i7326_2_lut_3_lut_4_lut.init = 16'hf040;
    PFUMX i22457 (.BLUT(\csr_read_3__N_1443[0] ), .ALUT(\csr_read_3__N_1451[0] ), 
          .C0(\imm[6] ), .Z(n24800));
    LUT4 instr_complete_I_134_4_lut (.A(cycle[0]), .B(n27369), .C(n27292), 
         .D(n22788), .Z(instr_complete_N_1652)) /* synthesis lut_function=(A (B+((D)+!C))+!A !(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(226[34:58])
    defparam instr_complete_I_134_4_lut.init = 16'haa9a;
    LUT4 csr_read_3__N_1463_1__bdd_3_lut_24293 (.A(\cycle_count_wide[0] ), 
         .B(\instrret_count[0] ), .C(\imm[1] ), .Z(n26977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam csr_read_3__N_1463_1__bdd_3_lut_24293.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n8786), .B(n27279), .C(\debug_rd_3__N_405[28] ), 
         .D(interrupt_core), .Z(n23213)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut.init = 16'h0004;
    LUT4 i1_3_lut (.A(\debug_rd_3__N_405[30] ), .B(\debug_rd_3__N_405[29] ), 
         .C(\debug_rd_3__N_405[31] ), .Z(n8786)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(353[26:40])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 next_pc_for_core_22__bdd_3_lut_24547 (.A(\next_pc_for_core[14] ), 
         .B(\next_pc_for_core[10] ), .C(counter_hi[2]), .Z(n27489)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam next_pc_for_core_22__bdd_3_lut_24547.init = 16'hacac;
    LUT4 n5145_bdd_3_lut (.A(n27415), .B(n26978), .C(\imm[10] ), .Z(n26979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n5145_bdd_3_lut.init = 16'hcaca;
    LUT4 n8162_bdd_4_lut (.A(\time_count[2] ), .B(n26968), .C(\imm[0] ), 
         .D(\imm[1] ), .Z(n27021)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C)+!B))) */ ;
    defparam n8162_bdd_4_lut.init = 16'h0cac;
    LUT4 i23242_4_lut_4_lut (.A(n27348), .B(n15), .C(n196[0]), .D(n191[0]), 
         .Z(debug_rd_3__N_1559[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;
    defparam i23242_4_lut_4_lut.init = 16'hf4b0;
    FD1P3IX mip_reg__i16 (.D(n979[0]), .SP(clk_c_enable_350), .CD(n27218), 
            .CK(clk_c), .Q(mip_reg[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mip_reg__i16.GSR = "DISABLED";
    LUT4 csr_read_3__I_128_i4_4_lut (.A(mcause[3]), .B(n24216), .C(n27306), 
         .D(n27309), .Z(csr_read_3__N_1455[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(490[33] 493[57])
    defparam csr_read_3__I_128_i4_4_lut.init = 16'hca0a;
    LUT4 n8162_bdd_3_lut (.A(n8162), .B(n27021), .C(\imm[10] ), .Z(n27022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n8162_bdd_3_lut.init = 16'hcaca;
    LUT4 n27019_bdd_3_lut (.A(n27019), .B(n27409), .C(\imm[0] ), .Z(n27020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27019_bdd_3_lut.init = 16'hcaca;
    LUT4 next_pc_for_core_22__bdd_4_lut_24546 (.A(\next_pc_for_core[22] ), 
         .B(\next_pc_for_core[18] ), .C(counter_hi[3]), .D(counter_hi[2]), 
         .Z(n27488)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam next_pc_for_core_22__bdd_4_lut_24546.init = 16'h0a0c;
    FD1P3IX mcause__i0 (.D(n611[0]), .SP(clk_c_enable_367), .CD(n27326), 
            .CK(clk_c), .Q(mcause[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i0.GSR = "DISABLED";
    LUT4 n5135_bdd_3_lut (.A(n26855), .B(n4521), .C(\imm[6] ), .Z(n27019)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam n5135_bdd_3_lut.init = 16'h0808;
    LUT4 i2841_4_lut_4_lut_4_lut (.A(n27112), .B(n27106), .C(n23738), 
         .D(n27109), .Z(n2123)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i2841_4_lut_4_lut_4_lut.init = 16'hffbf;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n27112), .B(n27106), .C(n23798), .D(n27109), 
         .Z(n22721)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_242 (.A(n27112), .B(n27106), .C(n23750), 
         .D(n27109), .Z(n22745)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_242.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_243 (.A(n27112), .B(n27106), .C(n23718), 
         .D(n27109), .Z(n22551)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_243.init = 16'h0040;
    LUT4 i12200_4_lut_4_lut (.A(n27348), .B(n24822), .C(\debug_branch_N_442[28] ), 
         .D(n157), .Z(alu_a_in[0])) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam i12200_4_lut_4_lut.init = 16'h5410;
    LUT4 i1_4_lut_4_lut_4_lut_adj_244 (.A(n27112), .B(n27106), .C(n23704), 
         .D(n27109), .Z(n22559)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_244.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_245 (.A(n27112), .B(n27106), .C(n23774), 
         .D(n27109), .Z(n22733)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_245.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_246 (.A(n27112), .B(n27106), .C(n23450), 
         .D(n27109), .Z(n22700)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_246.init = 16'h0040;
    LUT4 i23474_4_lut (.A(n27218), .B(n24242), .C(n27195), .D(n8), .Z(clk_c_enable_421)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i23474_4_lut.init = 16'hfbfa;
    LUT4 n10_bdd_4_lut_23982_4_lut (.A(n27112), .B(n23820), .C(n26), .D(n27106), 
         .Z(n26345)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam n10_bdd_4_lut_23982_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_4_lut_4_lut_adj_247 (.A(n27112), .B(n27106), .C(n23690), 
         .D(n27109), .Z(n2322)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_247.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_248 (.A(n27112), .B(n27106), .C(n23810), 
         .D(n27109), .Z(n22715)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_248.init = 16'h0040;
    LUT4 i1_4_lut_adj_249 (.A(n19988), .B(debug_rd_3__N_1575), .C(counter_hi[4]), 
         .D(n24034), .Z(load_top_bit_next_N_1731)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_249.init = 16'h0400;
    LUT4 i17774_2_lut (.A(counter_hi[3]), .B(mem_op[0]), .Z(n19988)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17774_2_lut.init = 16'h6666;
    LUT4 i1_3_lut_adj_250 (.A(mem_op[2]), .B(mem_op[1]), .C(counter_hi[2]), 
         .Z(n24034)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_adj_250.init = 16'h1010;
    LUT4 i1_4_lut_4_lut (.A(n27112), .B(n24516), .C(n8274), .D(n24), 
         .Z(n23838)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_4_lut_4_lut_adj_251 (.A(n27112), .B(n27106), .C(n23824), 
         .D(n27109), .Z(n3295)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_251.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_252 (.A(n27112), .B(n27106), .C(n23762), 
         .D(n27109), .Z(n22739)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_252.init = 16'h0040;
    LUT4 i1_3_lut_rep_655_4_lut (.A(\imm[4] ), .B(n27329), .C(n24360), 
         .D(n27374), .Z(n27280)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i1_3_lut_rep_655_4_lut.init = 16'hfeff;
    LUT4 i1_4_lut_4_lut_adj_253 (.A(n27112), .B(n23842), .C(n12), .D(n8274), 
         .Z(n23848)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_253.init = 16'h0040;
    LUT4 i10344_3_lut (.A(tmp_data_c[1]), .B(\tmp_data[30] ), .C(alu_op[2]), 
         .Z(a_for_shift_right[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    defparam i10344_3_lut.init = 16'hcaca;
    LUT4 i22229_4_lut_4_lut_4_lut (.A(n27112), .B(n27106), .C(n24601), 
         .D(n27109), .Z(n24505)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i22229_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i10331_3_lut (.A(tmp_data_c[0]), .B(\tmp_data[31] ), .C(alu_op[2]), 
         .Z(\a_for_shift_right[31] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    defparam i10331_3_lut.init = 16'hcaca;
    LUT4 i10351_3_lut (.A(tmp_data_c[2]), .B(tmp_data[29]), .C(alu_op[2]), 
         .Z(a_for_shift_right[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    defparam i10351_3_lut.init = 16'hcaca;
    LUT4 mux_251_i4_3_lut (.A(mepc[3]), .B(data_rs1[3]), .C(n652), .Z(n653[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i4_3_lut.init = 16'hcaca;
    LUT4 mux_251_i1_3_lut (.A(\mepc[0] ), .B(data_rs1[0]), .C(n652), .Z(n653[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_4_lut_adj_254 (.A(n27112), .B(n27106), .C(n23894), 
         .D(n27109), .Z(n22784)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_254.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_255 (.A(n27112), .B(n23650), .C(n27122), .D(n8274), 
         .Z(n23656)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_255.init = 16'h0040;
    LUT4 i1_3_lut_3_lut (.A(n27112), .B(n27391), .C(n8274), .Z(n23498)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_3_lut_3_lut.init = 16'h0404;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n27112), .B(n23594), .C(n27114), .D(n27108), 
         .Z(n23598)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 i23464_2_lut_3_lut_4_lut (.A(n14470), .B(n27110), .C(rst_reg_n), 
         .D(n27342), .Z(clk_c_enable_68)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A ((D)+!C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(208[14] 211[12])
    defparam i23464_2_lut_3_lut_4_lut.init = 16'hdf0f;
    LUT4 n26060_bdd_3_lut (.A(n26060), .B(load_top_bit), .C(data_out_3__N_1385), 
         .Z(n26061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26060_bdd_3_lut.init = 16'hcaca;
    LUT4 i12506_4_lut_4_lut (.A(n27348), .B(alu_a_in_3__N_1552), .C(\debug_branch_N_442[29] ), 
         .D(data_rs1[1]), .Z(\alu_a_in[1] )) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i12506_4_lut_4_lut.init = 16'h5140;
    LUT4 debug_branch_N_840_29__bdd_3_lut_24086 (.A(\debug_branch_N_840[29] ), 
         .B(\timer_data[1] ), .C(is_timer_addr), .Z(n26060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam debug_branch_N_840_29__bdd_3_lut_24086.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_256 (.A(alu_op[2]), .B(n27347), .C(n27346), 
         .D(n27369), .Z(clk_c_enable_321)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam i1_3_lut_4_lut_adj_256.init = 16'h0fef;
    LUT4 dr_3__N_1864_32__bdd_3_lut_24097_4_lut (.A(alu_op[2]), .B(n27347), 
         .C(\mul_out[2] ), .D(alu_out[2]), .Z(n26684)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam dr_3__N_1864_32__bdd_3_lut_24097_4_lut.init = 16'hfe10;
    LUT4 mux_72_i4_3_lut_4_lut (.A(alu_op[2]), .B(n27347), .C(alu_out[3]), 
         .D(\mul_out[3] ), .Z(n191[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam mux_72_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_72_i2_3_lut_4_lut (.A(alu_op[2]), .B(n27347), .C(alu_out[1]), 
         .D(\mul_out[1] ), .Z(n191[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(61[19:40])
    defparam mux_72_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12588_4_lut (.A(mip_reg[17]), .B(n27290), .C(\ui_in_sync[1] ), 
         .D(last_interrupt_req[1]), .Z(n948[1])) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(447[18] 459[12])
    defparam i12588_4_lut.init = 16'h88c8;
    LUT4 i1_4_lut_adj_257 (.A(n1167), .B(n5), .C(data_rs1[1]), .D(n27276), 
         .Z(n822[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_4_lut_adj_257.init = 16'ha088;
    PFUMX i24392 (.BLUT(n27489), .ALUT(n27488), .C0(counter_hi[4]), .Z(n27490));
    LUT4 i12254_4_lut (.A(mip_reg[16]), .B(n27290), .C(\next_fsm_state_3__N_2499[3] ), 
         .D(last_interrupt_req[0]), .Z(n948[0])) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(447[18] 459[12])
    defparam i12254_4_lut.init = 16'h88c8;
    LUT4 i12249_4_lut (.A(n809[0]), .B(n1167), .C(data_rs1[0]), .D(n27276), 
         .Z(n822[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(434[22] 438[16])
    defparam i12249_4_lut.init = 16'hc088;
    LUT4 is_csr_write_bdd_4_lut (.A(\mie[1] ), .B(data_rs1[1]), .C(n27249), 
         .D(n27248), .Z(n26327)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B (D))) */ ;
    defparam is_csr_write_bdd_4_lut.init = 16'hee2a;
    LUT4 counter_hi_4__bdd_4_lut_24187 (.A(counter_hi[4]), .B(mie[11]), 
         .C(mie[3]), .D(counter_hi[3]), .Z(n26343)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (B)) */ ;
    defparam counter_hi_4__bdd_4_lut_24187.init = 16'hcce4;
    PFUMX i24098 (.BLUT(n26686), .ALUT(n26684), .C0(n27302), .Z(n26687));
    LUT4 n26341_bdd_3_lut_24284 (.A(n26341), .B(mie[15]), .C(counter_hi[3]), 
         .Z(n26342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26341_bdd_3_lut_24284.init = 16'hcaca;
    LUT4 counter_hi_4__bdd_3_lut_24186 (.A(counter_hi[4]), .B(mie[7]), .C(mie[16]), 
         .Z(n26341)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam counter_hi_4__bdd_3_lut_24186.init = 16'hd8d8;
    LUT4 n27473_bdd_3_lut (.A(n27473), .B(n27475), .C(n25069), .Z(n28360)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n27473_bdd_3_lut.init = 16'hacac;
    LUT4 n192_bdd_4_lut (.A(n191[3]), .B(n26049), .C(n15), .D(n27302), 
         .Z(n28358)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(((D)+!C)+!B)) */ ;
    defparam n192_bdd_4_lut.init = 16'ha0c0;
    LUT4 i1_3_lut_4_lut_adj_258 (.A(instr_complete_N_1647), .B(clk_c_enable_276), 
         .C(cycle[1]), .D(cycle[0]), .Z(n20944)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_4_lut_adj_258.init = 16'h0770;
    LUT4 mie_4__bdd_4_lut (.A(mie[8]), .B(counter_hi[3]), .C(mie[0]), 
         .D(counter_hi[4]), .Z(n26360)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B+!(C (D)))) */ ;
    defparam mie_4__bdd_4_lut.init = 16'hb8aa;
    LUT4 n26062_bdd_3_lut (.A(n26062), .B(n26059), .C(debug_rd_3__N_1400), 
         .Z(debug_rd[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26062_bdd_3_lut.init = 16'hcaca;
    FD1P3AX shift_amt__i2 (.D(n92[1]), .SP(clk_c_enable_289), .CK(clk_c), 
            .Q(\shift_amt[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i2.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(stall_core), .B(instr_complete_N_1647), .C(n27263), 
         .D(is_load), .Z(n856)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_4_lut.init = 16'h40ff;
    FD1P3AX shift_amt__i3 (.D(n92[2]), .SP(clk_c_enable_289), .CK(clk_c), 
            .Q(shift_amt[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i3.GSR = "DISABLED";
    FD1P3AX shift_amt__i4 (.D(n92[3]), .SP(clk_c_enable_289), .CK(clk_c), 
            .Q(shift_amt[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i4.GSR = "DISABLED";
    FD1P3AX shift_amt__i5 (.D(n92[0]), .SP(clk_c_enable_290), .CK(clk_c), 
            .Q(shift_amt[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i5.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut_adj_259 (.A(stall_core), .B(instr_complete_N_1647), 
         .C(n27263), .D(n22226), .Z(clk_c_enable_423)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_4_lut_adj_259.init = 16'hff40;
    LUT4 interrupt_core_I_32_2_lut_rep_483_4_lut (.A(stall_core), .B(instr_complete_N_1647), 
         .C(n27263), .D(n22898), .Z(n27108)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam interrupt_core_I_32_2_lut_rep_483_4_lut.init = 16'h40ff;
    LUT4 i2_rep_487 (.A(any_additional_mem_ops), .B(clk_c_enable_276), .C(instr_complete_N_1647), 
         .D(n23326), .Z(n27112)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i2_rep_487.init = 16'h4000;
    LUT4 mie_4__bdd_4_lut_23910 (.A(mie[4]), .B(counter_hi[3]), .C(mie[12]), 
         .D(counter_hi[4]), .Z(n26359)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (C))) */ ;
    defparam mie_4__bdd_4_lut_23910.init = 16'he2c0;
    LUT4 i1_2_lut_rep_484_4_lut (.A(stall_core), .B(instr_complete_N_1647), 
         .C(clk_c_enable_276), .D(any_additional_mem_ops), .Z(n27109)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_rep_484_4_lut.init = 16'h4000;
    FD1P3AX tmp_data_i0_i1 (.D(tmp_data_c[5]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i1.GSR = "DISABLED";
    LUT4 i2_1_lut_rep_479_2_lut_4_lut (.A(stall_core), .B(instr_complete_N_1647), 
         .C(clk_c_enable_276), .D(any_additional_mem_ops), .Z(clk_c_enable_275)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i2_1_lut_rep_479_2_lut_4_lut.init = 16'hbfff;
    FD1P3IX mepc_i0_i22 (.D(n658[2]), .SP(clk_c_enable_424), .CD(n9675), 
            .CK(clk_c), .Q(mepc[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i22.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i2 (.D(tmp_data_c[6]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i2.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i3 (.D(tmp_data_c[7]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i3.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i4 (.D(tmp_data_c[8]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i4.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i5 (.D(tmp_data_c[9]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i5.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i6 (.D(tmp_data_c[10]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i6.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i7 (.D(tmp_data_c[11]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i7.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i8 (.D(tmp_data_c[12]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i8.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i9 (.D(tmp_data_c[13]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i9.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i10 (.D(tmp_data_c[14]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i10.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i11 (.D(tmp_data_c[15]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i11.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i12 (.D(tmp_data_c[16]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i12.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i13 (.D(tmp_data_c[17]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i13.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i14 (.D(tmp_data_c[18]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i14.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i15 (.D(tmp_data_c[19]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i15.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i16 (.D(tmp_data_c[20]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i16.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i17 (.D(tmp_data_c[21]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i17.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i18 (.D(tmp_data_c[22]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i18.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i19 (.D(tmp_data_c[23]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i19.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i20 (.D(tmp_data_c[24]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i20.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i21 (.D(tmp_data_c[25]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i21.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i22 (.D(tmp_data_c[26]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i22.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i23 (.D(tmp_data_c[27]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i23.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i24 (.D(tmp_data[28]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i24.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i25 (.D(tmp_data[29]), .SP(clk_c_enable_321), .CK(clk_c), 
            .Q(tmp_data_c[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i25.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i26 (.D(\tmp_data[30] ), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i26.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i27 (.D(\tmp_data[31] ), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(tmp_data_c[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i27.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i30 (.D(tmp_data_in[2]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(\tmp_data[30] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i30.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i31 (.D(tmp_data_in[3]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(\tmp_data[31] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i31.GSR = "DISABLED";
    FD1P3AX mepc_i0_i1 (.D(mepc[5]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i1.GSR = "DISABLED";
    FD1P3AX mepc_i0_i2 (.D(mepc[6]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i2.GSR = "DISABLED";
    FD1P3AX mepc_i0_i3 (.D(mepc[7]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i3.GSR = "DISABLED";
    FD1P3AX mepc_i0_i4 (.D(mepc[8]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i4.GSR = "DISABLED";
    FD1P3AX mepc_i0_i5 (.D(mepc[9]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i5.GSR = "DISABLED";
    FD1P3AX mepc_i0_i6 (.D(mepc[10]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i6.GSR = "DISABLED";
    FD1P3AX mepc_i0_i7 (.D(mepc[11]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i7.GSR = "DISABLED";
    FD1P3AX mepc_i0_i8 (.D(mepc[12]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i8.GSR = "DISABLED";
    FD1P3AX mepc_i0_i9 (.D(mepc[13]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i9.GSR = "DISABLED";
    FD1P3AX mepc_i0_i10 (.D(mepc[14]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i10.GSR = "DISABLED";
    FD1P3AX mepc_i0_i11 (.D(mepc[15]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i11.GSR = "DISABLED";
    FD1P3AX mepc_i0_i12 (.D(mepc[16]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i12.GSR = "DISABLED";
    FD1P3AX mepc_i0_i13 (.D(mepc[17]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i13.GSR = "DISABLED";
    FD1P3AX mepc_i0_i14 (.D(mepc[18]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i14.GSR = "DISABLED";
    FD1P3AX mepc_i0_i15 (.D(mepc[19]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i15.GSR = "DISABLED";
    FD1P3AX mepc_i0_i16 (.D(mepc[20]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i16.GSR = "DISABLED";
    FD1P3AX mepc_i0_i17 (.D(mepc[21]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i17.GSR = "DISABLED";
    FD1P3AX mepc_i0_i18 (.D(mepc[22]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i18.GSR = "DISABLED";
    FD1P3AX mepc_i0_i19 (.D(mepc[23]), .SP(clk_c_enable_424), .CK(clk_c), 
            .Q(mepc[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i19.GSR = "DISABLED";
    LUT4 mux_73_i1_4_lut (.A(cmp), .B(tmp_data_c[0]), .C(n27348), .D(n27346), 
         .Z(n196[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(170[18] 174[35])
    defparam mux_73_i1_4_lut.init = 16'hca0a;
    LUT4 mux_72_i1_4_lut (.A(accum[0]), .B(alu_out[0]), .C(n27292), .D(d_3__N_1868[0]), 
         .Z(n191[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(174[17:35])
    defparam mux_72_i1_4_lut.init = 16'hc5ca;
    LUT4 i23254_3_lut_4_lut (.A(n27369), .B(n27346), .C(n191[1]), .D(\shift_out[1] ), 
         .Z(n196[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam i23254_3_lut_4_lut.init = 16'hf870;
    FD1P3AX last_interrupt_req_i0_i1 (.D(\ui_in_sync[1] ), .SP(clk_c_enable_345), 
            .CK(clk_c), .Q(last_interrupt_req[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam last_interrupt_req_i0_i1.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_260 (.A(n27368), .B(n27366), .C(\imm[7] ), 
         .D(n46), .Z(n7717)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(75[19:52])
    defparam i1_3_lut_4_lut_adj_260.init = 16'h0800;
    LUT4 mux_87_i1_3_lut (.A(n26733), .B(\debug_branch_N_450[0] ), .C(n25053), 
         .Z(debug_rd_3__N_1571[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam mux_87_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_261 (.A(debug_instr_valid), .B(debug_rd_3__N_1575), 
         .C(n27367), .D(n7590), .Z(debug_reg_wen_N_1689)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(184[18] 194[12])
    defparam i1_4_lut_adj_261.init = 16'hfefc;
    LUT4 n26343_bdd_4_lut_24570 (.A(n26343), .B(n26342), .C(counter_hi[2]), 
         .D(n4521), .Z(csr_read_3__N_1447[3])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n26343_bdd_4_lut_24570.init = 16'hca00;
    LUT4 i1_4_lut_adj_262 (.A(n24410), .B(n27346), .C(n27376), .D(alu_op[1]), 
         .Z(n15)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_4_lut_adj_262.init = 16'hfbff;
    LUT4 i1_3_lut_adj_263 (.A(counter_hi[2]), .B(alu_op[2]), .C(alu_op[3]), 
         .Z(n24410)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_3_lut_adj_263.init = 16'hfefe;
    LUT4 tmp_data_in_3__I_124_i3_4_lut (.A(data_rs1[2]), .B(mstatus_mte), 
         .C(n27242), .D(n27256), .Z(tmp_data_in_3__N_1514[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_124_i3_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_rep_653_4_lut (.A(alu_op[2]), .B(n27366), .C(n27368), 
         .D(n27374), .Z(n27278)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_653_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_654_4_lut (.A(alu_op[2]), .B(n27366), .C(n27368), 
         .D(n27332), .Z(n27279)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_654_4_lut.init = 16'h0010;
    LUT4 i12569_2_lut (.A(n26687), .B(n15), .Z(debug_rd_3__N_1559[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[18] 174[35])
    defparam i12569_2_lut.init = 16'h8888;
    LUT4 imm_3__I_0_i1_3_lut (.A(\debug_rd_3__N_405[28] ), .B(data_rs2[0]), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 i4698_3_lut (.A(debug_instr_valid), .B(is_auipc), .C(is_jal), 
         .Z(alu_a_in_3__N_1552)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(108[27:47])
    defparam i4698_3_lut.init = 16'ha8a8;
    LUT4 imm_3__I_0_i3_3_lut (.A(\debug_rd_3__N_405[30] ), .B(data_rs2[2]), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 imm_3__I_0_i2_3_lut (.A(\debug_rd_3__N_405[29] ), .B(data_rs2[1]), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 n26360_bdd_4_lut (.A(n26360), .B(n26359), .C(counter_hi[2]), 
         .D(n4521), .Z(csr_read_3__N_1447[0])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n26360_bdd_4_lut.init = 16'hca00;
    LUT4 i1_3_lut_adj_264 (.A(\tmp_data[30] ), .B(\tmp_data[31] ), .C(cycle[0]), 
         .Z(instr_complete_N_1656)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_adj_264.init = 16'hf7f7;
    LUT4 cycle_0__I_0_548_3_lut (.A(cycle[0]), .B(cmp_out), .C(alu_op[0]), 
         .Z(instr_complete_N_1654)) /* synthesis lut_function=(A+!(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(224[34:67])
    defparam cycle_0__I_0_548_3_lut.init = 16'hbebe;
    LUT4 mux_3207_i1_3_lut (.A(n26979), .B(n24801), .C(n5160), .Z(n5171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3207_i1_3_lut.init = 16'hcaca;
    FD1P3IX mip_reg__i17 (.D(n979[1]), .SP(clk_c_enable_350), .CD(n27218), 
            .CK(clk_c), .Q(mip_reg[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mip_reg__i17.GSR = "DISABLED";
    LUT4 i10349_3_lut (.A(tmp_data[29]), .B(tmp_data_c[2]), .C(alu_op[2]), 
         .Z(a_for_shift_right[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    defparam i10349_3_lut.init = 16'hcaca;
    LUT4 mux_351_i2_3_lut_4_lut (.A(clk_c_enable_276), .B(n22499), .C(n4575[1]), 
         .D(n1766), .Z(\instr_write_offset_3__N_934[1] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_351_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_351_i1_3_lut_4_lut (.A(clk_c_enable_276), .B(n22499), .C(n4575[0]), 
         .D(n1767), .Z(\instr_write_offset_3__N_934[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_351_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 interrupt_core_I_31_2_lut_rep_481_3_lut_4_lut (.A(clk_c_enable_276), 
         .B(n22499), .C(n27111), .D(n22898), .Z(n27106)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (C+!(D))) */ ;
    defparam interrupt_core_I_31_2_lut_rep_481_3_lut_4_lut.init = 16'hf8ff;
    LUT4 i1_4_lut_adj_265 (.A(n27279), .B(instr_complete_N_1648), .C(n27288), 
         .D(n23264), .Z(instr_complete_N_1647)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i1_4_lut_adj_265.init = 16'hfffe;
    LUT4 mux_352_i2_3_lut_4_lut (.A(clk_c_enable_276), .B(n22499), .C(n4575[1]), 
         .D(n1768[1]), .Z(pc_2__N_932[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_352_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_352_i1_3_lut_4_lut (.A(clk_c_enable_276), .B(n22499), .C(n4575[0]), 
         .D(n1768[0]), .Z(pc_2__N_932[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_352_i1_3_lut_4_lut.init = 16'hf780;
    FD1P3IX mcause__i1 (.D(n616), .SP(clk_c_enable_367), .CD(n27326), 
            .CK(clk_c), .Q(\mcause[1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i1.GSR = "DISABLED";
    FD1P3IX mcause__i2 (.D(n27308), .SP(clk_c_enable_367), .CD(n27326), 
            .CK(clk_c), .Q(\mcause[2] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i2.GSR = "DISABLED";
    FD1P3IX mcause__i3 (.D(n23213), .SP(clk_c_enable_367), .CD(n27326), 
            .CK(clk_c), .Q(mcause[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i3.GSR = "DISABLED";
    FD1P3IX mcause__i4 (.D(n611[4]), .SP(clk_c_enable_367), .CD(n27326), 
            .CK(clk_c), .Q(mcause[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i4.GSR = "DISABLED";
    FD1P3IX mcause__i5 (.D(interrupt_core), .SP(clk_c_enable_367), .CD(n27326), 
            .CK(clk_c), .Q(\mcause[5] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i5.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_266 (.A(debug_instr_valid), .B(interrupt_core), .C(n24018), 
         .D(n24014), .Z(n23264)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i1_4_lut_adj_266.init = 16'heeec;
    LUT4 i1_4_lut_adj_267 (.A(is_branch), .B(is_jalr), .C(is_auipc), .D(is_system), 
         .Z(n24018)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(218[17:110])
    defparam i1_4_lut_adj_267.init = 16'hfffe;
    LUT4 i5872_3_lut_4_lut (.A(is_alu_imm), .B(is_alu_reg), .C(is_auipc), 
         .D(debug_instr_valid), .Z(debug_rd_3__N_1400)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(225[22:46])
    defparam i5872_3_lut_4_lut.init = 16'hfe00;
    FD1P3AX mstatus_mie_524 (.D(mstatus_mie_N_1707), .SP(clk_c_enable_421), 
            .CK(clk_c), .Q(mstatus_mie)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam mstatus_mie_524.GSR = "DISABLED";
    FD1P3IX load_top_bit_513 (.D(\debug_branch_N_450[3] ), .SP(clk_c_enable_422), 
            .CD(n15206), .CK(clk_c), .Q(load_top_bit)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(156[12] 157[43])
    defparam load_top_bit_513.GSR = "DISABLED";
    FD1P3IX mepc_i0_i23 (.D(n658[3]), .SP(clk_c_enable_424), .CD(n9675), 
            .CK(clk_c), .Q(mepc[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i23.GSR = "DISABLED";
    LUT4 i4714_2_lut_3_lut (.A(is_alu_imm), .B(is_alu_reg), .C(debug_instr_valid), 
         .Z(debug_rd_3__N_1401)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(225[22:46])
    defparam i4714_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut (.A(is_lui), .B(is_jal), .Z(n24014)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(218[17:110])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 mie_0__bdd_4_lut (.A(mie[0]), .B(data_rs1[0]), .C(n27249), .D(n27248), 
         .Z(n26532)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B (D))) */ ;
    defparam mie_0__bdd_4_lut.init = 16'hee2a;
    LUT4 i1_4_lut_adj_268 (.A(n23318), .B(cmp_out), .C(n27350), .D(mem_op[0]), 
         .Z(n22499)) /* synthesis lut_function=(A+!(B ((D)+!C)+!B !(C (D)))) */ ;
    defparam i1_4_lut_adj_268.init = 16'hbaea;
    LUT4 i12508_4_lut_4_lut (.A(n27348), .B(alu_a_in_3__N_1552), .C(\debug_branch_N_442[31] ), 
         .D(data_rs1[3]), .Z(alu_a_in[3])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i12508_4_lut_4_lut.init = 16'h5140;
    LUT4 i1_4_lut_adj_269 (.A(n27279), .B(n27278), .C(n27293), .D(interrupt_core), 
         .Z(n23318)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_269.init = 16'hfffe;
    LUT4 i1_2_lut_rep_697 (.A(cycle[0]), .B(cycle[1]), .Z(n27322)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam i1_2_lut_rep_697.init = 16'heeee;
    LUT4 i23549_2_lut_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(counter_hi[2]), 
         .D(n27376), .Z(clk_c_enable_289)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam i23549_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i23563_2_lut_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(n27376), 
         .D(counter_hi[2]), .Z(clk_c_enable_290)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam i23563_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i4475_2_lut (.A(time_hi[0]), .B(clk_c_enable_73), .Z(n1[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam i4475_2_lut.init = 16'h6666;
    LUT4 imm_3__I_0_i4_3_lut (.A(\debug_rd_3__N_405[31] ), .B(data_rs2[3]), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 i4699_3_lut (.A(debug_instr_valid), .B(is_alu_reg), .C(is_branch), 
         .Z(alu_b_in_3__N_1504)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:52])
    defparam i4699_3_lut.init = 16'ha8a8;
    LUT4 i1_3_lut_adj_270 (.A(interrupt_pending_N_1671), .B(no_write_in_progress), 
         .C(mstatus_mie), .Z(n23326)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_adj_270.init = 16'h8080;
    LUT4 mux_3207_i4_3_lut (.A(n24789), .B(n5155[3]), .C(n5160), .Z(n5168)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3207_i4_3_lut.init = 16'hcaca;
    LUT4 mux_3203_i4_4_lut (.A(n5123[3]), .B(mepc[3]), .C(\imm[0] ), .D(n22121), 
         .Z(n5155[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3203_i4_4_lut.init = 16'hca0a;
    LUT4 tmp_data_in_3__I_124_i2_3_lut (.A(tmp_data_in_3__N_1582[1]), .B(data_rs1[1]), 
         .C(n5215), .Z(tmp_data_in_3__N_1514[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_124_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_704 (.A(\imm[3] ), .B(\imm[5] ), .Z(n27329)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i1_2_lut_rep_704.init = 16'heeee;
    LUT4 i9805_4_lut (.A(alu_op[0]), .B(alu_op[2]), .C(alu_op[1]), .D(alu_op[3]), 
         .Z(n5215)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    defparam i9805_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_rep_662_3_lut (.A(\imm[3] ), .B(\imm[5] ), .C(\imm[4] ), 
         .Z(n27287)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i1_2_lut_rep_662_3_lut.init = 16'hfefe;
    LUT4 i23581_2_lut_3_lut (.A(\imm[3] ), .B(\imm[5] ), .C(\imm[2] ), 
         .Z(n22178)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i23581_2_lut_3_lut.init = 16'h0101;
    LUT4 and_454_i1_2_lut (.A(mip_reg[16]), .B(mie[0]), .Z(interrupt_pending_N_1672[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[48:59])
    defparam and_454_i1_2_lut.init = 16'h8888;
    LUT4 mux_327_i1_4_lut (.A(n27249), .B(data_rs1[0]), .C(n27248), .D(mip_reg[16]), 
         .Z(n809[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(437[22:76])
    defparam mux_327_i1_4_lut.init = 16'hf2c0;
    LUT4 i11310_4_lut (.A(data_rs1[1]), .B(n27248), .C(n27249), .D(mip_reg[17]), 
         .Z(n5)) /* synthesis lut_function=(A (B)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(78[10:20])
    defparam i11310_4_lut.init = 16'hdc88;
    FD1S3AX cycle__i0 (.D(n26802), .CK(clk_c), .Q(cycle[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam cycle__i0.GSR = "DISABLED";
    LUT4 i12714_2_lut_rep_707 (.A(\imm[8] ), .B(\imm[9] ), .Z(n27332)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12714_2_lut_rep_707.init = 16'heeee;
    LUT4 i12507_4_lut_4_lut (.A(n27348), .B(alu_a_in_3__N_1552), .C(\debug_branch_N_442[30] ), 
         .D(data_rs1[2]), .Z(alu_a_in[2])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i12507_4_lut_4_lut.init = 16'h5140;
    LUT4 i12241_2_lut_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), .C(n8786), 
         .D(n27305), .Z(n4674[0])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i12241_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 is_trap_I_0_586_2_lut_rep_617_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), 
         .C(interrupt_core), .D(n27305), .Z(n27242)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam is_trap_I_0_586_2_lut_rep_617_3_lut_4_lut.init = 16'hf1f0;
    PFUMX i23998 (.BLUT(n26532), .ALUT(n28580), .C0(n27276), .Z(n26533));
    LUT4 i1_4_lut_4_lut_adj_271 (.A(\imm[6] ), .B(\imm[10] ), .C(n26318), 
         .D(n22178), .Z(n23101)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam i1_4_lut_4_lut_adj_271.init = 16'h4000;
    LUT4 i4299_1_lut_rep_713 (.A(counter_hi[2]), .Z(n27338)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i4299_1_lut_rep_713.init = 16'h5555;
    LUT4 i1_3_lut_4_lut_adj_272 (.A(n28573), .B(counter_hi[2]), .C(debug_instr_valid), 
         .D(n28571), .Z(n22898)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_272.init = 16'hf7ff;
    LUT4 i17744_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(counter_hi[4]), 
         .Z(n18)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i17744_2_lut_3_lut.init = 16'h7878;
    L6MUX21 i24394 (.D0(n234[2]), .D1(n27490), .SD(n25069), .Z(n27491));
    LUT4 i1_3_lut_4_lut_adj_273 (.A(mip_reg[17]), .B(\mie[1] ), .C(n27343), 
         .D(interrupt_pending_N_1672[0]), .Z(interrupt_pending_N_1671)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam i1_3_lut_4_lut_adj_273.init = 16'hfff8;
    LUT4 reduce_or_226_i5_3_lut_4_lut (.A(mip_reg[17]), .B(\mie[1] ), .C(n27343), 
         .D(interrupt_pending_N_1672[0]), .Z(n5_adj_2620)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam reduce_or_226_i5_3_lut_4_lut.init = 16'hf0f8;
    LUT4 i1_2_lut_rep_718 (.A(mie[16]), .B(timer_interrupt), .Z(n27343)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam i1_2_lut_rep_718.init = 16'h8888;
    LUT4 i12586_2_lut_3_lut (.A(mie[16]), .B(timer_interrupt), .C(interrupt_core), 
         .Z(n611[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam i12586_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_683_3_lut (.A(mie[16]), .B(timer_interrupt), .C(interrupt_core), 
         .Z(n27308)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam i1_2_lut_rep_683_3_lut.init = 16'h8080;
    LUT4 i23452_2_lut_rep_721 (.A(cycle[1]), .B(cycle[0]), .Z(n27346)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i23452_2_lut_rep_721.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(cycle[1]), .B(cycle[0]), .C(tmp_data_c[1]), 
         .Z(debug_rd_3__N_1563[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_274 (.A(cycle[1]), .B(cycle[0]), .C(tmp_data_c[2]), 
         .Z(debug_rd_3__N_1563[2])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_274.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_275 (.A(cycle[1]), .B(cycle[0]), .C(tmp_data_c[3]), 
         .Z(debug_rd_3__N_1563[3])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_275.init = 16'h4040;
    LUT4 tmp_data_in_3__I_124_i1_3_lut (.A(tmp_data_in_3__N_1582[0]), .B(data_rs1[0]), 
         .C(n5215), .Z(tmp_data_in_3__N_1514[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_124_i1_3_lut.init = 16'hcaca;
    LUT4 is_jal_I_0_2_lut_rep_724 (.A(is_jal), .B(is_jalr), .Z(n27349)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam is_jal_I_0_2_lut_rep_724.init = 16'heeee;
    LUT4 i22799_2_lut_3_lut_4_lut (.A(is_jal), .B(is_jalr), .C(n27362), 
         .D(debug_instr_valid), .Z(n25142)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam i22799_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i4709_2_lut_rep_668_3_lut (.A(is_jal), .B(is_jalr), .C(debug_instr_valid), 
         .Z(n27293)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam i4709_2_lut_rep_668_3_lut.init = 16'he0e0;
    LUT4 i4705_2_lut_3_lut (.A(is_jal), .B(is_jalr), .C(is_lui), .Z(n7590)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam i4705_2_lut_3_lut.init = 16'hfefe;
    LUT4 i23662_2_lut_3_lut_3_lut_4_lut (.A(is_jal), .B(is_jalr), .C(debug_instr_valid), 
         .D(is_lui), .Z(n25072)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam i23662_2_lut_3_lut_3_lut_4_lut.init = 16'hff1f;
    LUT4 i1_3_lut_4_lut_adj_276 (.A(data_rs1[1]), .B(n27231), .C(n20), 
         .D(\mie[13] ), .Z(n21454)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(450[22] 451[75])
    defparam i1_3_lut_4_lut_adj_276.init = 16'h8f88;
    LUT4 mux_251_i2_3_lut (.A(mepc[1]), .B(data_rs1[1]), .C(n652), .Z(n653[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i2_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_277 (.A(data_rs1[1]), .B(n27231), .C(n20), 
         .D(\mie[9] ), .Z(n21452)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(450[22] 451[75])
    defparam i1_3_lut_4_lut_adj_277.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_278 (.A(data_rs1[1]), .B(n27231), .C(n20), 
         .D(\mie[5] ), .Z(n21450)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(450[22] 451[75])
    defparam i1_3_lut_4_lut_adj_278.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_279 (.A(n27231), .B(data_rs1[3]), .C(n14), 
         .D(mie[15]), .Z(n21490)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_279.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_280 (.A(n27231), .B(data_rs1[3]), .C(n14), 
         .D(mie[11]), .Z(n21488)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_280.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_281 (.A(n27231), .B(data_rs1[3]), .C(n14), 
         .D(mie[16]), .Z(n21486)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_281.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_282 (.A(n27231), .B(data_rs1[3]), .C(n14), 
         .D(mie[7]), .Z(n21484)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_282.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_283 (.A(n27231), .B(data_rs1[3]), .C(n14), 
         .D(mie[3]), .Z(n21482)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_283.init = 16'h8f88;
    LUT4 i12169_2_lut (.A(cycle[1]), .B(cycle[0]), .Z(n14470)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12169_2_lut.init = 16'h8888;
    LUT4 mstatus_mie_I_153_3_lut_4_lut (.A(n27231), .B(data_rs1[3]), .C(n27278), 
         .D(mstatus_mpie), .Z(mstatus_mie_N_1709)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam mstatus_mie_I_153_3_lut_4_lut.init = 16'hf808;
    LUT4 n27491_bdd_3_lut_24400 (.A(n27491), .B(debug_rd_3__N_1396[2]), 
         .C(debug_rd_3__N_1400), .Z(debug_rd_3__N_1392[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27491_bdd_3_lut_24400.init = 16'hcaca;
    LUT4 i3889_3_lut (.A(time_hi[2]), .B(time_hi[1]), .C(time_hi[0]), 
         .Z(n498[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(295[55:71])
    defparam i3889_3_lut.init = 16'h6a6a;
    LUT4 i3882_2_lut (.A(time_hi[1]), .B(time_hi[0]), .Z(n498[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(295[55:71])
    defparam i3882_2_lut.init = 16'h6666;
    L6MUX21 instr_complete_I_131 (.D0(instr_complete_N_1650), .D1(instr_complete_N_1649), 
            .SD(n24838), .Z(instr_complete_N_1648)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX instr_complete_I_132 (.BLUT(instr_complete_N_1654), .ALUT(instr_complete_N_1656), 
          .C0(debug_rd_3__N_413), .Z(instr_complete_N_1649)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX tmp_data_in_3__I_0_i4 (.BLUT(tmp_data_in_3__N_1582[3]), .ALUT(\tmp_data_in_3__N_1514[3] ), 
          .C0(n25081), .Z(tmp_data_in[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX debug_rd_3__I_121_i3 (.BLUT(debug_rd_3__N_1563[2]), .ALUT(debug_rd_3__N_1559[2]), 
          .C0(n27274), .Z(debug_rd_3__N_1396[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX tmp_data_in_3__I_0_i3 (.BLUT(tmp_data_in_3__N_1582[2]), .ALUT(tmp_data_in_3__N_1514[2]), 
          .C0(n25081), .Z(tmp_data_in[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_adj_284 (.A(alu_op[3]), .B(alu_op[2]), .C(alu_op[1]), 
         .Z(n22788)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_adj_284.init = 16'h1010;
    PFUMX debug_rd_3__I_122_i1 (.BLUT(\debug_rd_3__N_1567[0] ), .ALUT(debug_rd_3__N_1571[0]), 
          .C0(debug_rd_3__N_1575), .Z(debug_rd_3__N_1392[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX debug_reg_wen_I_0 (.BLUT(debug_reg_wen_N_1689), .ALUT(debug_reg_wen_N_1692), 
          .C0(debug_rd_3__N_1400), .Z(debug_reg_wen)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX debug_rd_3__I_121_i1 (.BLUT(\shift_out[0] ), .ALUT(debug_rd_3__N_1559[0]), 
          .C0(n25132), .Z(debug_rd_3__N_1396[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i23601_2_lut (.A(\imm[1] ), .B(\imm[0] ), .Z(n25119)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i23601_2_lut.init = 16'hbbbb;
    LUT4 c_2__N_1861_1__bdd_4_lut_4_lut (.A(n28573), .B(counter_hi[2]), 
         .C(\pc[21] ), .D(\pc[17] ), .Z(n26200)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam c_2__N_1861_1__bdd_4_lut_4_lut.init = 16'h5140;
    LUT4 i12321_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[20] ), 
         .D(\next_pc_for_core[16] ), .Z(n225)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i12321_4_lut_4_lut.init = 16'h5140;
    LUT4 c_2__N_1861_1__bdd_4_lut_23807_4_lut (.A(n28573), .B(counter_hi[2]), 
         .C(\pc[23] ), .D(\pc[19] ), .Z(n26175)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam c_2__N_1861_1__bdd_4_lut_23807_4_lut.init = 16'h5140;
    LUT4 i12303_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\pc[20] ), 
         .D(\pc[16] ), .Z(n225_adj_4)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i12303_4_lut_4_lut.init = 16'h5140;
    LUT4 i1_3_lut_3_lut_adj_285 (.A(counter_hi[3]), .B(counter_hi[2]), .C(counter_hi[4]), 
         .Z(n4521)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_3_lut_3_lut_adj_285.init = 16'hf4f4;
    LUT4 i12322_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[21] ), 
         .D(\next_pc_for_core[17] ), .Z(n226)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i12322_4_lut_4_lut.init = 16'h5140;
    LUT4 c_2__N_1861_1__bdd_4_lut_23811_4_lut (.A(n28573), .B(counter_hi[2]), 
         .C(\pc[22] ), .D(\pc[18] ), .Z(n26195)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam c_2__N_1861_1__bdd_4_lut_23811_4_lut.init = 16'h5140;
    LUT4 dr_3__N_1864_32__bdd_3_lut_24475 (.A(dr_3__N_1864[32]), .B(dr_3__N_1864[33]), 
         .C(alu_op[2]), .Z(n26685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam dr_3__N_1864_32__bdd_3_lut_24475.init = 16'hcaca;
    LUT4 i12580_2_lut (.A(data_rs2[2]), .B(data_out_3__N_1385), .Z(\data_out_slice[2] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i12580_2_lut.init = 16'h2222;
    LUT4 i23683_4_lut (.A(n27280), .B(n27367), .C(\imm[6] ), .D(\imm[2] ), 
         .Z(n1167)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i23683_4_lut.init = 16'h4000;
    LUT4 i12581_2_lut_rep_589 (.A(data_rs2[3]), .B(data_out_3__N_1385), 
         .Z(n27214)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i12581_2_lut_rep_589.init = 16'h2222;
    LUT4 mtimecmp_7__I_0_3_lut_4_lut (.A(data_rs2[3]), .B(data_out_3__N_1385), 
         .C(n27223), .D(\mtimecmp[7] ), .Z(mtimecmp_3__N_1935)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam mtimecmp_7__I_0_3_lut_4_lut.init = 16'h2f20;
    L6MUX21 i24863 (.D0(n28361), .D1(n28359), .SD(debug_rd_3__N_1400), 
            .Z(debug_rd[3]));
    PFUMX i24861 (.BLUT(n28360), .ALUT(debug_rd_3__N_1571[3]), .C0(debug_rd_3__N_1575), 
          .Z(n28361));
    LUT4 i12248_3_lut_4_lut (.A(rst_reg_n), .B(n27234), .C(n27235), .D(mstatus_mie_N_1709), 
         .Z(mstatus_mie_N_1707)) /* synthesis lut_function=((B+!(C+!(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(395[13:37])
    defparam i12248_3_lut_4_lut.init = 16'hdfdd;
    PFUMX i24859 (.BLUT(debug_rd_3__N_1563[3]), .ALUT(n28358), .C0(n27274), 
          .Z(n28359));
    LUT4 i1_3_lut_4_lut_adj_286 (.A(rst_reg_n), .B(n27234), .C(n27309), 
         .D(n27290), .Z(clk_c_enable_345)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(395[13:37])
    defparam i1_3_lut_4_lut_adj_286.init = 16'h2000;
    PFUMX mux_91_i2 (.BLUT(n24772), .ALUT(\debug_branch_N_446[29] ), .C0(n25072), 
          .Z(n234[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX i23740 (.BLUT(debug_rd_3__N_1567[1]), .ALUT(n26061), .C0(debug_rd_3__N_1575), 
          .Z(n26062));
    LUT4 i12579_2_lut_rep_597 (.A(data_rs2[1]), .B(data_out_3__N_1385), 
         .Z(n27222)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i12579_2_lut_rep_597.init = 16'h2222;
    LUT4 mtimecmp_5__I_0_3_lut_4_lut (.A(data_rs2[1]), .B(data_out_3__N_1385), 
         .C(n27223), .D(\mtimecmp[5] ), .Z(mtimecmp_1__N_1941)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam mtimecmp_5__I_0_3_lut_4_lut.init = 16'h2f20;
    LUT4 i6738_4_lut (.A(mem_op[1]), .B(mem_op[0]), .C(counter_hi[4]), 
         .D(counter_hi[3]), .Z(data_out_3__N_1385)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[13] 272[50])
    defparam i6738_4_lut.init = 16'h5150;
    LUT4 i2_2_lut_3_lut_4_lut (.A(\imm[2] ), .B(n27247), .C(n27290), .D(n27309), 
         .Z(clk_c_enable_87)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\imm[2] ), .B(n27247), .C(n27296), .D(n27309), 
         .Z(clk_c_enable_91)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0200;
    PFUMX mux_443_i1 (.BLUT(n822[0]), .ALUT(n948[0]), .C0(n27296), .Z(n979[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    L6MUX21 debug_rd_3__I_0_i1 (.D0(debug_rd_3__N_1392[0]), .D1(debug_rd_3__N_1396[0]), 
            .SD(debug_rd_3__N_1400), .Z(debug_rd[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX i23888 (.BLUT(n26327), .ALUT(n28581), .C0(n27276), .Z(n26328));
    LUT4 mux_251_i3_3_lut (.A(mepc[2]), .B(data_rs1[2]), .C(n652), .Z(n653[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i3_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_287 (.A(n27322), .B(clk_c_enable_276), .C(n8197), 
         .D(n27321), .Z(address_ready)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_287.init = 16'h4000;
    LUT4 rstn_N_1579_I_0_2_lut_rep_593_4_lut (.A(mstatus_mte), .B(is_double_fault_r), 
         .C(n27256), .D(n28575), .Z(n27218)) /* synthesis lut_function=(A (B+!(D))+!A (B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(365[28:90])
    defparam rstn_N_1579_I_0_2_lut_rep_593_4_lut.init = 16'hdcff;
    PFUMX mux_443_i2 (.BLUT(n822[1]), .ALUT(n948[1]), .C0(n27296), .Z(n979[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX mux_91_i3 (.BLUT(n24775), .ALUT(\debug_branch_N_446[30] ), .C0(n25072), 
          .Z(n234[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i12244_2_lut_4_lut (.A(mstatus_mte), .B(is_double_fault_r), .C(n27256), 
         .D(n27235), .Z(mstatus_mte_N_1703)) /* synthesis lut_function=(A (B+!(D))+!A (B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(365[28:90])
    defparam i12244_2_lut_4_lut.init = 16'hdcff;
    LUT4 i1_2_lut_3_lut_4_lut_adj_288 (.A(n27306), .B(n27242), .C(n27234), 
         .D(n27278), .Z(clk_c_enable_101)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(398[22:52])
    defparam i1_2_lut_3_lut_4_lut_adj_288.init = 16'hfff4;
    LUT4 i1_2_lut_3_lut_4_lut_adj_289 (.A(n27306), .B(n27242), .C(n27234), 
         .D(n28575), .Z(n24290)) /* synthesis lut_function=(A (C+!(D))+!A (B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(398[22:52])
    defparam i1_2_lut_3_lut_4_lut_adj_289.init = 16'hf4ff;
    LUT4 n26336_bdd_4_lut (.A(n26336), .B(n26335), .C(counter_hi[2]), 
         .D(n4521), .Z(csr_read_3__N_1447[1])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n26336_bdd_4_lut.init = 16'hca00;
    LUT4 i3740_2_lut_4_lut (.A(tmp_data_c[6]), .B(mepc[2]), .C(n27278), 
         .D(\addr_offset[2] ), .Z(n701)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(267[23:65])
    defparam i3740_2_lut_4_lut.init = 16'h35ca;
    LUT4 is_load_I_0_2_lut (.A(is_load), .B(is_store), .Z(n8197)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(237[58:79])
    defparam is_load_I_0_2_lut.init = 16'heeee;
    LUT4 i22291_2_lut_rep_570_3_lut_4_lut (.A(n27279), .B(interrupt_core), 
         .C(n27278), .D(n27306), .Z(n27195)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i22291_2_lut_rep_570_3_lut_4_lut.init = 16'hf0fe;
    LUT4 mux_252_i2_3_lut_4_lut (.A(n27279), .B(interrupt_core), .C(\debug_branch_N_442[29] ), 
         .D(n653[1]), .Z(n658[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_290 (.A(n24290), .B(n27278), .C(n8), .D(n24607), 
         .Z(clk_c_enable_3)) /* synthesis lut_function=(A+!(B+((D)+!C))) */ ;
    defparam i1_4_lut_adj_290.init = 16'haaba;
    LUT4 mux_252_i4_3_lut_4_lut (.A(n27279), .B(interrupt_core), .C(\debug_branch_N_442[31] ), 
         .D(n653[3]), .Z(n658[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i3_3_lut_4_lut (.A(n27279), .B(interrupt_core), .C(\debug_branch_N_442[30] ), 
         .D(n653[2]), .Z(n658[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i3_3_lut_4_lut.init = 16'hf1e0;
    PFUMX mux_252_i1 (.BLUT(n653[0]), .ALUT(n24611), .C0(n27242), .Z(n658[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 debug_rd_3__I_0_i3_4_lut (.A(debug_rd_3__N_1571[2]), .B(debug_rd_3__N_1392[2]), 
         .C(debug_rd_3__N_1400), .D(debug_rd_3__N_1575), .Z(debug_rd[2])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(176[18] 194[12])
    defparam debug_rd_3__I_0_i3_4_lut.init = 16'hcacc;
    LUT4 mux_87_i3_3_lut (.A(n26717), .B(\debug_branch_N_450[2] ), .C(n25053), 
         .Z(debug_rd_3__N_1571[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam mux_87_i3_3_lut.init = 16'hcaca;
    LUT4 i23669_3_lut (.A(data_out_3__N_1385), .B(is_timer_addr), .C(n28571), 
         .Z(n25053)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam i23669_3_lut.init = 16'hfefe;
    LUT4 mux_93_i2_3_lut (.A(n24774), .B(n234[1]), .C(n25069), .Z(debug_rd_3__N_1567[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(187[18] 194[12])
    defparam mux_93_i2_3_lut.init = 16'hacac;
    LUT4 i1_3_lut_4_lut_adj_291 (.A(\imm[6] ), .B(n27280), .C(\imm[2] ), 
         .D(n27306), .Z(n24242)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_3_lut_4_lut_adj_291.init = 16'hfffe;
    L6MUX21 i22446 (.D0(n24787), .D1(n24788), .SD(\imm[10] ), .Z(n24789));
    LUT4 i1_2_lut_rep_605_3_lut (.A(\imm[6] ), .B(n27280), .C(\imm[2] ), 
         .Z(n27230)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_2_lut_rep_605_3_lut.init = 16'hefef;
    LUT4 i23634_2_lut_3_lut_4_lut (.A(\imm[6] ), .B(n27280), .C(n27309), 
         .D(\imm[2] ), .Z(clk_c_enable_74)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i23634_2_lut_3_lut_4_lut.init = 16'h0100;
    L6MUX21 i22458 (.D0(n24799), .D1(n24800), .SD(\imm[0] ), .Z(n24801));
    PFUMX mux_233_i1 (.BLUT(n4674[0]), .ALUT(n5_adj_2620), .C0(interrupt_core), 
          .Z(n611[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX i22456 (.BLUT(csr_read_3__N_1447[0]), .ALUT(\csr_read_3__N_1459[0] ), 
          .C0(\imm[6] ), .Z(n24799));
    LUT4 mux_87_i4_3_lut_4_lut (.A(data_out_3__N_1385), .B(is_timer_addr), 
         .C(n24616), .D(\debug_branch_N_840[31] ), .Z(debug_rd_3__N_1571[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam mux_87_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12235_2_lut (.A(data_rs2[0]), .B(data_out_3__N_1385), .Z(\data_out_slice[0] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i12235_2_lut.init = 16'h2222;
    LUT4 is_double_fault_I_0_3_lut_rep_609_4_lut (.A(n27306), .B(n27279), 
         .C(is_double_fault_r), .D(mstatus_mte), .Z(n27234)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam is_double_fault_I_0_3_lut_rep_609_4_lut.init = 16'hf0f4;
    PFUMX mux_3187_i4 (.BLUT(csr_read_3__N_1447[3]), .ALUT(\csr_read_3__N_1459[3] ), 
          .C0(\imm[6] ), .Z(n5123[3]));
    PFUMX i24304 (.BLUT(n27022), .ALUT(n27020), .C0(n5160), .Z(n27023));
    PFUMX mux_3187_i2 (.BLUT(csr_read_3__N_1447[1]), .ALUT(\csr_read_3__N_1459[1] ), 
          .C0(\imm[6] ), .Z(n5123[1]));
    LUT4 csr_read_3__N_1463_1__bdd_3_lut_24242 (.A(\cycle_count_wide[1] ), 
         .B(instrret_count[1]), .C(\imm[1] ), .Z(n26928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam csr_read_3__N_1463_1__bdd_3_lut_24242.init = 16'hcaca;
    PFUMX i22444 (.BLUT(\csr_read_3__N_1439[3] ), .ALUT(csr_read_3__N_1455[3]), 
          .C0(\imm[1] ), .Z(n24787));
    LUT4 data_rs1_3__I_0_i1_2_lut (.A(data_rs1[0]), .B(cycle[0]), .Z(mul_out_3__N_1510[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i1_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_rep_486_4_lut (.A(clk_c_enable_276), .B(any_additional_mem_ops), 
         .C(instr_complete_N_1647), .D(stall_core), .Z(n27111)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_rep_486_4_lut.init = 16'h0020;
    LUT4 data_rs1_3__I_0_i2_2_lut (.A(data_rs1[1]), .B(cycle[0]), .Z(mul_out_3__N_1510[1])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i2_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i3_2_lut (.A(data_rs1[2]), .B(cycle[0]), .Z(mul_out_3__N_1510[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i3_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i4_2_lut (.A(data_rs1[3]), .B(cycle[0]), .Z(mul_out_3__N_1510[3])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i4_2_lut.init = 16'h8888;
    PFUMX i66 (.BLUT(n22090), .ALUT(n23101), .C0(\imm[11] ), .Z(n46));
    PFUMX i24282 (.BLUT(n26977), .ALUT(n26976), .C0(\imm[0] ), .Z(n26978));
    LUT4 mux_149_i1_3_lut_4_lut (.A(n27322), .B(n27292), .C(alu_out[0]), 
         .D(data_rs2[0]), .Z(tmp_data_in_3__N_1582[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_149_i2_3_lut_4_lut (.A(n27322), .B(n27292), .C(alu_out[1]), 
         .D(data_rs2[1]), .Z(tmp_data_in_3__N_1582[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_149_i4_3_lut_4_lut (.A(n27322), .B(n27292), .C(alu_out[3]), 
         .D(data_rs2[3]), .Z(tmp_data_in_3__N_1582[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_149_i3_3_lut_4_lut (.A(n27322), .B(n27292), .C(alu_out[2]), 
         .D(data_rs2[2]), .Z(tmp_data_in_3__N_1582[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i3_3_lut_4_lut.init = 16'hfb40;
    PFUMX instr_complete_I_133 (.BLUT(instr_complete_N_1651), .ALUT(instr_complete_N_1652), 
          .C0(debug_rd_3__N_1401), .Z(instr_complete_N_1650)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 n26484_bdd_3_lut_4_lut (.A(n27348), .B(alu_op[0]), .C(n26482), 
         .D(n26484), .Z(cmp_out)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam n26484_bdd_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_2756_i3_3_lut_4_lut (.A(n27348), .B(alu_op[0]), .C(alu_b_in[2]), 
         .D(alu_a_in[2]), .Z(n4528[2])) /* synthesis lut_function=(A (C+(D))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam mux_2756_i3_3_lut_4_lut.init = 16'hfbb0;
    LUT4 mux_2756_i2_3_lut_4_lut (.A(n27348), .B(alu_op[0]), .C(alu_b_in[1]), 
         .D(\alu_a_in[1] ), .Z(n4528[1])) /* synthesis lut_function=(A (C+(D))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam mux_2756_i2_3_lut_4_lut.init = 16'hfbb0;
    LUT4 mux_2756_i1_3_lut_4_lut (.A(n27348), .B(alu_op[0]), .C(alu_b_in[0]), 
         .D(alu_a_in[0]), .Z(n4528[0])) /* synthesis lut_function=(A (C+(D))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam mux_2756_i1_3_lut_4_lut.init = 16'hfbb0;
    LUT4 mux_2756_i4_3_lut_4_lut (.A(n27348), .B(alu_op[0]), .C(alu_b_in[3]), 
         .D(alu_a_in[3]), .Z(n4528[3])) /* synthesis lut_function=(A (C+(D))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(62[21:42])
    defparam mux_2756_i4_3_lut_4_lut.init = 16'hfbb0;
    PFUMX i24358 (.BLUT(n27413), .ALUT(n27414), .C0(counter_hi[2]), .Z(n27415));
    PFUMX i24381 (.BLUT(n27472), .ALUT(n27471), .C0(counter_hi[4]), .Z(n27473));
    PFUMX i24354 (.BLUT(n27407), .ALUT(n27408), .C0(counter_hi[3]), .Z(n27409));
    PFUMX i22445 (.BLUT(\time_count[3] ), .ALUT(n5115), .C0(n25119), .Z(n24788));
    PFUMX i24243 (.BLUT(n26931), .ALUT(n5155[1]), .C0(n5160), .Z(n26932));
    tinyqv_mul multiplier (.accum({accum}), .\next_accum[5] (\next_accum[5] ), 
            .\next_accum[6] (\next_accum[6] ), .clk_c(clk_c), .\next_accum[7] (\next_accum[7] ), 
            .mul_out_3__N_1510({mul_out_3__N_1510}), .\tmp_data[0] (tmp_data_c[0]), 
            .\tmp_data[1] (tmp_data_c[1]), .\tmp_data[2] (tmp_data_c[2]), 
            .\tmp_data[3] (tmp_data_c[3]), .\tmp_data[4] (tmp_data_c[4]), 
            .\tmp_data[5] (tmp_data_c[5]), .\tmp_data[6] (tmp_data_c[6]), 
            .\tmp_data[7] (tmp_data_c[7]), .\tmp_data[8] (tmp_data_c[8]), 
            .\tmp_data[9] (tmp_data_c[9]), .\tmp_data[10] (tmp_data_c[10]), 
            .\tmp_data[11] (tmp_data_c[11]), .\tmp_data[12] (tmp_data_c[12]), 
            .\tmp_data[13] (tmp_data_c[13]), .\tmp_data[14] (tmp_data_c[14]), 
            .\tmp_data[15] (tmp_data_c[15]), .d_3__N_1868({d_3__N_1868}), 
            .GND_net(GND_net), .VCC_net(VCC_net), .\next_accum[8] (\next_accum[8] ), 
            .\next_accum[9] (\next_accum[9] ), .\next_accum[10] (\next_accum[10] ), 
            .\next_accum[11] (\next_accum[11] ), .\next_accum[12] (\next_accum[12] ), 
            .\next_accum[13] (\next_accum[13] ), .\next_accum[14] (\next_accum[14] ), 
            .\next_accum[15] (\next_accum[15] ), .\next_accum[16] (\next_accum[16] ), 
            .\next_accum[17] (\next_accum[17] ), .\next_accum[18] (\next_accum[18] ), 
            .\next_accum[19] (\next_accum[19] ), .\next_accum[4] (\next_accum[4] ), 
            .\cycle[0] (cycle[0]), .data_rs1({data_rs1})) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[31:97])
    tinyqv_shifter i_shift (.a_for_shift_right({Open_35, Open_36, Open_37, 
            Open_38, Open_39, Open_40, Open_41, Open_42, Open_43, 
            Open_44, Open_45, Open_46, Open_47, Open_48, Open_49, 
            Open_50, Open_51, Open_52, Open_53, Open_54, Open_55, 
            Open_56, Open_57, Open_58, Open_59, Open_60, Open_61, 
            Open_62, Open_63, Open_64, a_for_shift_right[1:0]}), .shift_amt({Open_65, 
            Open_66, Open_67, Open_68, Open_69, \shift_amt[0] }), 
            .\shift_amt[2]_adj_1 (shift_amt[2]), .\shift_amt[3]_adj_2 (shift_amt[3]), 
            .\tmp_data[5] (tmp_data_c[5]), .\tmp_data[26] (tmp_data_c[26]), 
            .\alu_op[2] (alu_op[2]), .\tmp_data[4] (tmp_data_c[4]), .\tmp_data[27] (tmp_data_c[27]), 
            .\a_for_shift_right[29] (a_for_shift_right[29]), .\a_for_shift_right[30] (a_for_shift_right[30]), 
            .\a_for_shift_right[31] (\a_for_shift_right[31] ), .n62(n62), 
            .\tmp_data[3] (tmp_data_c[3]), .\tmp_data[28] (tmp_data[28]), 
            .\a_for_shift_right[2] (a_for_shift_right[2]), .\tmp_data[16] (tmp_data_c[16]), 
            .\tmp_data[15] (tmp_data_c[15]), .n27377(n27377), .\shift_amt[1] (\shift_amt[1] ), 
            .n8157(n8157), .\dr_3__N_1864[33] (dr_3__N_1864[33]), .\dr_3__N_1864[32] (dr_3__N_1864[32]), 
            .n8153(n8153), .n7278(n7278), .n25292(n25292), .n63(n63), 
            .\counter_hi[2] (counter_hi[2]), .\tmp_data[25] (tmp_data_c[25]), 
            .\tmp_data[6] (tmp_data_c[6]), .\tmp_data[22] (tmp_data_c[22]), 
            .\tmp_data[9] (tmp_data_c[9]), .\tmp_data[21] (tmp_data_c[21]), 
            .\tmp_data[10] (tmp_data_c[10]), .\tmp_data[24] (tmp_data_c[24]), 
            .\tmp_data[7] (tmp_data_c[7]), .\tmp_data[23] (tmp_data_c[23]), 
            .\tmp_data[8] (tmp_data_c[8]), .n28571(n28571), .\shift_amt[4]_adj_3 (shift_amt[4]), 
            .\shift_amt[5] (\shift_amt[5] ), .\counter_hi[4] (counter_hi[4]), 
            .n28573(n28573), .\tmp_data[19] (tmp_data_c[19]), .\tmp_data[12] (tmp_data_c[12]), 
            .\tmp_data[18] (tmp_data_c[18]), .\tmp_data[13] (tmp_data_c[13]), 
            .\tmp_data[20] (tmp_data_c[20]), .\tmp_data[11] (tmp_data_c[11]), 
            .\tmp_data[14] (tmp_data_c[14]), .\tmp_data[17] (tmp_data_c[17])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(133[20:81])
    tinyqv_registers i_registers (.rs1({rs1}), .rd({rd}), .debug_reg_wen(debug_reg_wen), 
            .rs2({rs2}), .clk_c(clk_c), .return_addr({return_addr}), .debug_rd({debug_rd}), 
            .\reg_access[4][3] (\reg_access[4][3] ), .data_rs1({data_rs1}), 
            .n28571(n28571), .n28573(n28573), .\counter_hi[2] (counter_hi[2]), 
            .data_rs2({data_rs2}), .n28580(n28580), .n27231(n27231), .n24605(n24605), 
            .\mie[12] (mie[12]), .n928(n928), .\reg_access[3][2] (\reg_access[3][2] ), 
            .n28581(n28581), .n27205(n27205), .n27113(n27113), .any_additional_mem_ops(any_additional_mem_ops), 
            .n2356(n2356), .\mie[8] (mie[8]), .n895(n895), .\mie[4] (mie[4]), 
            .n862(n862)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(91[9:103])
    tinyqv_counter_U0 i_instrret (.cy(cy_adj_5), .clk_c(clk_c), .n27326(n27326), 
            .\increment_result_3__N_1925[0] (\increment_result_3__N_1925[0] ), 
            .instrret_count({\instrret_count[3] , instrret_count[2:1], \instrret_count[0] }), 
            .n27229(n27229), .n27246(n27246)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(307[20] 315[6])
    \tinyqv_counter(OUTPUT_WIDTH=7)  i_cycles (.cy(cy_adj_6), .clk_c(clk_c), 
            .n27326(n27326), .\increment_result_3__N_1911[1] (\increment_result_3__N_1911[1] ), 
            .\increment_result_3__N_1911[0] (\increment_result_3__N_1911[0] ), 
            .cycle_count_wide({\cycle_count_wide[6] , \cycle_count_wide[5] , 
            \cycle_count_wide[4] , \cycle_count_wide[3] , cycle_count_wide[2], 
            \cycle_count_wide[1] , \cycle_count_wide[0] }), .n27228(n27228), 
            .n27245(n27245), .n27180(n27180)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(281[40] 290[6])
    tinyqv_alu i_alu (.alu_a_in({alu_a_in[3:2], \alu_a_in[1] , alu_a_in[0]}), 
            .n27187(n27187), .n24124(n24124), .alu_b_in({alu_b_in}), .\alu_op[2] (alu_op[2]), 
            .n27188(n27188), .n27252(n27252), .n27215(n27215), .n27154(n27154), 
            .n27181(n27181), .n23342(n23342), .n26482(n26482), .n27267(n27267), 
            .cy_out(cy_out), .n27266(n27266), .n26484(n26484), .n4528({n4528}), 
            .n27270(n27270), .alu_out({alu_out})) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(115[16:93])
    
endmodule
//
// Verilog Description of module tinyqv_mul
//

module tinyqv_mul (accum, \next_accum[5] , \next_accum[6] , clk_c, \next_accum[7] , 
            mul_out_3__N_1510, \tmp_data[0] , \tmp_data[1] , \tmp_data[2] , 
            \tmp_data[3] , \tmp_data[4] , \tmp_data[5] , \tmp_data[6] , 
            \tmp_data[7] , \tmp_data[8] , \tmp_data[9] , \tmp_data[10] , 
            \tmp_data[11] , \tmp_data[12] , \tmp_data[13] , \tmp_data[14] , 
            \tmp_data[15] , d_3__N_1868, GND_net, VCC_net, \next_accum[8] , 
            \next_accum[9] , \next_accum[10] , \next_accum[11] , \next_accum[12] , 
            \next_accum[13] , \next_accum[14] , \next_accum[15] , \next_accum[16] , 
            \next_accum[17] , \next_accum[18] , \next_accum[19] , \next_accum[4] , 
            \cycle[0] , data_rs1) /* synthesis syn_module_defined=1 */ ;
    output [15:0]accum;
    input \next_accum[5] ;
    input \next_accum[6] ;
    input clk_c;
    input \next_accum[7] ;
    input [3:0]mul_out_3__N_1510;
    input \tmp_data[0] ;
    input \tmp_data[1] ;
    input \tmp_data[2] ;
    input \tmp_data[3] ;
    input \tmp_data[4] ;
    input \tmp_data[5] ;
    input \tmp_data[6] ;
    input \tmp_data[7] ;
    input \tmp_data[8] ;
    input \tmp_data[9] ;
    input \tmp_data[10] ;
    input \tmp_data[11] ;
    input \tmp_data[12] ;
    input \tmp_data[13] ;
    input \tmp_data[14] ;
    input \tmp_data[15] ;
    output [19:0]d_3__N_1868;
    input GND_net;
    input VCC_net;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[4] ;
    input \cycle[0] ;
    input [3:0]data_rs1;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n7;
    wire [15:0]accum_15__N_1888;
    
    wire n24326;
    
    LUT4 accum_15__I_0_i2_3_lut (.A(accum[5]), .B(\next_accum[5] ), .C(n7), 
         .Z(accum_15__N_1888[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i2_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i3_3_lut (.A(accum[6]), .B(\next_accum[6] ), .C(n7), 
         .Z(accum_15__N_1888[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i3_3_lut.init = 16'hacac;
    FD1S3AX accum_i0 (.D(accum_15__N_1888[0]), .CK(clk_c), .Q(accum[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i0.GSR = "DISABLED";
    LUT4 accum_15__I_0_i4_3_lut (.A(accum[7]), .B(\next_accum[7] ), .C(n7), 
         .Z(accum_15__N_1888[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i4_3_lut.init = 16'hacac;
    MULT18X18D a_3__I_0_11_mult_2 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(mul_out_3__N_1510[3]), 
            .A2(mul_out_3__N_1510[2]), .A1(mul_out_3__N_1510[1]), .A0(mul_out_3__N_1510[0]), 
            .B17(GND_net), .B16(GND_net), .B15(\tmp_data[15] ), .B14(\tmp_data[14] ), 
            .B13(\tmp_data[13] ), .B12(\tmp_data[12] ), .B11(\tmp_data[11] ), 
            .B10(\tmp_data[10] ), .B9(\tmp_data[9] ), .B8(\tmp_data[8] ), 
            .B7(\tmp_data[7] ), .B6(\tmp_data[6] ), .B5(\tmp_data[5] ), 
            .B4(\tmp_data[4] ), .B3(\tmp_data[3] ), .B2(\tmp_data[2] ), 
            .B1(\tmp_data[1] ), .B0(\tmp_data[0] ), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .P19(d_3__N_1868[19]), .P18(d_3__N_1868[18]), .P17(d_3__N_1868[17]), 
            .P16(d_3__N_1868[16]), .P15(d_3__N_1868[15]), .P14(d_3__N_1868[14]), 
            .P13(d_3__N_1868[13]), .P12(d_3__N_1868[12]), .P11(d_3__N_1868[11]), 
            .P10(d_3__N_1868[10]), .P9(d_3__N_1868[9]), .P8(d_3__N_1868[8]), 
            .P7(d_3__N_1868[7]), .P6(d_3__N_1868[6]), .P5(d_3__N_1868[5]), 
            .P4(d_3__N_1868[4]), .P3(d_3__N_1868[3]), .P2(d_3__N_1868[2]), 
            .P1(d_3__N_1868[1]), .P0(d_3__N_1868[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[52:83])
    defparam a_3__I_0_11_mult_2.REG_INPUTA_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTA_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTA_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_RST = "RST0";
    defparam a_3__I_0_11_mult_2.CLK0_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK1_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK2_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK3_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.HIGHSPEED_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.GSR = "DISABLED";
    defparam a_3__I_0_11_mult_2.CAS_MATCH_REG = "FALSE";
    defparam a_3__I_0_11_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam a_3__I_0_11_mult_2.MULT_BYPASS = "DISABLED";
    defparam a_3__I_0_11_mult_2.RESETMODE = "SYNC";
    LUT4 accum_15__I_0_i5_3_lut (.A(accum[8]), .B(\next_accum[8] ), .C(n7), 
         .Z(accum_15__N_1888[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i5_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i6_3_lut (.A(accum[9]), .B(\next_accum[9] ), .C(n7), 
         .Z(accum_15__N_1888[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i6_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i7_3_lut (.A(accum[10]), .B(\next_accum[10] ), .C(n7), 
         .Z(accum_15__N_1888[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i7_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i8_3_lut (.A(accum[11]), .B(\next_accum[11] ), .C(n7), 
         .Z(accum_15__N_1888[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i8_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i9_3_lut (.A(accum[12]), .B(\next_accum[12] ), .C(n7), 
         .Z(accum_15__N_1888[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i9_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i10_3_lut (.A(accum[13]), .B(\next_accum[13] ), .C(n7), 
         .Z(accum_15__N_1888[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i10_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i11_3_lut (.A(accum[14]), .B(\next_accum[14] ), .C(n7), 
         .Z(accum_15__N_1888[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i11_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i12_3_lut (.A(accum[15]), .B(\next_accum[15] ), .C(n7), 
         .Z(accum_15__N_1888[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i12_3_lut.init = 16'hacac;
    FD1S3IX accum_i12 (.D(\next_accum[16] ), .CK(clk_c), .CD(n7), .Q(accum[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i12.GSR = "DISABLED";
    FD1S3AX accum_i1 (.D(accum_15__N_1888[1]), .CK(clk_c), .Q(accum[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i1.GSR = "DISABLED";
    FD1S3AX accum_i2 (.D(accum_15__N_1888[2]), .CK(clk_c), .Q(accum[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i2.GSR = "DISABLED";
    FD1S3AX accum_i3 (.D(accum_15__N_1888[3]), .CK(clk_c), .Q(accum[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i3.GSR = "DISABLED";
    FD1S3AX accum_i4 (.D(accum_15__N_1888[4]), .CK(clk_c), .Q(accum[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i4.GSR = "DISABLED";
    FD1S3AX accum_i5 (.D(accum_15__N_1888[5]), .CK(clk_c), .Q(accum[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i5.GSR = "DISABLED";
    FD1S3AX accum_i6 (.D(accum_15__N_1888[6]), .CK(clk_c), .Q(accum[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i6.GSR = "DISABLED";
    FD1S3AX accum_i7 (.D(accum_15__N_1888[7]), .CK(clk_c), .Q(accum[7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i7.GSR = "DISABLED";
    FD1S3AX accum_i8 (.D(accum_15__N_1888[8]), .CK(clk_c), .Q(accum[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i8.GSR = "DISABLED";
    FD1S3AX accum_i9 (.D(accum_15__N_1888[9]), .CK(clk_c), .Q(accum[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i9.GSR = "DISABLED";
    FD1S3AX accum_i10 (.D(accum_15__N_1888[10]), .CK(clk_c), .Q(accum[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i10.GSR = "DISABLED";
    FD1S3AX accum_i11 (.D(accum_15__N_1888[11]), .CK(clk_c), .Q(accum[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i11.GSR = "DISABLED";
    FD1S3IX accum_i13 (.D(\next_accum[17] ), .CK(clk_c), .CD(n7), .Q(accum[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i13.GSR = "DISABLED";
    FD1S3IX accum_i14 (.D(\next_accum[18] ), .CK(clk_c), .CD(n7), .Q(accum[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i14.GSR = "DISABLED";
    FD1S3IX accum_i15 (.D(\next_accum[19] ), .CK(clk_c), .CD(n7), .Q(accum[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i15.GSR = "DISABLED";
    LUT4 accum_15__I_0_i1_3_lut (.A(accum[4]), .B(\next_accum[4] ), .C(n7), 
         .Z(accum_15__N_1888[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i1_3_lut.init = 16'hacac;
    LUT4 i23631_4_lut (.A(\cycle[0] ), .B(n24326), .C(data_rs1[3]), .D(data_rs1[0]), 
         .Z(n7)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:32])
    defparam i23631_4_lut.init = 16'h5557;
    LUT4 i1_2_lut (.A(data_rs1[2]), .B(data_rs1[1]), .Z(n24326)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:32])
    defparam i1_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module tinyqv_shifter
//

module tinyqv_shifter (a_for_shift_right, shift_amt, \shift_amt[2]_adj_1 , 
            \shift_amt[3]_adj_2 , \tmp_data[5] , \tmp_data[26] , \alu_op[2] , 
            \tmp_data[4] , \tmp_data[27] , \a_for_shift_right[29] , \a_for_shift_right[30] , 
            \a_for_shift_right[31] , n62, \tmp_data[3] , \tmp_data[28] , 
            \a_for_shift_right[2] , \tmp_data[16] , \tmp_data[15] , n27377, 
            \shift_amt[1] , n8157, \dr_3__N_1864[33] , \dr_3__N_1864[32] , 
            n8153, n7278, n25292, n63, \counter_hi[2] , \tmp_data[25] , 
            \tmp_data[6] , \tmp_data[22] , \tmp_data[9] , \tmp_data[21] , 
            \tmp_data[10] , \tmp_data[24] , \tmp_data[7] , \tmp_data[23] , 
            \tmp_data[8] , n28571, \shift_amt[4]_adj_3 , \shift_amt[5] , 
            \counter_hi[4] , n28573, \tmp_data[19] , \tmp_data[12] , 
            \tmp_data[18] , \tmp_data[13] , \tmp_data[20] , \tmp_data[11] , 
            \tmp_data[14] , \tmp_data[17] ) /* synthesis syn_module_defined=1 */ ;
    input [31:0]a_for_shift_right;
    input [5:0]shift_amt;
    input \shift_amt[2]_adj_1 ;
    input \shift_amt[3]_adj_2 ;
    input \tmp_data[5] ;
    input \tmp_data[26] ;
    input \alu_op[2] ;
    input \tmp_data[4] ;
    input \tmp_data[27] ;
    input \a_for_shift_right[29] ;
    input \a_for_shift_right[30] ;
    input \a_for_shift_right[31] ;
    output n62;
    input \tmp_data[3] ;
    input \tmp_data[28] ;
    input \a_for_shift_right[2] ;
    input \tmp_data[16] ;
    input \tmp_data[15] ;
    input n27377;
    input \shift_amt[1] ;
    output n8157;
    output \dr_3__N_1864[33] ;
    output \dr_3__N_1864[32] ;
    output n8153;
    output n7278;
    input n25292;
    input n63;
    input \counter_hi[2] ;
    input \tmp_data[25] ;
    input \tmp_data[6] ;
    input \tmp_data[22] ;
    input \tmp_data[9] ;
    input \tmp_data[21] ;
    input \tmp_data[10] ;
    input \tmp_data[24] ;
    input \tmp_data[7] ;
    input \tmp_data[23] ;
    input \tmp_data[8] ;
    input n28571;
    input \shift_amt[4]_adj_3 ;
    output \shift_amt[5] ;
    input \counter_hi[4] ;
    input n28573;
    input \tmp_data[19] ;
    input \tmp_data[12] ;
    input \tmp_data[18] ;
    input \tmp_data[13] ;
    input \tmp_data[20] ;
    input \tmp_data[11] ;
    input \tmp_data[14] ;
    input \tmp_data[17] ;
    
    
    wire n101, n105, n25701, n25300, n32, n27336, n25387;
    wire [5:0]shift_amt_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[16:25])
    
    wire n4;
    wire [31:0]a_for_shift_right_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[17:34])
    
    wire n58, n60, n25263, n25264, n25267, n33, n25265, n25266, 
        n25268, n43, n45, n47, n25278, n25279, n25282, n25280, 
        n25281, n25283, n25285, n25286, n25293, n49, n51, n53, 
        n55, n57, n59, n61, n34, n129, n125;
    wire [65:0]dr_3__N_1864;
    
    wire n25287, n25288, n25700, n25294, n121, n117, n25289, n25290, 
        n25295, n36, n25255, n25256, n113, n109, n25257, n25258, 
        n25259, n25260, n25261, n25262, n25270, n25271, n38, n25291, 
        n25699, n25296, n25272, n25273, n25274, n25275, n25276, 
        n25277, n41, n54, n56, n37, n39, n35, n25301, n52, 
        n48, n50, n44, n46, n40, n42, n25302, n25303, n25297, 
        n25298, n25304, n25305;
    
    PFUMX i22957 (.BLUT(n101), .ALUT(n105), .C0(n25701), .Z(n25300));
    LUT4 top_bit_I_0_i32_3_lut (.A(a_for_shift_right[0]), .B(a_for_shift_right[1]), 
         .C(shift_amt[0]), .Z(n32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i32_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(\shift_amt[2]_adj_1 ), .B(n27336), .C(n25387), 
         .D(\shift_amt[3]_adj_2 ), .Z(shift_amt_c[3])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[28:55])
    defparam i2_3_lut_4_lut.init = 16'hd22d;
    LUT4 i4040_3_lut_4_lut (.A(\shift_amt[2]_adj_1 ), .B(n27336), .C(n25387), 
         .D(\shift_amt[3]_adj_2 ), .Z(n4)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[28:55])
    defparam i4040_3_lut_4_lut.init = 16'h2f02;
    LUT4 top_bit_I_0_i58_3_lut (.A(a_for_shift_right_c[26]), .B(a_for_shift_right_c[27]), 
         .C(shift_amt[0]), .Z(n58)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i58_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i27_3_lut (.A(\tmp_data[5] ), .B(\tmp_data[26] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i28_3_lut (.A(\tmp_data[4] ), .B(\tmp_data[27] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i60_3_lut (.A(a_for_shift_right_c[28]), .B(\a_for_shift_right[29] ), 
         .C(shift_amt[0]), .Z(n60)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i60_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i62_3_lut (.A(\a_for_shift_right[30] ), .B(\a_for_shift_right[31] ), 
         .C(shift_amt[0]), .Z(n62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i62_3_lut.init = 16'hcaca;
    L6MUX21 i22924 (.D0(n25263), .D1(n25264), .SD(shift_amt_c[3]), .Z(n25267));
    LUT4 a_0__I_0_i29_3_lut (.A(\tmp_data[3] ), .B(\tmp_data[28] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i33_3_lut (.A(a_for_shift_right[1]), .B(\a_for_shift_right[2] ), 
         .C(shift_amt[0]), .Z(n33)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i33_3_lut.init = 16'hcaca;
    L6MUX21 i22925 (.D0(n25265), .D1(n25266), .SD(shift_amt_c[3]), .Z(n25268));
    LUT4 top_bit_I_0_i43_3_lut (.A(a_for_shift_right_c[11]), .B(a_for_shift_right_c[12]), 
         .C(shift_amt[0]), .Z(n43)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i43_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i45_3_lut (.A(a_for_shift_right_c[13]), .B(a_for_shift_right_c[14]), 
         .C(shift_amt[0]), .Z(n45)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i45_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i47_4_lut (.A(\tmp_data[16] ), .B(\tmp_data[15] ), 
         .C(\alu_op[2] ), .D(shift_amt[0]), .Z(n47)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A !((C (D)+!C !(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i47_4_lut.init = 16'hacca;
    L6MUX21 i22939 (.D0(n25278), .D1(n25279), .SD(shift_amt_c[3]), .Z(n25282));
    L6MUX21 i22940 (.D0(n25280), .D1(n25281), .SD(shift_amt_c[3]), .Z(n25283));
    PFUMX i22950 (.BLUT(n25285), .ALUT(n25286), .C0(n25701), .Z(n25293));
    LUT4 top_bit_I_0_i49_3_lut (.A(a_for_shift_right_c[17]), .B(a_for_shift_right_c[18]), 
         .C(shift_amt[0]), .Z(n49)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i49_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i51_3_lut (.A(a_for_shift_right_c[19]), .B(a_for_shift_right_c[20]), 
         .C(shift_amt[0]), .Z(n51)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i51_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i53_3_lut (.A(a_for_shift_right_c[21]), .B(a_for_shift_right_c[22]), 
         .C(shift_amt[0]), .Z(n53)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i53_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i55_3_lut (.A(a_for_shift_right_c[23]), .B(a_for_shift_right_c[24]), 
         .C(shift_amt[0]), .Z(n55)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i55_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i57_3_lut (.A(a_for_shift_right_c[25]), .B(a_for_shift_right_c[26]), 
         .C(shift_amt[0]), .Z(n57)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i57_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i59_3_lut (.A(a_for_shift_right_c[27]), .B(a_for_shift_right_c[28]), 
         .C(shift_amt[0]), .Z(n59)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i59_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i61_3_lut (.A(\a_for_shift_right[29] ), .B(\a_for_shift_right[30] ), 
         .C(shift_amt[0]), .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i61_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i34_3_lut (.A(\a_for_shift_right[2] ), .B(a_for_shift_right_c[3]), 
         .C(shift_amt[0]), .Z(n34)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i34_3_lut.init = 16'hcaca;
    LUT4 i5108_4_lut (.A(\a_for_shift_right[31] ), .B(n27377), .C(shift_amt[0]), 
         .D(\shift_amt[1] ), .Z(n129)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam i5108_4_lut.init = 16'hccca;
    LUT4 top_bit_I_0_i125_3_lut (.A(n59), .B(n61), .C(\shift_amt[1] ), 
         .Z(n125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i125_3_lut.init = 16'hcaca;
    LUT4 i5839_3_lut (.A(dr_3__N_1864[31]), .B(dr_3__N_1864[34]), .C(\alu_op[2] ), 
         .Z(n8157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i5839_3_lut.init = 16'hcaca;
    PFUMX i22951 (.BLUT(n25287), .ALUT(n25288), .C0(n25700), .Z(n25294));
    LUT4 i5835_3_lut (.A(\dr_3__N_1864[33] ), .B(\dr_3__N_1864[32] ), .C(\alu_op[2] ), 
         .Z(n8153)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i5835_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i121_3_lut (.A(n55), .B(n57), .C(\shift_amt[1] ), 
         .Z(n121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i121_3_lut.init = 16'hcaca;
    LUT4 i4962_3_lut (.A(dr_3__N_1864[34]), .B(dr_3__N_1864[31]), .C(\alu_op[2] ), 
         .Z(n7278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i4962_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i117_3_lut (.A(n51), .B(n53), .C(\shift_amt[1] ), 
         .Z(n117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i117_3_lut.init = 16'hcaca;
    PFUMX i22952 (.BLUT(n25289), .ALUT(n25290), .C0(n25700), .Z(n25295));
    LUT4 top_bit_I_0_i36_3_lut (.A(a_for_shift_right_c[4]), .B(a_for_shift_right_c[5]), 
         .C(shift_amt[0]), .Z(n36)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i36_3_lut.init = 16'hcaca;
    PFUMX i22920 (.BLUT(n25255), .ALUT(n25256), .C0(shift_amt_c[2]), .Z(n25263));
    LUT4 top_bit_I_0_i113_3_lut (.A(n47), .B(n49), .C(\shift_amt[1] ), 
         .Z(n113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i113_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i109_3_lut (.A(n43), .B(n45), .C(\shift_amt[1] ), 
         .Z(n109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i109_3_lut.init = 16'hcaca;
    PFUMX i22921 (.BLUT(n25257), .ALUT(n25258), .C0(shift_amt_c[2]), .Z(n25264));
    PFUMX i22922 (.BLUT(n25259), .ALUT(n25260), .C0(shift_amt_c[2]), .Z(n25265));
    PFUMX i22923 (.BLUT(n25261), .ALUT(n25262), .C0(shift_amt_c[2]), .Z(n25266));
    PFUMX i22935 (.BLUT(n25270), .ALUT(n25271), .C0(n25701), .Z(n25278));
    LUT4 top_bit_I_0_i38_3_lut (.A(a_for_shift_right_c[6]), .B(a_for_shift_right_c[7]), 
         .C(shift_amt[0]), .Z(n38)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i38_3_lut.init = 16'hcaca;
    PFUMX i22953 (.BLUT(n25291), .ALUT(n25292), .C0(n25699), .Z(n25296));
    PFUMX i22936 (.BLUT(n25272), .ALUT(n25273), .C0(n25701), .Z(n25279));
    PFUMX i22937 (.BLUT(n25274), .ALUT(n25275), .C0(n25700), .Z(n25280));
    PFUMX i22938 (.BLUT(n25276), .ALUT(n25277), .C0(n25700), .Z(n25281));
    LUT4 i22934_3_lut (.A(n61), .B(n63), .C(\shift_amt[1] ), .Z(n25277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22934_3_lut.init = 16'hcaca;
    LUT4 i22933_3_lut (.A(n57), .B(n59), .C(\shift_amt[1] ), .Z(n25276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22933_3_lut.init = 16'hcaca;
    LUT4 i22932_3_lut (.A(n53), .B(n55), .C(\shift_amt[1] ), .Z(n25275)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22932_3_lut.init = 16'hcaca;
    LUT4 i22931_3_lut (.A(n49), .B(n51), .C(\shift_amt[1] ), .Z(n25274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22931_3_lut.init = 16'hcaca;
    LUT4 i22930_3_lut (.A(n45), .B(n47), .C(\shift_amt[1] ), .Z(n25273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22930_3_lut.init = 16'hcaca;
    LUT4 i22929_3_lut (.A(n41), .B(n43), .C(\shift_amt[1] ), .Z(n25272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22929_3_lut.init = 16'hcaca;
    LUT4 i23409_2_lut_rep_711 (.A(\counter_hi[2] ), .B(\alu_op[2] ), .Z(n27336)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i23409_2_lut_rep_711.init = 16'h6666;
    LUT4 i4027_rep_132_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op[2] ), 
         .C(\shift_amt[2]_adj_1 ), .Z(n25701)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4027_rep_132_2_lut_3_lut.init = 16'h6969;
    LUT4 i4027_rep_131_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op[2] ), 
         .C(\shift_amt[2]_adj_1 ), .Z(n25700)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4027_rep_131_2_lut_3_lut.init = 16'h6969;
    LUT4 i4027_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op[2] ), .C(\shift_amt[2]_adj_1 ), 
         .Z(shift_amt_c[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4027_2_lut_3_lut.init = 16'h6969;
    LUT4 i4027_rep_130_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op[2] ), 
         .C(\shift_amt[2]_adj_1 ), .Z(n25699)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4027_rep_130_2_lut_3_lut.init = 16'h6969;
    LUT4 i22948_3_lut (.A(n58), .B(n60), .C(\shift_amt[1] ), .Z(n25291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22948_3_lut.init = 16'hcaca;
    LUT4 i22947_3_lut (.A(n54), .B(n56), .C(\shift_amt[1] ), .Z(n25290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22947_3_lut.init = 16'hcaca;
    LUT4 i22928_3_lut (.A(n37), .B(n39), .C(\shift_amt[1] ), .Z(n25271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22928_3_lut.init = 16'hcaca;
    LUT4 i22927_3_lut (.A(n33), .B(n35), .C(\shift_amt[1] ), .Z(n25270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22927_3_lut.init = 16'hcaca;
    LUT4 i22919_3_lut (.A(n60), .B(n62), .C(\shift_amt[1] ), .Z(n25262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22919_3_lut.init = 16'hcaca;
    LUT4 i22918_3_lut (.A(n56), .B(n58), .C(\shift_amt[1] ), .Z(n25261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22918_3_lut.init = 16'hcaca;
    PFUMX i22958 (.BLUT(n109), .ALUT(n113), .C0(n25699), .Z(n25301));
    LUT4 i22917_3_lut (.A(n52), .B(n54), .C(\shift_amt[1] ), .Z(n25260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22917_3_lut.init = 16'hcaca;
    LUT4 i22916_3_lut (.A(n48), .B(n50), .C(\shift_amt[1] ), .Z(n25259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22916_3_lut.init = 16'hcaca;
    LUT4 i22915_3_lut (.A(n44), .B(n46), .C(\shift_amt[1] ), .Z(n25258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22915_3_lut.init = 16'hcaca;
    LUT4 i22914_3_lut (.A(n40), .B(n42), .C(\shift_amt[1] ), .Z(n25257)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22914_3_lut.init = 16'hcaca;
    LUT4 i22913_3_lut (.A(n36), .B(n38), .C(\shift_amt[1] ), .Z(n25256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22913_3_lut.init = 16'hcaca;
    LUT4 i22912_3_lut (.A(n32), .B(n34), .C(\shift_amt[1] ), .Z(n25255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22912_3_lut.init = 16'hcaca;
    LUT4 i22946_3_lut (.A(n50), .B(n52), .C(\shift_amt[1] ), .Z(n25289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22946_3_lut.init = 16'hcaca;
    PFUMX i22959 (.BLUT(n117), .ALUT(n121), .C0(n25699), .Z(n25302));
    LUT4 i22945_3_lut (.A(n46), .B(n48), .C(\shift_amt[1] ), .Z(n25288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22945_3_lut.init = 16'hcaca;
    LUT4 i22944_3_lut (.A(n42), .B(n44), .C(\shift_amt[1] ), .Z(n25287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22944_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i40_3_lut (.A(a_for_shift_right_c[8]), .B(a_for_shift_right_c[9]), 
         .C(shift_amt[0]), .Z(n40)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i40_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i35_3_lut (.A(a_for_shift_right_c[3]), .B(a_for_shift_right_c[4]), 
         .C(shift_amt[0]), .Z(n35)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i35_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i37_3_lut (.A(a_for_shift_right_c[5]), .B(a_for_shift_right_c[6]), 
         .C(shift_amt[0]), .Z(n37)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i37_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i6_3_lut (.A(\tmp_data[26] ), .B(\tmp_data[5] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i7_3_lut (.A(\tmp_data[25] ), .B(\tmp_data[6] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i4_3_lut (.A(\tmp_data[28] ), .B(\tmp_data[3] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i5_3_lut (.A(\tmp_data[27] ), .B(\tmp_data[4] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i39_3_lut (.A(a_for_shift_right_c[7]), .B(a_for_shift_right_c[8]), 
         .C(shift_amt[0]), .Z(n39)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i39_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i41_3_lut (.A(a_for_shift_right_c[9]), .B(a_for_shift_right_c[10]), 
         .C(shift_amt[0]), .Z(n41)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i41_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i10_3_lut (.A(\tmp_data[22] ), .B(\tmp_data[9] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i11_3_lut (.A(\tmp_data[21] ), .B(\tmp_data[10] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i8_3_lut (.A(\tmp_data[24] ), .B(\tmp_data[7] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i9_3_lut (.A(\tmp_data[23] ), .B(\tmp_data[8] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i9_3_lut.init = 16'hcaca;
    PFUMX i22960 (.BLUT(n125), .ALUT(n129), .C0(n25699), .Z(n25303));
    LUT4 i4047_3_lut_4_lut (.A(n28571), .B(\alu_op[2] ), .C(n4), .D(\shift_amt[4]_adj_3 ), 
         .Z(\shift_amt[5] )) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4047_3_lut_4_lut.init = 16'hf990;
    LUT4 i2_3_lut_4_lut_adj_241 (.A(\counter_hi[4] ), .B(\alu_op[2] ), .C(n4), 
         .D(\shift_amt[4]_adj_3 ), .Z(shift_amt_c[4])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i2_3_lut_4_lut_adj_241.init = 16'h9669;
    LUT4 i22943_3_lut (.A(n38), .B(n40), .C(\shift_amt[1] ), .Z(n25286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22943_3_lut.init = 16'hcaca;
    LUT4 i22942_3_lut (.A(n34), .B(n36), .C(\shift_amt[1] ), .Z(n25285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22942_3_lut.init = 16'hcaca;
    LUT4 i23411_2_lut (.A(n28573), .B(\alu_op[2] ), .Z(n25387)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i23411_2_lut.init = 16'h6666;
    LUT4 top_bit_I_0_i105_3_lut (.A(n39), .B(n41), .C(\shift_amt[1] ), 
         .Z(n105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i105_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i101_3_lut (.A(n35), .B(n37), .C(\shift_amt[1] ), 
         .Z(n101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i101_3_lut.init = 16'hcaca;
    L6MUX21 i22956 (.D0(n25297), .D1(n25298), .SD(shift_amt_c[4]), .Z(\dr_3__N_1864[33] ));
    L6MUX21 i22963 (.D0(n25304), .D1(n25305), .SD(shift_amt_c[4]), .Z(dr_3__N_1864[34]));
    L6MUX21 i22926 (.D0(n25267), .D1(n25268), .SD(shift_amt_c[4]), .Z(dr_3__N_1864[31]));
    L6MUX21 i22941 (.D0(n25282), .D1(n25283), .SD(shift_amt_c[4]), .Z(\dr_3__N_1864[32] ));
    LUT4 top_bit_I_0_i42_3_lut (.A(a_for_shift_right_c[10]), .B(a_for_shift_right_c[11]), 
         .C(shift_amt[0]), .Z(n42)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i42_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i44_3_lut (.A(a_for_shift_right_c[12]), .B(a_for_shift_right_c[13]), 
         .C(shift_amt[0]), .Z(n44)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i44_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i13_3_lut (.A(\tmp_data[19] ), .B(\tmp_data[12] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i14_3_lut (.A(\tmp_data[18] ), .B(\tmp_data[13] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i12_3_lut (.A(\tmp_data[20] ), .B(\tmp_data[11] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i46_3_lut (.A(a_for_shift_right_c[14]), .B(a_for_shift_right_c[15]), 
         .C(shift_amt[0]), .Z(n46)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i46_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i16_3_lut (.A(\tmp_data[16] ), .B(\tmp_data[15] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i16_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i48_3_lut (.A(a_for_shift_right_c[16]), .B(a_for_shift_right_c[17]), 
         .C(shift_amt[0]), .Z(n48)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i48_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i17_3_lut (.A(\tmp_data[15] ), .B(\tmp_data[16] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i18_3_lut (.A(\tmp_data[14] ), .B(\tmp_data[17] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i15_3_lut (.A(\tmp_data[17] ), .B(\tmp_data[14] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i50_3_lut (.A(a_for_shift_right_c[18]), .B(a_for_shift_right_c[19]), 
         .C(shift_amt[0]), .Z(n50)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i50_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i52_3_lut (.A(a_for_shift_right_c[20]), .B(a_for_shift_right_c[21]), 
         .C(shift_amt[0]), .Z(n52)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i52_3_lut.init = 16'hcaca;
    L6MUX21 i22954 (.D0(n25293), .D1(n25294), .SD(shift_amt_c[3]), .Z(n25297));
    LUT4 a_0__I_0_i21_3_lut (.A(\tmp_data[11] ), .B(\tmp_data[20] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i21_3_lut.init = 16'hcaca;
    L6MUX21 i22955 (.D0(n25295), .D1(n25296), .SD(shift_amt_c[3]), .Z(n25298));
    LUT4 a_0__I_0_i22_3_lut (.A(\tmp_data[10] ), .B(\tmp_data[21] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i19_3_lut (.A(\tmp_data[13] ), .B(\tmp_data[18] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i20_3_lut (.A(\tmp_data[12] ), .B(\tmp_data[19] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i20_3_lut.init = 16'hcaca;
    L6MUX21 i22961 (.D0(n25300), .D1(n25301), .SD(shift_amt_c[3]), .Z(n25304));
    LUT4 top_bit_I_0_i54_3_lut (.A(a_for_shift_right_c[22]), .B(a_for_shift_right_c[23]), 
         .C(shift_amt[0]), .Z(n54)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i54_3_lut.init = 16'hcaca;
    L6MUX21 i22962 (.D0(n25302), .D1(n25303), .SD(shift_amt_c[3]), .Z(n25305));
    LUT4 top_bit_I_0_i56_3_lut (.A(a_for_shift_right_c[24]), .B(a_for_shift_right_c[25]), 
         .C(shift_amt[0]), .Z(n56)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i56_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i25_3_lut (.A(\tmp_data[7] ), .B(\tmp_data[24] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i26_3_lut (.A(\tmp_data[6] ), .B(\tmp_data[25] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i23_3_lut (.A(\tmp_data[9] ), .B(\tmp_data[22] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i24_3_lut (.A(\tmp_data[8] ), .B(\tmp_data[23] ), .C(\alu_op[2] ), 
         .Z(a_for_shift_right_c[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i24_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module tinyqv_registers
//

module tinyqv_registers (rs1, rd, debug_reg_wen, rs2, clk_c, return_addr, 
            debug_rd, \reg_access[4][3] , data_rs1, n28571, n28573, 
            \counter_hi[2] , data_rs2, n28580, n27231, n24605, \mie[12] , 
            n928, \reg_access[3][2] , n28581, n27205, n27113, any_additional_mem_ops, 
            n2356, \mie[8] , n895, \mie[4] , n862) /* synthesis syn_module_defined=1 */ ;
    input [3:0]rs1;
    input [3:0]rd;
    input debug_reg_wen;
    input [3:0]rs2;
    input clk_c;
    output [23:1]return_addr;
    input [3:0]debug_rd;
    output \reg_access[4][3] ;
    output [3:0]data_rs1;
    input n28571;
    input n28573;
    input \counter_hi[2] ;
    output [3:0]data_rs2;
    output n28580;
    input n27231;
    input n24605;
    input \mie[12] ;
    output n928;
    output \reg_access[3][2] ;
    output n28581;
    input n27205;
    input n27113;
    input any_additional_mem_ops;
    output n2356;
    input \mie[8] ;
    output n895;
    input \mie[4] ;
    output n862;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [31:0]\registers[14] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[15] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n25247, n27118, n27117, n27116, n27115;
    wire [31:0]\registers[12] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[13] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n25246;
    wire [31:0]\registers[10] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[11] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n25245;
    wire [31:0]\registers[8] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[9] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n25244;
    wire [31:0]\registers[6] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[7] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n25243;
    wire [31:0]\registers[5] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n25242, n25225, n25224, n25223, n25222, n25221, n25220, 
        n25210, n25209, n25208, n25207, n25206, n25205, n25160, 
        n25161, n25168, n25203, n25204, n25211, n25218, n25219, 
        n25226;
    wire [31:0]\registers[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_1__2__N_1756, registers_1__1__N_1757, registers_1__0__N_1758;
    wire [31:0]\registers[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_2__3__N_1759, registers_2__2__N_1762, registers_2__1__N_1763, 
        registers_2__0__N_1764, registers_5__3__N_1765, registers_5__2__N_1768, 
        registers_5__1__N_1769, registers_5__0__N_1770, registers_6__3__N_1771, 
        registers_6__2__N_1774, registers_6__1__N_1775, registers_6__0__N_1776, 
        registers_7__3__N_1777, registers_7__2__N_1780, registers_7__1__N_1781, 
        registers_7__0__N_1782, registers_8__3__N_1783, registers_8__2__N_1786, 
        registers_8__1__N_1787, registers_8__0__N_1788, registers_9__3__N_1789, 
        registers_9__2__N_1792, registers_9__1__N_1793, registers_9__0__N_1794, 
        registers_10__3__N_1795, registers_10__2__N_1798, registers_10__1__N_1799, 
        registers_10__0__N_1800, registers_11__3__N_1801, registers_11__2__N_1804, 
        registers_11__1__N_1805, registers_11__0__N_1806, registers_12__3__N_1807, 
        registers_12__2__N_1810, registers_12__1__N_1811, registers_12__0__N_1812, 
        registers_13__3__N_1813, registers_13__2__N_1816, registers_13__1__N_1817, 
        registers_13__0__N_1818, registers_14__3__N_1819, registers_14__2__N_1822, 
        registers_14__1__N_1823, registers_14__0__N_1824, registers_15__3__N_1825, 
        registers_15__2__N_1828, registers_15__1__N_1829, registers_15__0__N_1830, 
        registers_1__3__N_1753, n25167, n25166, n25165, n25164, n25163, 
        n25162, n12, n11, n9, n8, n5, n5_adj_2600, n12_adj_2601, 
        n11_adj_2602, n9_adj_2603, n8_adj_2604, n5_adj_2605, n27315, 
        n4, n25315, n5_adj_2606, n25311, n25312, n27316, n4_adj_2607, 
        n25308, n12_adj_2608, n11_adj_2609, n9_adj_2610, n8_adj_2611, 
        n12_adj_2612, n27317, n11_adj_2613, n9_adj_2614, n8_adj_2615, 
        n25240, n25241, n25248, n27318, n25230, n25231, n25318, 
        n25319, n25309, n25310, n25316, n25317, n25314, n25307, 
        n25146, n25147, n25150, n25148, n25149, n25151, n25153, 
        n25154, n25157, n25155, n25156, n25158, n25170, n25171, 
        n25173, n25213, n25214, n25216, n25228, n25229, n25250, 
        n25251, n25253, n25169, n25212, n25227, n25172, n25215, 
        n25252, n25249;
    
    LUT4 i22904_3_lut (.A(\registers[14] [6]), .B(\registers[15] [6]), .C(rs1[0]), 
         .Z(n25247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22904_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_493_3_lut (.A(rd[0]), .B(debug_reg_wen), .C(rd[1]), 
         .Z(n27118)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_493_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_492_3_lut (.A(rd[0]), .B(rd[1]), .C(debug_reg_wen), 
         .Z(n27117)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_rep_492_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_491_3_lut (.A(rd[0]), .B(rd[1]), .C(debug_reg_wen), 
         .Z(n27116)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_491_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_490_3_lut (.A(rd[0]), .B(debug_reg_wen), .C(rd[1]), 
         .Z(n27115)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_rep_490_3_lut.init = 16'h0404;
    LUT4 i22903_3_lut (.A(\registers[12] [6]), .B(\registers[13] [6]), .C(rs1[0]), 
         .Z(n25246)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22903_3_lut.init = 16'hcaca;
    LUT4 i22902_3_lut (.A(\registers[10] [6]), .B(\registers[11] [6]), .C(rs1[0]), 
         .Z(n25245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22902_3_lut.init = 16'hcaca;
    LUT4 i22901_3_lut (.A(\registers[8] [6]), .B(\registers[9] [6]), .C(rs1[0]), 
         .Z(n25244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22901_3_lut.init = 16'hcaca;
    LUT4 i22900_3_lut (.A(\registers[6] [6]), .B(\registers[7] [6]), .C(rs1[0]), 
         .Z(n25243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22900_3_lut.init = 16'hcaca;
    LUT4 i22899_3_lut (.A(\registers[5] [6]), .B(rs1[0]), .Z(n25242)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22899_3_lut.init = 16'h8888;
    LUT4 i22882_3_lut (.A(\registers[14] [4]), .B(\registers[15] [4]), .C(rs1[0]), 
         .Z(n25225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22882_3_lut.init = 16'hcaca;
    LUT4 i22881_3_lut (.A(\registers[12] [4]), .B(\registers[13] [4]), .C(rs1[0]), 
         .Z(n25224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22881_3_lut.init = 16'hcaca;
    LUT4 i22880_3_lut (.A(\registers[10] [4]), .B(\registers[11] [4]), .C(rs1[0]), 
         .Z(n25223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22880_3_lut.init = 16'hcaca;
    LUT4 i22879_3_lut (.A(\registers[8] [4]), .B(\registers[9] [4]), .C(rs1[0]), 
         .Z(n25222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22879_3_lut.init = 16'hcaca;
    LUT4 i22878_3_lut (.A(\registers[6] [4]), .B(\registers[7] [4]), .C(rs1[0]), 
         .Z(n25221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22878_3_lut.init = 16'hcaca;
    LUT4 i22877_3_lut (.A(\registers[5] [4]), .B(rs1[0]), .Z(n25220)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22877_3_lut.init = 16'h8888;
    LUT4 i22867_3_lut (.A(\registers[14] [4]), .B(\registers[15] [4]), .C(rs2[0]), 
         .Z(n25210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22867_3_lut.init = 16'hcaca;
    LUT4 i22866_3_lut (.A(\registers[12] [4]), .B(\registers[13] [4]), .C(rs2[0]), 
         .Z(n25209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22866_3_lut.init = 16'hcaca;
    LUT4 i22865_3_lut (.A(\registers[10] [4]), .B(\registers[11] [4]), .C(rs2[0]), 
         .Z(n25208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22865_3_lut.init = 16'hcaca;
    LUT4 i22864_3_lut (.A(\registers[8] [4]), .B(\registers[9] [4]), .C(rs2[0]), 
         .Z(n25207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22864_3_lut.init = 16'hcaca;
    LUT4 i22863_3_lut (.A(\registers[6] [4]), .B(\registers[7] [4]), .C(rs2[0]), 
         .Z(n25206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22863_3_lut.init = 16'hcaca;
    LUT4 i22862_3_lut (.A(\registers[5] [4]), .B(rs2[0]), .Z(n25205)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22862_3_lut.init = 16'h8888;
    PFUMX i22825 (.BLUT(n25160), .ALUT(n25161), .C0(rs2[1]), .Z(n25168));
    PFUMX i22868 (.BLUT(n25203), .ALUT(n25204), .C0(rs2[1]), .Z(n25211));
    PFUMX i22883 (.BLUT(n25218), .ALUT(n25219), .C0(rs1[1]), .Z(n25226));
    FD1S3AX \registers_1[[2__504  (.D(registers_1__2__N_1756), .CK(clk_c), 
            .Q(\registers[1] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[2__504 .GSR = "DISABLED";
    FD1S3AX \registers_1[[1__505  (.D(registers_1__1__N_1757), .CK(clk_c), 
            .Q(\registers[1] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[1__505 .GSR = "DISABLED";
    FD1S3AX \registers_1[[0__506  (.D(registers_1__0__N_1758), .CK(clk_c), 
            .Q(\registers[1] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[0__506 .GSR = "DISABLED";
    FD1S3AX \registers_1[[31__507  (.D(\registers[1] [3]), .CK(clk_c), .Q(return_addr[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[31__507 .GSR = "DISABLED";
    FD1S3AX \registers_1[[30__508  (.D(\registers[1] [2]), .CK(clk_c), .Q(return_addr[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[30__508 .GSR = "DISABLED";
    FD1S3AX \registers_1[[29__509  (.D(\registers[1] [1]), .CK(clk_c), .Q(return_addr[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[29__509 .GSR = "DISABLED";
    FD1S3AX \registers_1[[28__510  (.D(\registers[1] [0]), .CK(clk_c), .Q(return_addr[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[28__510 .GSR = "DISABLED";
    FD1S3AX \registers_1[[27__511  (.D(return_addr[23]), .CK(clk_c), .Q(return_addr[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[27__511 .GSR = "DISABLED";
    FD1S3AX \registers_1[[26__512  (.D(return_addr[22]), .CK(clk_c), .Q(return_addr[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[26__512 .GSR = "DISABLED";
    FD1S3AX \registers_1[[25__513  (.D(return_addr[21]), .CK(clk_c), .Q(return_addr[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[25__513 .GSR = "DISABLED";
    FD1S3AX \registers_1[[24__514  (.D(return_addr[20]), .CK(clk_c), .Q(return_addr[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[24__514 .GSR = "DISABLED";
    FD1S3AX \registers_1[[23__515  (.D(return_addr[19]), .CK(clk_c), .Q(return_addr[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[23__515 .GSR = "DISABLED";
    FD1S3AX \registers_1[[22__516  (.D(return_addr[18]), .CK(clk_c), .Q(return_addr[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[22__516 .GSR = "DISABLED";
    FD1S3AX \registers_1[[21__517  (.D(return_addr[17]), .CK(clk_c), .Q(return_addr[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[21__517 .GSR = "DISABLED";
    FD1S3AX \registers_1[[20__518  (.D(return_addr[16]), .CK(clk_c), .Q(return_addr[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[20__518 .GSR = "DISABLED";
    FD1S3AX \registers_1[[19__519  (.D(return_addr[15]), .CK(clk_c), .Q(return_addr[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[19__519 .GSR = "DISABLED";
    FD1S3AX \registers_1[[18__520  (.D(return_addr[14]), .CK(clk_c), .Q(return_addr[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[18__520 .GSR = "DISABLED";
    FD1S3AX \registers_1[[17__521  (.D(return_addr[13]), .CK(clk_c), .Q(return_addr[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[17__521 .GSR = "DISABLED";
    FD1S3AX \registers_1[[16__522  (.D(return_addr[12]), .CK(clk_c), .Q(return_addr[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[16__522 .GSR = "DISABLED";
    FD1S3AX \registers_1[[15__523  (.D(return_addr[11]), .CK(clk_c), .Q(return_addr[7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[15__523 .GSR = "DISABLED";
    FD1S3AX \registers_1[[14__524  (.D(return_addr[10]), .CK(clk_c), .Q(return_addr[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[14__524 .GSR = "DISABLED";
    FD1S3AX \registers_1[[13__525  (.D(return_addr[9]), .CK(clk_c), .Q(return_addr[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[13__525 .GSR = "DISABLED";
    FD1S3AX \registers_1[[12__526  (.D(return_addr[8]), .CK(clk_c), .Q(return_addr[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[12__526 .GSR = "DISABLED";
    FD1S3AX \registers_1[[11__527  (.D(return_addr[7]), .CK(clk_c), .Q(return_addr[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[11__527 .GSR = "DISABLED";
    FD1S3AX \registers_1[[10__528  (.D(return_addr[6]), .CK(clk_c), .Q(return_addr[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[10__528 .GSR = "DISABLED";
    FD1S3AX \registers_1[[9__529  (.D(return_addr[5]), .CK(clk_c), .Q(return_addr[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[9__529 .GSR = "DISABLED";
    FD1S3AX \registers_1[[8__530  (.D(return_addr[4]), .CK(clk_c), .Q(\registers[1] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[8__530 .GSR = "DISABLED";
    FD1S3AX \registers_1[[7__531  (.D(return_addr[3]), .CK(clk_c), .Q(\registers[1] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[7__531 .GSR = "DISABLED";
    FD1S3AX \registers_1[[6__532  (.D(return_addr[2]), .CK(clk_c), .Q(\registers[1] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[6__532 .GSR = "DISABLED";
    FD1S3AX \registers_1[[5__533  (.D(return_addr[1]), .CK(clk_c), .Q(\registers[1] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[5__533 .GSR = "DISABLED";
    FD1S3AX \registers_1[[4__534  (.D(\registers[1] [8]), .CK(clk_c), .Q(\registers[1] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[4__534 .GSR = "DISABLED";
    FD1S3AX \registers_2[[3__535  (.D(registers_2__3__N_1759), .CK(clk_c), 
            .Q(\registers[2] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[3__535 .GSR = "DISABLED";
    FD1S3AX \registers_2[[2__536  (.D(registers_2__2__N_1762), .CK(clk_c), 
            .Q(\registers[2] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[2__536 .GSR = "DISABLED";
    FD1S3AX \registers_2[[1__537  (.D(registers_2__1__N_1763), .CK(clk_c), 
            .Q(\registers[2] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[1__537 .GSR = "DISABLED";
    FD1S3AX \registers_2[[0__538  (.D(registers_2__0__N_1764), .CK(clk_c), 
            .Q(\registers[2] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[0__538 .GSR = "DISABLED";
    FD1S3AX \registers_2[[31__539  (.D(\registers[2] [3]), .CK(clk_c), .Q(\registers[2] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[31__539 .GSR = "DISABLED";
    FD1S3AX \registers_2[[30__540  (.D(\registers[2] [2]), .CK(clk_c), .Q(\registers[2] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[30__540 .GSR = "DISABLED";
    FD1S3AX \registers_2[[29__541  (.D(\registers[2] [1]), .CK(clk_c), .Q(\registers[2] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[29__541 .GSR = "DISABLED";
    FD1S3AX \registers_2[[28__542  (.D(\registers[2] [0]), .CK(clk_c), .Q(\registers[2] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[28__542 .GSR = "DISABLED";
    FD1S3AX \registers_2[[27__543  (.D(\registers[2] [31]), .CK(clk_c), 
            .Q(\registers[2] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[27__543 .GSR = "DISABLED";
    FD1S3AX \registers_2[[26__544  (.D(\registers[2] [30]), .CK(clk_c), 
            .Q(\registers[2] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[26__544 .GSR = "DISABLED";
    FD1S3AX \registers_2[[25__545  (.D(\registers[2] [29]), .CK(clk_c), 
            .Q(\registers[2] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[25__545 .GSR = "DISABLED";
    FD1S3AX \registers_2[[24__546  (.D(\registers[2] [28]), .CK(clk_c), 
            .Q(\registers[2] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[24__546 .GSR = "DISABLED";
    FD1S3AX \registers_2[[23__547  (.D(\registers[2] [27]), .CK(clk_c), 
            .Q(\registers[2] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[23__547 .GSR = "DISABLED";
    FD1S3AX \registers_2[[22__548  (.D(\registers[2] [26]), .CK(clk_c), 
            .Q(\registers[2] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[22__548 .GSR = "DISABLED";
    FD1S3AX \registers_2[[21__549  (.D(\registers[2] [25]), .CK(clk_c), 
            .Q(\registers[2] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[21__549 .GSR = "DISABLED";
    FD1S3AX \registers_2[[20__550  (.D(\registers[2] [24]), .CK(clk_c), 
            .Q(\registers[2] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[20__550 .GSR = "DISABLED";
    FD1S3AX \registers_2[[19__551  (.D(\registers[2] [23]), .CK(clk_c), 
            .Q(\registers[2] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[19__551 .GSR = "DISABLED";
    FD1S3AX \registers_2[[18__552  (.D(\registers[2] [22]), .CK(clk_c), 
            .Q(\registers[2] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[18__552 .GSR = "DISABLED";
    FD1S3AX \registers_2[[17__553  (.D(\registers[2] [21]), .CK(clk_c), 
            .Q(\registers[2] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[17__553 .GSR = "DISABLED";
    FD1S3AX \registers_2[[16__554  (.D(\registers[2] [20]), .CK(clk_c), 
            .Q(\registers[2] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[16__554 .GSR = "DISABLED";
    FD1S3AX \registers_2[[15__555  (.D(\registers[2] [19]), .CK(clk_c), 
            .Q(\registers[2] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[15__555 .GSR = "DISABLED";
    FD1S3AX \registers_2[[14__556  (.D(\registers[2] [18]), .CK(clk_c), 
            .Q(\registers[2] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[14__556 .GSR = "DISABLED";
    FD1S3AX \registers_2[[13__557  (.D(\registers[2] [17]), .CK(clk_c), 
            .Q(\registers[2] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[13__557 .GSR = "DISABLED";
    FD1S3AX \registers_2[[12__558  (.D(\registers[2] [16]), .CK(clk_c), 
            .Q(\registers[2] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[12__558 .GSR = "DISABLED";
    FD1S3AX \registers_2[[11__559  (.D(\registers[2] [15]), .CK(clk_c), 
            .Q(\registers[2] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[11__559 .GSR = "DISABLED";
    FD1S3AX \registers_2[[10__560  (.D(\registers[2] [14]), .CK(clk_c), 
            .Q(\registers[2] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[10__560 .GSR = "DISABLED";
    FD1S3AX \registers_2[[9__561  (.D(\registers[2] [13]), .CK(clk_c), .Q(\registers[2] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[9__561 .GSR = "DISABLED";
    FD1S3AX \registers_2[[8__562  (.D(\registers[2] [12]), .CK(clk_c), .Q(\registers[2] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[8__562 .GSR = "DISABLED";
    FD1S3AX \registers_2[[7__563  (.D(\registers[2] [11]), .CK(clk_c), .Q(\registers[2] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[7__563 .GSR = "DISABLED";
    FD1S3AX \registers_2[[6__564  (.D(\registers[2] [10]), .CK(clk_c), .Q(\registers[2] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[6__564 .GSR = "DISABLED";
    FD1S3AX \registers_2[[5__565  (.D(\registers[2] [9]), .CK(clk_c), .Q(\registers[2] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[5__565 .GSR = "DISABLED";
    FD1S3AX \registers_2[[4__566  (.D(\registers[2] [8]), .CK(clk_c), .Q(\registers[2] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[4__566 .GSR = "DISABLED";
    FD1S3AX \registers_5[[3__567  (.D(registers_5__3__N_1765), .CK(clk_c), 
            .Q(\registers[5] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[3__567 .GSR = "DISABLED";
    FD1S3AX \registers_5[[2__568  (.D(registers_5__2__N_1768), .CK(clk_c), 
            .Q(\registers[5] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[2__568 .GSR = "DISABLED";
    FD1S3AX \registers_5[[1__569  (.D(registers_5__1__N_1769), .CK(clk_c), 
            .Q(\registers[5] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[1__569 .GSR = "DISABLED";
    FD1S3AX \registers_5[[0__570  (.D(registers_5__0__N_1770), .CK(clk_c), 
            .Q(\registers[5] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[0__570 .GSR = "DISABLED";
    FD1S3AX \registers_5[[31__571  (.D(\registers[5] [3]), .CK(clk_c), .Q(\registers[5] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[31__571 .GSR = "DISABLED";
    FD1S3AX \registers_5[[30__572  (.D(\registers[5] [2]), .CK(clk_c), .Q(\registers[5] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[30__572 .GSR = "DISABLED";
    FD1S3AX \registers_5[[29__573  (.D(\registers[5] [1]), .CK(clk_c), .Q(\registers[5] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[29__573 .GSR = "DISABLED";
    FD1S3AX \registers_5[[28__574  (.D(\registers[5] [0]), .CK(clk_c), .Q(\registers[5] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[28__574 .GSR = "DISABLED";
    FD1S3AX \registers_5[[27__575  (.D(\registers[5] [31]), .CK(clk_c), 
            .Q(\registers[5] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[27__575 .GSR = "DISABLED";
    FD1S3AX \registers_5[[26__576  (.D(\registers[5] [30]), .CK(clk_c), 
            .Q(\registers[5] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[26__576 .GSR = "DISABLED";
    FD1S3AX \registers_5[[25__577  (.D(\registers[5] [29]), .CK(clk_c), 
            .Q(\registers[5] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[25__577 .GSR = "DISABLED";
    FD1S3AX \registers_5[[24__578  (.D(\registers[5] [28]), .CK(clk_c), 
            .Q(\registers[5] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[24__578 .GSR = "DISABLED";
    FD1S3AX \registers_5[[23__579  (.D(\registers[5] [27]), .CK(clk_c), 
            .Q(\registers[5] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[23__579 .GSR = "DISABLED";
    FD1S3AX \registers_5[[22__580  (.D(\registers[5] [26]), .CK(clk_c), 
            .Q(\registers[5] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[22__580 .GSR = "DISABLED";
    FD1S3AX \registers_5[[21__581  (.D(\registers[5] [25]), .CK(clk_c), 
            .Q(\registers[5] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[21__581 .GSR = "DISABLED";
    FD1S3AX \registers_5[[20__582  (.D(\registers[5] [24]), .CK(clk_c), 
            .Q(\registers[5] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[20__582 .GSR = "DISABLED";
    FD1S3AX \registers_5[[19__583  (.D(\registers[5] [23]), .CK(clk_c), 
            .Q(\registers[5] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[19__583 .GSR = "DISABLED";
    FD1S3AX \registers_5[[18__584  (.D(\registers[5] [22]), .CK(clk_c), 
            .Q(\registers[5] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[18__584 .GSR = "DISABLED";
    FD1S3AX \registers_5[[17__585  (.D(\registers[5] [21]), .CK(clk_c), 
            .Q(\registers[5] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[17__585 .GSR = "DISABLED";
    FD1S3AX \registers_5[[16__586  (.D(\registers[5] [20]), .CK(clk_c), 
            .Q(\registers[5] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[16__586 .GSR = "DISABLED";
    FD1S3AX \registers_5[[15__587  (.D(\registers[5] [19]), .CK(clk_c), 
            .Q(\registers[5] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[15__587 .GSR = "DISABLED";
    FD1S3AX \registers_5[[14__588  (.D(\registers[5] [18]), .CK(clk_c), 
            .Q(\registers[5] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[14__588 .GSR = "DISABLED";
    FD1S3AX \registers_5[[13__589  (.D(\registers[5] [17]), .CK(clk_c), 
            .Q(\registers[5] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[13__589 .GSR = "DISABLED";
    FD1S3AX \registers_5[[12__590  (.D(\registers[5] [16]), .CK(clk_c), 
            .Q(\registers[5] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[12__590 .GSR = "DISABLED";
    FD1S3AX \registers_5[[11__591  (.D(\registers[5] [15]), .CK(clk_c), 
            .Q(\registers[5] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[11__591 .GSR = "DISABLED";
    FD1S3AX \registers_5[[10__592  (.D(\registers[5] [14]), .CK(clk_c), 
            .Q(\registers[5] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[10__592 .GSR = "DISABLED";
    FD1S3AX \registers_5[[9__593  (.D(\registers[5] [13]), .CK(clk_c), .Q(\registers[5] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[9__593 .GSR = "DISABLED";
    FD1S3AX \registers_5[[8__594  (.D(\registers[5] [12]), .CK(clk_c), .Q(\registers[5] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[8__594 .GSR = "DISABLED";
    FD1S3AX \registers_5[[7__595  (.D(\registers[5] [11]), .CK(clk_c), .Q(\registers[5] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[7__595 .GSR = "DISABLED";
    FD1S3AX \registers_5[[6__596  (.D(\registers[5] [10]), .CK(clk_c), .Q(\registers[5] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[6__596 .GSR = "DISABLED";
    FD1S3AX \registers_5[[5__597  (.D(\registers[5] [9]), .CK(clk_c), .Q(\registers[5] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[5__597 .GSR = "DISABLED";
    FD1S3AX \registers_5[[4__598  (.D(\registers[5] [8]), .CK(clk_c), .Q(\registers[5] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[4__598 .GSR = "DISABLED";
    FD1S3AX \registers_6[[3__599  (.D(registers_6__3__N_1771), .CK(clk_c), 
            .Q(\registers[6] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[3__599 .GSR = "DISABLED";
    FD1S3AX \registers_6[[2__600  (.D(registers_6__2__N_1774), .CK(clk_c), 
            .Q(\registers[6] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[2__600 .GSR = "DISABLED";
    FD1S3AX \registers_6[[1__601  (.D(registers_6__1__N_1775), .CK(clk_c), 
            .Q(\registers[6] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[1__601 .GSR = "DISABLED";
    FD1S3AX \registers_6[[0__602  (.D(registers_6__0__N_1776), .CK(clk_c), 
            .Q(\registers[6] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[0__602 .GSR = "DISABLED";
    FD1S3AX \registers_6[[31__603  (.D(\registers[6] [3]), .CK(clk_c), .Q(\registers[6] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[31__603 .GSR = "DISABLED";
    FD1S3AX \registers_6[[30__604  (.D(\registers[6] [2]), .CK(clk_c), .Q(\registers[6] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[30__604 .GSR = "DISABLED";
    FD1S3AX \registers_6[[29__605  (.D(\registers[6] [1]), .CK(clk_c), .Q(\registers[6] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[29__605 .GSR = "DISABLED";
    FD1S3AX \registers_6[[28__606  (.D(\registers[6] [0]), .CK(clk_c), .Q(\registers[6] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[28__606 .GSR = "DISABLED";
    FD1S3AX \registers_6[[27__607  (.D(\registers[6] [31]), .CK(clk_c), 
            .Q(\registers[6] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[27__607 .GSR = "DISABLED";
    FD1S3AX \registers_6[[26__608  (.D(\registers[6] [30]), .CK(clk_c), 
            .Q(\registers[6] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[26__608 .GSR = "DISABLED";
    FD1S3AX \registers_6[[25__609  (.D(\registers[6] [29]), .CK(clk_c), 
            .Q(\registers[6] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[25__609 .GSR = "DISABLED";
    FD1S3AX \registers_6[[24__610  (.D(\registers[6] [28]), .CK(clk_c), 
            .Q(\registers[6] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[24__610 .GSR = "DISABLED";
    FD1S3AX \registers_6[[23__611  (.D(\registers[6] [27]), .CK(clk_c), 
            .Q(\registers[6] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[23__611 .GSR = "DISABLED";
    FD1S3AX \registers_6[[22__612  (.D(\registers[6] [26]), .CK(clk_c), 
            .Q(\registers[6] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[22__612 .GSR = "DISABLED";
    FD1S3AX \registers_6[[21__613  (.D(\registers[6] [25]), .CK(clk_c), 
            .Q(\registers[6] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[21__613 .GSR = "DISABLED";
    FD1S3AX \registers_6[[20__614  (.D(\registers[6] [24]), .CK(clk_c), 
            .Q(\registers[6] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[20__614 .GSR = "DISABLED";
    FD1S3AX \registers_6[[19__615  (.D(\registers[6] [23]), .CK(clk_c), 
            .Q(\registers[6] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[19__615 .GSR = "DISABLED";
    FD1S3AX \registers_6[[18__616  (.D(\registers[6] [22]), .CK(clk_c), 
            .Q(\registers[6] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[18__616 .GSR = "DISABLED";
    FD1S3AX \registers_6[[17__617  (.D(\registers[6] [21]), .CK(clk_c), 
            .Q(\registers[6] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[17__617 .GSR = "DISABLED";
    FD1S3AX \registers_6[[16__618  (.D(\registers[6] [20]), .CK(clk_c), 
            .Q(\registers[6] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[16__618 .GSR = "DISABLED";
    FD1S3AX \registers_6[[15__619  (.D(\registers[6] [19]), .CK(clk_c), 
            .Q(\registers[6] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[15__619 .GSR = "DISABLED";
    FD1S3AX \registers_6[[14__620  (.D(\registers[6] [18]), .CK(clk_c), 
            .Q(\registers[6] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[14__620 .GSR = "DISABLED";
    FD1S3AX \registers_6[[13__621  (.D(\registers[6] [17]), .CK(clk_c), 
            .Q(\registers[6] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[13__621 .GSR = "DISABLED";
    FD1S3AX \registers_6[[12__622  (.D(\registers[6] [16]), .CK(clk_c), 
            .Q(\registers[6] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[12__622 .GSR = "DISABLED";
    FD1S3AX \registers_6[[11__623  (.D(\registers[6] [15]), .CK(clk_c), 
            .Q(\registers[6] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[11__623 .GSR = "DISABLED";
    FD1S3AX \registers_6[[10__624  (.D(\registers[6] [14]), .CK(clk_c), 
            .Q(\registers[6] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[10__624 .GSR = "DISABLED";
    FD1S3AX \registers_6[[9__625  (.D(\registers[6] [13]), .CK(clk_c), .Q(\registers[6] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[9__625 .GSR = "DISABLED";
    FD1S3AX \registers_6[[8__626  (.D(\registers[6] [12]), .CK(clk_c), .Q(\registers[6] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[8__626 .GSR = "DISABLED";
    FD1S3AX \registers_6[[7__627  (.D(\registers[6] [11]), .CK(clk_c), .Q(\registers[6] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[7__627 .GSR = "DISABLED";
    FD1S3AX \registers_6[[6__628  (.D(\registers[6] [10]), .CK(clk_c), .Q(\registers[6] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[6__628 .GSR = "DISABLED";
    FD1S3AX \registers_6[[5__629  (.D(\registers[6] [9]), .CK(clk_c), .Q(\registers[6] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[5__629 .GSR = "DISABLED";
    FD1S3AX \registers_6[[4__630  (.D(\registers[6] [8]), .CK(clk_c), .Q(\registers[6] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[4__630 .GSR = "DISABLED";
    FD1S3AX \registers_7[[3__631  (.D(registers_7__3__N_1777), .CK(clk_c), 
            .Q(\registers[7] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[3__631 .GSR = "DISABLED";
    FD1S3AX \registers_7[[2__632  (.D(registers_7__2__N_1780), .CK(clk_c), 
            .Q(\registers[7] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[2__632 .GSR = "DISABLED";
    FD1S3AX \registers_7[[1__633  (.D(registers_7__1__N_1781), .CK(clk_c), 
            .Q(\registers[7] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[1__633 .GSR = "DISABLED";
    FD1S3AX \registers_7[[0__634  (.D(registers_7__0__N_1782), .CK(clk_c), 
            .Q(\registers[7] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[0__634 .GSR = "DISABLED";
    FD1S3AX \registers_7[[31__635  (.D(\registers[7] [3]), .CK(clk_c), .Q(\registers[7] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[31__635 .GSR = "DISABLED";
    FD1S3AX \registers_7[[30__636  (.D(\registers[7] [2]), .CK(clk_c), .Q(\registers[7] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[30__636 .GSR = "DISABLED";
    FD1S3AX \registers_7[[29__637  (.D(\registers[7] [1]), .CK(clk_c), .Q(\registers[7] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[29__637 .GSR = "DISABLED";
    FD1S3AX \registers_7[[28__638  (.D(\registers[7] [0]), .CK(clk_c), .Q(\registers[7] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[28__638 .GSR = "DISABLED";
    FD1S3AX \registers_7[[27__639  (.D(\registers[7] [31]), .CK(clk_c), 
            .Q(\registers[7] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[27__639 .GSR = "DISABLED";
    FD1S3AX \registers_7[[26__640  (.D(\registers[7] [30]), .CK(clk_c), 
            .Q(\registers[7] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[26__640 .GSR = "DISABLED";
    FD1S3AX \registers_7[[25__641  (.D(\registers[7] [29]), .CK(clk_c), 
            .Q(\registers[7] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[25__641 .GSR = "DISABLED";
    FD1S3AX \registers_7[[24__642  (.D(\registers[7] [28]), .CK(clk_c), 
            .Q(\registers[7] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[24__642 .GSR = "DISABLED";
    FD1S3AX \registers_7[[23__643  (.D(\registers[7] [27]), .CK(clk_c), 
            .Q(\registers[7] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[23__643 .GSR = "DISABLED";
    FD1S3AX \registers_7[[22__644  (.D(\registers[7] [26]), .CK(clk_c), 
            .Q(\registers[7] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[22__644 .GSR = "DISABLED";
    FD1S3AX \registers_7[[21__645  (.D(\registers[7] [25]), .CK(clk_c), 
            .Q(\registers[7] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[21__645 .GSR = "DISABLED";
    FD1S3AX \registers_7[[20__646  (.D(\registers[7] [24]), .CK(clk_c), 
            .Q(\registers[7] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[20__646 .GSR = "DISABLED";
    FD1S3AX \registers_7[[19__647  (.D(\registers[7] [23]), .CK(clk_c), 
            .Q(\registers[7] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[19__647 .GSR = "DISABLED";
    FD1S3AX \registers_7[[18__648  (.D(\registers[7] [22]), .CK(clk_c), 
            .Q(\registers[7] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[18__648 .GSR = "DISABLED";
    FD1S3AX \registers_7[[17__649  (.D(\registers[7] [21]), .CK(clk_c), 
            .Q(\registers[7] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[17__649 .GSR = "DISABLED";
    FD1S3AX \registers_7[[16__650  (.D(\registers[7] [20]), .CK(clk_c), 
            .Q(\registers[7] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[16__650 .GSR = "DISABLED";
    FD1S3AX \registers_7[[15__651  (.D(\registers[7] [19]), .CK(clk_c), 
            .Q(\registers[7] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[15__651 .GSR = "DISABLED";
    FD1S3AX \registers_7[[14__652  (.D(\registers[7] [18]), .CK(clk_c), 
            .Q(\registers[7] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[14__652 .GSR = "DISABLED";
    FD1S3AX \registers_7[[13__653  (.D(\registers[7] [17]), .CK(clk_c), 
            .Q(\registers[7] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[13__653 .GSR = "DISABLED";
    FD1S3AX \registers_7[[12__654  (.D(\registers[7] [16]), .CK(clk_c), 
            .Q(\registers[7] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[12__654 .GSR = "DISABLED";
    FD1S3AX \registers_7[[11__655  (.D(\registers[7] [15]), .CK(clk_c), 
            .Q(\registers[7] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[11__655 .GSR = "DISABLED";
    FD1S3AX \registers_7[[10__656  (.D(\registers[7] [14]), .CK(clk_c), 
            .Q(\registers[7] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[10__656 .GSR = "DISABLED";
    FD1S3AX \registers_7[[9__657  (.D(\registers[7] [13]), .CK(clk_c), .Q(\registers[7] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[9__657 .GSR = "DISABLED";
    FD1S3AX \registers_7[[8__658  (.D(\registers[7] [12]), .CK(clk_c), .Q(\registers[7] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[8__658 .GSR = "DISABLED";
    FD1S3AX \registers_7[[7__659  (.D(\registers[7] [11]), .CK(clk_c), .Q(\registers[7] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[7__659 .GSR = "DISABLED";
    FD1S3AX \registers_7[[6__660  (.D(\registers[7] [10]), .CK(clk_c), .Q(\registers[7] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[6__660 .GSR = "DISABLED";
    FD1S3AX \registers_7[[5__661  (.D(\registers[7] [9]), .CK(clk_c), .Q(\registers[7] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[5__661 .GSR = "DISABLED";
    FD1S3AX \registers_7[[4__662  (.D(\registers[7] [8]), .CK(clk_c), .Q(\registers[7] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[4__662 .GSR = "DISABLED";
    FD1S3AX \registers_8[[3__663  (.D(registers_8__3__N_1783), .CK(clk_c), 
            .Q(\registers[8] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[3__663 .GSR = "DISABLED";
    FD1S3AX \registers_8[[2__664  (.D(registers_8__2__N_1786), .CK(clk_c), 
            .Q(\registers[8] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[2__664 .GSR = "DISABLED";
    FD1S3AX \registers_8[[1__665  (.D(registers_8__1__N_1787), .CK(clk_c), 
            .Q(\registers[8] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[1__665 .GSR = "DISABLED";
    FD1S3AX \registers_8[[0__666  (.D(registers_8__0__N_1788), .CK(clk_c), 
            .Q(\registers[8] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[0__666 .GSR = "DISABLED";
    FD1S3AX \registers_8[[31__667  (.D(\registers[8] [3]), .CK(clk_c), .Q(\registers[8] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[31__667 .GSR = "DISABLED";
    FD1S3AX \registers_8[[30__668  (.D(\registers[8] [2]), .CK(clk_c), .Q(\registers[8] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[30__668 .GSR = "DISABLED";
    FD1S3AX \registers_8[[29__669  (.D(\registers[8] [1]), .CK(clk_c), .Q(\registers[8] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[29__669 .GSR = "DISABLED";
    FD1S3AX \registers_8[[28__670  (.D(\registers[8] [0]), .CK(clk_c), .Q(\registers[8] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[28__670 .GSR = "DISABLED";
    FD1S3AX \registers_8[[27__671  (.D(\registers[8] [31]), .CK(clk_c), 
            .Q(\registers[8] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[27__671 .GSR = "DISABLED";
    FD1S3AX \registers_8[[26__672  (.D(\registers[8] [30]), .CK(clk_c), 
            .Q(\registers[8] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[26__672 .GSR = "DISABLED";
    FD1S3AX \registers_8[[25__673  (.D(\registers[8] [29]), .CK(clk_c), 
            .Q(\registers[8] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[25__673 .GSR = "DISABLED";
    FD1S3AX \registers_8[[24__674  (.D(\registers[8] [28]), .CK(clk_c), 
            .Q(\registers[8] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[24__674 .GSR = "DISABLED";
    FD1S3AX \registers_8[[23__675  (.D(\registers[8] [27]), .CK(clk_c), 
            .Q(\registers[8] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[23__675 .GSR = "DISABLED";
    FD1S3AX \registers_8[[22__676  (.D(\registers[8] [26]), .CK(clk_c), 
            .Q(\registers[8] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[22__676 .GSR = "DISABLED";
    FD1S3AX \registers_8[[21__677  (.D(\registers[8] [25]), .CK(clk_c), 
            .Q(\registers[8] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[21__677 .GSR = "DISABLED";
    FD1S3AX \registers_8[[20__678  (.D(\registers[8] [24]), .CK(clk_c), 
            .Q(\registers[8] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[20__678 .GSR = "DISABLED";
    FD1S3AX \registers_8[[19__679  (.D(\registers[8] [23]), .CK(clk_c), 
            .Q(\registers[8] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[19__679 .GSR = "DISABLED";
    FD1S3AX \registers_8[[18__680  (.D(\registers[8] [22]), .CK(clk_c), 
            .Q(\registers[8] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[18__680 .GSR = "DISABLED";
    FD1S3AX \registers_8[[17__681  (.D(\registers[8] [21]), .CK(clk_c), 
            .Q(\registers[8] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[17__681 .GSR = "DISABLED";
    FD1S3AX \registers_8[[16__682  (.D(\registers[8] [20]), .CK(clk_c), 
            .Q(\registers[8] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[16__682 .GSR = "DISABLED";
    FD1S3AX \registers_8[[15__683  (.D(\registers[8] [19]), .CK(clk_c), 
            .Q(\registers[8] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[15__683 .GSR = "DISABLED";
    FD1S3AX \registers_8[[14__684  (.D(\registers[8] [18]), .CK(clk_c), 
            .Q(\registers[8] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[14__684 .GSR = "DISABLED";
    FD1S3AX \registers_8[[13__685  (.D(\registers[8] [17]), .CK(clk_c), 
            .Q(\registers[8] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[13__685 .GSR = "DISABLED";
    FD1S3AX \registers_8[[12__686  (.D(\registers[8] [16]), .CK(clk_c), 
            .Q(\registers[8] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[12__686 .GSR = "DISABLED";
    FD1S3AX \registers_8[[11__687  (.D(\registers[8] [15]), .CK(clk_c), 
            .Q(\registers[8] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[11__687 .GSR = "DISABLED";
    FD1S3AX \registers_8[[10__688  (.D(\registers[8] [14]), .CK(clk_c), 
            .Q(\registers[8] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[10__688 .GSR = "DISABLED";
    FD1S3AX \registers_8[[9__689  (.D(\registers[8] [13]), .CK(clk_c), .Q(\registers[8] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[9__689 .GSR = "DISABLED";
    FD1S3AX \registers_8[[8__690  (.D(\registers[8] [12]), .CK(clk_c), .Q(\registers[8] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[8__690 .GSR = "DISABLED";
    FD1S3AX \registers_8[[7__691  (.D(\registers[8] [11]), .CK(clk_c), .Q(\registers[8] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[7__691 .GSR = "DISABLED";
    FD1S3AX \registers_8[[6__692  (.D(\registers[8] [10]), .CK(clk_c), .Q(\registers[8] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[6__692 .GSR = "DISABLED";
    FD1S3AX \registers_8[[5__693  (.D(\registers[8] [9]), .CK(clk_c), .Q(\registers[8] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[5__693 .GSR = "DISABLED";
    FD1S3AX \registers_8[[4__694  (.D(\registers[8] [8]), .CK(clk_c), .Q(\registers[8] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[4__694 .GSR = "DISABLED";
    FD1S3AX \registers_9[[3__695  (.D(registers_9__3__N_1789), .CK(clk_c), 
            .Q(\registers[9] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[3__695 .GSR = "DISABLED";
    FD1S3AX \registers_9[[2__696  (.D(registers_9__2__N_1792), .CK(clk_c), 
            .Q(\registers[9] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[2__696 .GSR = "DISABLED";
    FD1S3AX \registers_9[[1__697  (.D(registers_9__1__N_1793), .CK(clk_c), 
            .Q(\registers[9] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[1__697 .GSR = "DISABLED";
    FD1S3AX \registers_9[[0__698  (.D(registers_9__0__N_1794), .CK(clk_c), 
            .Q(\registers[9] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[0__698 .GSR = "DISABLED";
    FD1S3AX \registers_9[[31__699  (.D(\registers[9] [3]), .CK(clk_c), .Q(\registers[9] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[31__699 .GSR = "DISABLED";
    FD1S3AX \registers_9[[30__700  (.D(\registers[9] [2]), .CK(clk_c), .Q(\registers[9] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[30__700 .GSR = "DISABLED";
    FD1S3AX \registers_9[[29__701  (.D(\registers[9] [1]), .CK(clk_c), .Q(\registers[9] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[29__701 .GSR = "DISABLED";
    FD1S3AX \registers_9[[28__702  (.D(\registers[9] [0]), .CK(clk_c), .Q(\registers[9] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[28__702 .GSR = "DISABLED";
    FD1S3AX \registers_9[[27__703  (.D(\registers[9] [31]), .CK(clk_c), 
            .Q(\registers[9] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[27__703 .GSR = "DISABLED";
    FD1S3AX \registers_9[[26__704  (.D(\registers[9] [30]), .CK(clk_c), 
            .Q(\registers[9] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[26__704 .GSR = "DISABLED";
    FD1S3AX \registers_9[[25__705  (.D(\registers[9] [29]), .CK(clk_c), 
            .Q(\registers[9] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[25__705 .GSR = "DISABLED";
    FD1S3AX \registers_9[[24__706  (.D(\registers[9] [28]), .CK(clk_c), 
            .Q(\registers[9] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[24__706 .GSR = "DISABLED";
    FD1S3AX \registers_9[[23__707  (.D(\registers[9] [27]), .CK(clk_c), 
            .Q(\registers[9] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[23__707 .GSR = "DISABLED";
    FD1S3AX \registers_9[[22__708  (.D(\registers[9] [26]), .CK(clk_c), 
            .Q(\registers[9] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[22__708 .GSR = "DISABLED";
    FD1S3AX \registers_9[[21__709  (.D(\registers[9] [25]), .CK(clk_c), 
            .Q(\registers[9] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[21__709 .GSR = "DISABLED";
    FD1S3AX \registers_9[[20__710  (.D(\registers[9] [24]), .CK(clk_c), 
            .Q(\registers[9] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[20__710 .GSR = "DISABLED";
    FD1S3AX \registers_9[[19__711  (.D(\registers[9] [23]), .CK(clk_c), 
            .Q(\registers[9] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[19__711 .GSR = "DISABLED";
    FD1S3AX \registers_9[[18__712  (.D(\registers[9] [22]), .CK(clk_c), 
            .Q(\registers[9] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[18__712 .GSR = "DISABLED";
    FD1S3AX \registers_9[[17__713  (.D(\registers[9] [21]), .CK(clk_c), 
            .Q(\registers[9] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[17__713 .GSR = "DISABLED";
    FD1S3AX \registers_9[[16__714  (.D(\registers[9] [20]), .CK(clk_c), 
            .Q(\registers[9] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[16__714 .GSR = "DISABLED";
    FD1S3AX \registers_9[[15__715  (.D(\registers[9] [19]), .CK(clk_c), 
            .Q(\registers[9] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[15__715 .GSR = "DISABLED";
    FD1S3AX \registers_9[[14__716  (.D(\registers[9] [18]), .CK(clk_c), 
            .Q(\registers[9] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[14__716 .GSR = "DISABLED";
    FD1S3AX \registers_9[[13__717  (.D(\registers[9] [17]), .CK(clk_c), 
            .Q(\registers[9] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[13__717 .GSR = "DISABLED";
    FD1S3AX \registers_9[[12__718  (.D(\registers[9] [16]), .CK(clk_c), 
            .Q(\registers[9] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[12__718 .GSR = "DISABLED";
    FD1S3AX \registers_9[[11__719  (.D(\registers[9] [15]), .CK(clk_c), 
            .Q(\registers[9] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[11__719 .GSR = "DISABLED";
    FD1S3AX \registers_9[[10__720  (.D(\registers[9] [14]), .CK(clk_c), 
            .Q(\registers[9] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[10__720 .GSR = "DISABLED";
    FD1S3AX \registers_9[[9__721  (.D(\registers[9] [13]), .CK(clk_c), .Q(\registers[9] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[9__721 .GSR = "DISABLED";
    FD1S3AX \registers_9[[8__722  (.D(\registers[9] [12]), .CK(clk_c), .Q(\registers[9] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[8__722 .GSR = "DISABLED";
    FD1S3AX \registers_9[[7__723  (.D(\registers[9] [11]), .CK(clk_c), .Q(\registers[9] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[7__723 .GSR = "DISABLED";
    FD1S3AX \registers_9[[6__724  (.D(\registers[9] [10]), .CK(clk_c), .Q(\registers[9] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[6__724 .GSR = "DISABLED";
    FD1S3AX \registers_9[[5__725  (.D(\registers[9] [9]), .CK(clk_c), .Q(\registers[9] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[5__725 .GSR = "DISABLED";
    FD1S3AX \registers_9[[4__726  (.D(\registers[9] [8]), .CK(clk_c), .Q(\registers[9] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[4__726 .GSR = "DISABLED";
    FD1S3AX \registers_10[[3__727  (.D(registers_10__3__N_1795), .CK(clk_c), 
            .Q(\registers[10] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[3__727 .GSR = "DISABLED";
    FD1S3AX \registers_10[[2__728  (.D(registers_10__2__N_1798), .CK(clk_c), 
            .Q(\registers[10] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[2__728 .GSR = "DISABLED";
    FD1S3AX \registers_10[[1__729  (.D(registers_10__1__N_1799), .CK(clk_c), 
            .Q(\registers[10] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[1__729 .GSR = "DISABLED";
    FD1S3AX \registers_10[[0__730  (.D(registers_10__0__N_1800), .CK(clk_c), 
            .Q(\registers[10] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[0__730 .GSR = "DISABLED";
    FD1S3AX \registers_10[[31__731  (.D(\registers[10] [3]), .CK(clk_c), 
            .Q(\registers[10] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[31__731 .GSR = "DISABLED";
    FD1S3AX \registers_10[[30__732  (.D(\registers[10] [2]), .CK(clk_c), 
            .Q(\registers[10] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[30__732 .GSR = "DISABLED";
    FD1S3AX \registers_10[[29__733  (.D(\registers[10] [1]), .CK(clk_c), 
            .Q(\registers[10] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[29__733 .GSR = "DISABLED";
    FD1S3AX \registers_10[[28__734  (.D(\registers[10] [0]), .CK(clk_c), 
            .Q(\registers[10] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[28__734 .GSR = "DISABLED";
    FD1S3AX \registers_10[[27__735  (.D(\registers[10] [31]), .CK(clk_c), 
            .Q(\registers[10] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[27__735 .GSR = "DISABLED";
    FD1S3AX \registers_10[[26__736  (.D(\registers[10] [30]), .CK(clk_c), 
            .Q(\registers[10] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[26__736 .GSR = "DISABLED";
    FD1S3AX \registers_10[[25__737  (.D(\registers[10] [29]), .CK(clk_c), 
            .Q(\registers[10] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[25__737 .GSR = "DISABLED";
    FD1S3AX \registers_10[[24__738  (.D(\registers[10] [28]), .CK(clk_c), 
            .Q(\registers[10] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[24__738 .GSR = "DISABLED";
    FD1S3AX \registers_10[[23__739  (.D(\registers[10] [27]), .CK(clk_c), 
            .Q(\registers[10] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[23__739 .GSR = "DISABLED";
    FD1S3AX \registers_10[[22__740  (.D(\registers[10] [26]), .CK(clk_c), 
            .Q(\registers[10] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[22__740 .GSR = "DISABLED";
    FD1S3AX \registers_10[[21__741  (.D(\registers[10] [25]), .CK(clk_c), 
            .Q(\registers[10] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[21__741 .GSR = "DISABLED";
    FD1S3AX \registers_10[[20__742  (.D(\registers[10] [24]), .CK(clk_c), 
            .Q(\registers[10] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[20__742 .GSR = "DISABLED";
    FD1S3AX \registers_10[[19__743  (.D(\registers[10] [23]), .CK(clk_c), 
            .Q(\registers[10] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[19__743 .GSR = "DISABLED";
    FD1S3AX \registers_10[[18__744  (.D(\registers[10] [22]), .CK(clk_c), 
            .Q(\registers[10] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[18__744 .GSR = "DISABLED";
    FD1S3AX \registers_10[[17__745  (.D(\registers[10] [21]), .CK(clk_c), 
            .Q(\registers[10] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[17__745 .GSR = "DISABLED";
    FD1S3AX \registers_10[[16__746  (.D(\registers[10] [20]), .CK(clk_c), 
            .Q(\registers[10] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[16__746 .GSR = "DISABLED";
    FD1S3AX \registers_10[[15__747  (.D(\registers[10] [19]), .CK(clk_c), 
            .Q(\registers[10] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[15__747 .GSR = "DISABLED";
    FD1S3AX \registers_10[[14__748  (.D(\registers[10] [18]), .CK(clk_c), 
            .Q(\registers[10] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[14__748 .GSR = "DISABLED";
    FD1S3AX \registers_10[[13__749  (.D(\registers[10] [17]), .CK(clk_c), 
            .Q(\registers[10] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[13__749 .GSR = "DISABLED";
    FD1S3AX \registers_10[[12__750  (.D(\registers[10] [16]), .CK(clk_c), 
            .Q(\registers[10] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[12__750 .GSR = "DISABLED";
    FD1S3AX \registers_10[[11__751  (.D(\registers[10] [15]), .CK(clk_c), 
            .Q(\registers[10] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[11__751 .GSR = "DISABLED";
    FD1S3AX \registers_10[[10__752  (.D(\registers[10] [14]), .CK(clk_c), 
            .Q(\registers[10] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[10__752 .GSR = "DISABLED";
    FD1S3AX \registers_10[[9__753  (.D(\registers[10] [13]), .CK(clk_c), 
            .Q(\registers[10] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[9__753 .GSR = "DISABLED";
    FD1S3AX \registers_10[[8__754  (.D(\registers[10] [12]), .CK(clk_c), 
            .Q(\registers[10] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[8__754 .GSR = "DISABLED";
    FD1S3AX \registers_10[[7__755  (.D(\registers[10] [11]), .CK(clk_c), 
            .Q(\registers[10] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[7__755 .GSR = "DISABLED";
    FD1S3AX \registers_10[[6__756  (.D(\registers[10] [10]), .CK(clk_c), 
            .Q(\registers[10] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[6__756 .GSR = "DISABLED";
    FD1S3AX \registers_10[[5__757  (.D(\registers[10] [9]), .CK(clk_c), 
            .Q(\registers[10] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[5__757 .GSR = "DISABLED";
    FD1S3AX \registers_10[[4__758  (.D(\registers[10] [8]), .CK(clk_c), 
            .Q(\registers[10] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[4__758 .GSR = "DISABLED";
    FD1S3AX \registers_11[[3__759  (.D(registers_11__3__N_1801), .CK(clk_c), 
            .Q(\registers[11] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[3__759 .GSR = "DISABLED";
    FD1S3AX \registers_11[[2__760  (.D(registers_11__2__N_1804), .CK(clk_c), 
            .Q(\registers[11] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[2__760 .GSR = "DISABLED";
    FD1S3AX \registers_11[[1__761  (.D(registers_11__1__N_1805), .CK(clk_c), 
            .Q(\registers[11] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[1__761 .GSR = "DISABLED";
    FD1S3AX \registers_11[[0__762  (.D(registers_11__0__N_1806), .CK(clk_c), 
            .Q(\registers[11] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[0__762 .GSR = "DISABLED";
    FD1S3AX \registers_11[[31__763  (.D(\registers[11] [3]), .CK(clk_c), 
            .Q(\registers[11] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[31__763 .GSR = "DISABLED";
    FD1S3AX \registers_11[[30__764  (.D(\registers[11] [2]), .CK(clk_c), 
            .Q(\registers[11] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[30__764 .GSR = "DISABLED";
    FD1S3AX \registers_11[[29__765  (.D(\registers[11] [1]), .CK(clk_c), 
            .Q(\registers[11] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[29__765 .GSR = "DISABLED";
    FD1S3AX \registers_11[[28__766  (.D(\registers[11] [0]), .CK(clk_c), 
            .Q(\registers[11] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[28__766 .GSR = "DISABLED";
    FD1S3AX \registers_11[[27__767  (.D(\registers[11] [31]), .CK(clk_c), 
            .Q(\registers[11] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[27__767 .GSR = "DISABLED";
    FD1S3AX \registers_11[[26__768  (.D(\registers[11] [30]), .CK(clk_c), 
            .Q(\registers[11] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[26__768 .GSR = "DISABLED";
    FD1S3AX \registers_11[[25__769  (.D(\registers[11] [29]), .CK(clk_c), 
            .Q(\registers[11] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[25__769 .GSR = "DISABLED";
    FD1S3AX \registers_11[[24__770  (.D(\registers[11] [28]), .CK(clk_c), 
            .Q(\registers[11] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[24__770 .GSR = "DISABLED";
    FD1S3AX \registers_11[[23__771  (.D(\registers[11] [27]), .CK(clk_c), 
            .Q(\registers[11] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[23__771 .GSR = "DISABLED";
    FD1S3AX \registers_11[[22__772  (.D(\registers[11] [26]), .CK(clk_c), 
            .Q(\registers[11] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[22__772 .GSR = "DISABLED";
    FD1S3AX \registers_11[[21__773  (.D(\registers[11] [25]), .CK(clk_c), 
            .Q(\registers[11] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[21__773 .GSR = "DISABLED";
    FD1S3AX \registers_11[[20__774  (.D(\registers[11] [24]), .CK(clk_c), 
            .Q(\registers[11] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[20__774 .GSR = "DISABLED";
    FD1S3AX \registers_11[[19__775  (.D(\registers[11] [23]), .CK(clk_c), 
            .Q(\registers[11] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[19__775 .GSR = "DISABLED";
    FD1S3AX \registers_11[[18__776  (.D(\registers[11] [22]), .CK(clk_c), 
            .Q(\registers[11] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[18__776 .GSR = "DISABLED";
    FD1S3AX \registers_11[[17__777  (.D(\registers[11] [21]), .CK(clk_c), 
            .Q(\registers[11] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[17__777 .GSR = "DISABLED";
    FD1S3AX \registers_11[[16__778  (.D(\registers[11] [20]), .CK(clk_c), 
            .Q(\registers[11] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[16__778 .GSR = "DISABLED";
    FD1S3AX \registers_11[[15__779  (.D(\registers[11] [19]), .CK(clk_c), 
            .Q(\registers[11] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[15__779 .GSR = "DISABLED";
    FD1S3AX \registers_11[[14__780  (.D(\registers[11] [18]), .CK(clk_c), 
            .Q(\registers[11] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[14__780 .GSR = "DISABLED";
    FD1S3AX \registers_11[[13__781  (.D(\registers[11] [17]), .CK(clk_c), 
            .Q(\registers[11] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[13__781 .GSR = "DISABLED";
    FD1S3AX \registers_11[[12__782  (.D(\registers[11] [16]), .CK(clk_c), 
            .Q(\registers[11] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[12__782 .GSR = "DISABLED";
    FD1S3AX \registers_11[[11__783  (.D(\registers[11] [15]), .CK(clk_c), 
            .Q(\registers[11] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[11__783 .GSR = "DISABLED";
    FD1S3AX \registers_11[[10__784  (.D(\registers[11] [14]), .CK(clk_c), 
            .Q(\registers[11] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[10__784 .GSR = "DISABLED";
    FD1S3AX \registers_11[[9__785  (.D(\registers[11] [13]), .CK(clk_c), 
            .Q(\registers[11] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[9__785 .GSR = "DISABLED";
    FD1S3AX \registers_11[[8__786  (.D(\registers[11] [12]), .CK(clk_c), 
            .Q(\registers[11] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[8__786 .GSR = "DISABLED";
    FD1S3AX \registers_11[[7__787  (.D(\registers[11] [11]), .CK(clk_c), 
            .Q(\registers[11] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[7__787 .GSR = "DISABLED";
    FD1S3AX \registers_11[[6__788  (.D(\registers[11] [10]), .CK(clk_c), 
            .Q(\registers[11] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[6__788 .GSR = "DISABLED";
    FD1S3AX \registers_11[[5__789  (.D(\registers[11] [9]), .CK(clk_c), 
            .Q(\registers[11] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[5__789 .GSR = "DISABLED";
    FD1S3AX \registers_11[[4__790  (.D(\registers[11] [8]), .CK(clk_c), 
            .Q(\registers[11] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[4__790 .GSR = "DISABLED";
    FD1S3AX \registers_12[[3__791  (.D(registers_12__3__N_1807), .CK(clk_c), 
            .Q(\registers[12] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[3__791 .GSR = "DISABLED";
    FD1S3AX \registers_12[[2__792  (.D(registers_12__2__N_1810), .CK(clk_c), 
            .Q(\registers[12] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[2__792 .GSR = "DISABLED";
    FD1S3AX \registers_12[[1__793  (.D(registers_12__1__N_1811), .CK(clk_c), 
            .Q(\registers[12] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[1__793 .GSR = "DISABLED";
    FD1S3AX \registers_12[[0__794  (.D(registers_12__0__N_1812), .CK(clk_c), 
            .Q(\registers[12] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[0__794 .GSR = "DISABLED";
    FD1S3AX \registers_12[[31__795  (.D(\registers[12] [3]), .CK(clk_c), 
            .Q(\registers[12] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[31__795 .GSR = "DISABLED";
    FD1S3AX \registers_12[[30__796  (.D(\registers[12] [2]), .CK(clk_c), 
            .Q(\registers[12] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[30__796 .GSR = "DISABLED";
    FD1S3AX \registers_12[[29__797  (.D(\registers[12] [1]), .CK(clk_c), 
            .Q(\registers[12] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[29__797 .GSR = "DISABLED";
    FD1S3AX \registers_12[[28__798  (.D(\registers[12] [0]), .CK(clk_c), 
            .Q(\registers[12] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[28__798 .GSR = "DISABLED";
    FD1S3AX \registers_12[[27__799  (.D(\registers[12] [31]), .CK(clk_c), 
            .Q(\registers[12] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[27__799 .GSR = "DISABLED";
    FD1S3AX \registers_12[[26__800  (.D(\registers[12] [30]), .CK(clk_c), 
            .Q(\registers[12] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[26__800 .GSR = "DISABLED";
    FD1S3AX \registers_12[[25__801  (.D(\registers[12] [29]), .CK(clk_c), 
            .Q(\registers[12] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[25__801 .GSR = "DISABLED";
    FD1S3AX \registers_12[[24__802  (.D(\registers[12] [28]), .CK(clk_c), 
            .Q(\registers[12] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[24__802 .GSR = "DISABLED";
    FD1S3AX \registers_12[[23__803  (.D(\registers[12] [27]), .CK(clk_c), 
            .Q(\registers[12] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[23__803 .GSR = "DISABLED";
    FD1S3AX \registers_12[[22__804  (.D(\registers[12] [26]), .CK(clk_c), 
            .Q(\registers[12] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[22__804 .GSR = "DISABLED";
    FD1S3AX \registers_12[[21__805  (.D(\registers[12] [25]), .CK(clk_c), 
            .Q(\registers[12] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[21__805 .GSR = "DISABLED";
    FD1S3AX \registers_12[[20__806  (.D(\registers[12] [24]), .CK(clk_c), 
            .Q(\registers[12] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[20__806 .GSR = "DISABLED";
    FD1S3AX \registers_12[[19__807  (.D(\registers[12] [23]), .CK(clk_c), 
            .Q(\registers[12] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[19__807 .GSR = "DISABLED";
    FD1S3AX \registers_12[[18__808  (.D(\registers[12] [22]), .CK(clk_c), 
            .Q(\registers[12] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[18__808 .GSR = "DISABLED";
    FD1S3AX \registers_12[[17__809  (.D(\registers[12] [21]), .CK(clk_c), 
            .Q(\registers[12] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[17__809 .GSR = "DISABLED";
    FD1S3AX \registers_12[[16__810  (.D(\registers[12] [20]), .CK(clk_c), 
            .Q(\registers[12] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[16__810 .GSR = "DISABLED";
    FD1S3AX \registers_12[[15__811  (.D(\registers[12] [19]), .CK(clk_c), 
            .Q(\registers[12] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[15__811 .GSR = "DISABLED";
    FD1S3AX \registers_12[[14__812  (.D(\registers[12] [18]), .CK(clk_c), 
            .Q(\registers[12] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[14__812 .GSR = "DISABLED";
    FD1S3AX \registers_12[[13__813  (.D(\registers[12] [17]), .CK(clk_c), 
            .Q(\registers[12] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[13__813 .GSR = "DISABLED";
    FD1S3AX \registers_12[[12__814  (.D(\registers[12] [16]), .CK(clk_c), 
            .Q(\registers[12] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[12__814 .GSR = "DISABLED";
    FD1S3AX \registers_12[[11__815  (.D(\registers[12] [15]), .CK(clk_c), 
            .Q(\registers[12] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[11__815 .GSR = "DISABLED";
    FD1S3AX \registers_12[[10__816  (.D(\registers[12] [14]), .CK(clk_c), 
            .Q(\registers[12] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[10__816 .GSR = "DISABLED";
    FD1S3AX \registers_12[[9__817  (.D(\registers[12] [13]), .CK(clk_c), 
            .Q(\registers[12] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[9__817 .GSR = "DISABLED";
    FD1S3AX \registers_12[[8__818  (.D(\registers[12] [12]), .CK(clk_c), 
            .Q(\registers[12] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[8__818 .GSR = "DISABLED";
    FD1S3AX \registers_12[[7__819  (.D(\registers[12] [11]), .CK(clk_c), 
            .Q(\registers[12] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[7__819 .GSR = "DISABLED";
    FD1S3AX \registers_12[[6__820  (.D(\registers[12] [10]), .CK(clk_c), 
            .Q(\registers[12] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[6__820 .GSR = "DISABLED";
    FD1S3AX \registers_12[[5__821  (.D(\registers[12] [9]), .CK(clk_c), 
            .Q(\registers[12] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[5__821 .GSR = "DISABLED";
    FD1S3AX \registers_12[[4__822  (.D(\registers[12] [8]), .CK(clk_c), 
            .Q(\registers[12] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[4__822 .GSR = "DISABLED";
    FD1S3AX \registers_13[[3__823  (.D(registers_13__3__N_1813), .CK(clk_c), 
            .Q(\registers[13] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[3__823 .GSR = "DISABLED";
    FD1S3AX \registers_13[[2__824  (.D(registers_13__2__N_1816), .CK(clk_c), 
            .Q(\registers[13] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[2__824 .GSR = "DISABLED";
    FD1S3AX \registers_13[[1__825  (.D(registers_13__1__N_1817), .CK(clk_c), 
            .Q(\registers[13] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[1__825 .GSR = "DISABLED";
    FD1S3AX \registers_13[[0__826  (.D(registers_13__0__N_1818), .CK(clk_c), 
            .Q(\registers[13] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[0__826 .GSR = "DISABLED";
    FD1S3AX \registers_13[[31__827  (.D(\registers[13] [3]), .CK(clk_c), 
            .Q(\registers[13] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[31__827 .GSR = "DISABLED";
    FD1S3AX \registers_13[[30__828  (.D(\registers[13] [2]), .CK(clk_c), 
            .Q(\registers[13] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[30__828 .GSR = "DISABLED";
    FD1S3AX \registers_13[[29__829  (.D(\registers[13] [1]), .CK(clk_c), 
            .Q(\registers[13] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[29__829 .GSR = "DISABLED";
    FD1S3AX \registers_13[[28__830  (.D(\registers[13] [0]), .CK(clk_c), 
            .Q(\registers[13] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[28__830 .GSR = "DISABLED";
    FD1S3AX \registers_13[[27__831  (.D(\registers[13] [31]), .CK(clk_c), 
            .Q(\registers[13] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[27__831 .GSR = "DISABLED";
    FD1S3AX \registers_13[[26__832  (.D(\registers[13] [30]), .CK(clk_c), 
            .Q(\registers[13] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[26__832 .GSR = "DISABLED";
    FD1S3AX \registers_13[[25__833  (.D(\registers[13] [29]), .CK(clk_c), 
            .Q(\registers[13] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[25__833 .GSR = "DISABLED";
    FD1S3AX \registers_13[[24__834  (.D(\registers[13] [28]), .CK(clk_c), 
            .Q(\registers[13] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[24__834 .GSR = "DISABLED";
    FD1S3AX \registers_13[[23__835  (.D(\registers[13] [27]), .CK(clk_c), 
            .Q(\registers[13] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[23__835 .GSR = "DISABLED";
    FD1S3AX \registers_13[[22__836  (.D(\registers[13] [26]), .CK(clk_c), 
            .Q(\registers[13] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[22__836 .GSR = "DISABLED";
    FD1S3AX \registers_13[[21__837  (.D(\registers[13] [25]), .CK(clk_c), 
            .Q(\registers[13] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[21__837 .GSR = "DISABLED";
    FD1S3AX \registers_13[[20__838  (.D(\registers[13] [24]), .CK(clk_c), 
            .Q(\registers[13] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[20__838 .GSR = "DISABLED";
    FD1S3AX \registers_13[[19__839  (.D(\registers[13] [23]), .CK(clk_c), 
            .Q(\registers[13] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[19__839 .GSR = "DISABLED";
    FD1S3AX \registers_13[[18__840  (.D(\registers[13] [22]), .CK(clk_c), 
            .Q(\registers[13] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[18__840 .GSR = "DISABLED";
    FD1S3AX \registers_13[[17__841  (.D(\registers[13] [21]), .CK(clk_c), 
            .Q(\registers[13] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[17__841 .GSR = "DISABLED";
    FD1S3AX \registers_13[[16__842  (.D(\registers[13] [20]), .CK(clk_c), 
            .Q(\registers[13] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[16__842 .GSR = "DISABLED";
    FD1S3AX \registers_13[[15__843  (.D(\registers[13] [19]), .CK(clk_c), 
            .Q(\registers[13] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[15__843 .GSR = "DISABLED";
    FD1S3AX \registers_13[[14__844  (.D(\registers[13] [18]), .CK(clk_c), 
            .Q(\registers[13] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[14__844 .GSR = "DISABLED";
    FD1S3AX \registers_13[[13__845  (.D(\registers[13] [17]), .CK(clk_c), 
            .Q(\registers[13] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[13__845 .GSR = "DISABLED";
    FD1S3AX \registers_13[[12__846  (.D(\registers[13] [16]), .CK(clk_c), 
            .Q(\registers[13] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[12__846 .GSR = "DISABLED";
    FD1S3AX \registers_13[[11__847  (.D(\registers[13] [15]), .CK(clk_c), 
            .Q(\registers[13] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[11__847 .GSR = "DISABLED";
    FD1S3AX \registers_13[[10__848  (.D(\registers[13] [14]), .CK(clk_c), 
            .Q(\registers[13] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[10__848 .GSR = "DISABLED";
    FD1S3AX \registers_13[[9__849  (.D(\registers[13] [13]), .CK(clk_c), 
            .Q(\registers[13] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[9__849 .GSR = "DISABLED";
    FD1S3AX \registers_13[[8__850  (.D(\registers[13] [12]), .CK(clk_c), 
            .Q(\registers[13] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[8__850 .GSR = "DISABLED";
    FD1S3AX \registers_13[[7__851  (.D(\registers[13] [11]), .CK(clk_c), 
            .Q(\registers[13] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[7__851 .GSR = "DISABLED";
    FD1S3AX \registers_13[[6__852  (.D(\registers[13] [10]), .CK(clk_c), 
            .Q(\registers[13] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[6__852 .GSR = "DISABLED";
    FD1S3AX \registers_13[[5__853  (.D(\registers[13] [9]), .CK(clk_c), 
            .Q(\registers[13] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[5__853 .GSR = "DISABLED";
    FD1S3AX \registers_13[[4__854  (.D(\registers[13] [8]), .CK(clk_c), 
            .Q(\registers[13] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[4__854 .GSR = "DISABLED";
    FD1S3AX \registers_14[[3__855  (.D(registers_14__3__N_1819), .CK(clk_c), 
            .Q(\registers[14] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[3__855 .GSR = "DISABLED";
    FD1S3AX \registers_14[[2__856  (.D(registers_14__2__N_1822), .CK(clk_c), 
            .Q(\registers[14] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[2__856 .GSR = "DISABLED";
    FD1S3AX \registers_14[[1__857  (.D(registers_14__1__N_1823), .CK(clk_c), 
            .Q(\registers[14] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[1__857 .GSR = "DISABLED";
    FD1S3AX \registers_14[[0__858  (.D(registers_14__0__N_1824), .CK(clk_c), 
            .Q(\registers[14] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[0__858 .GSR = "DISABLED";
    FD1S3AX \registers_14[[31__859  (.D(\registers[14] [3]), .CK(clk_c), 
            .Q(\registers[14] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[31__859 .GSR = "DISABLED";
    FD1S3AX \registers_14[[30__860  (.D(\registers[14] [2]), .CK(clk_c), 
            .Q(\registers[14] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[30__860 .GSR = "DISABLED";
    FD1S3AX \registers_14[[29__861  (.D(\registers[14] [1]), .CK(clk_c), 
            .Q(\registers[14] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[29__861 .GSR = "DISABLED";
    FD1S3AX \registers_14[[28__862  (.D(\registers[14] [0]), .CK(clk_c), 
            .Q(\registers[14] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[28__862 .GSR = "DISABLED";
    FD1S3AX \registers_14[[27__863  (.D(\registers[14] [31]), .CK(clk_c), 
            .Q(\registers[14] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[27__863 .GSR = "DISABLED";
    FD1S3AX \registers_14[[26__864  (.D(\registers[14] [30]), .CK(clk_c), 
            .Q(\registers[14] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[26__864 .GSR = "DISABLED";
    FD1S3AX \registers_14[[25__865  (.D(\registers[14] [29]), .CK(clk_c), 
            .Q(\registers[14] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[25__865 .GSR = "DISABLED";
    FD1S3AX \registers_14[[24__866  (.D(\registers[14] [28]), .CK(clk_c), 
            .Q(\registers[14] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[24__866 .GSR = "DISABLED";
    FD1S3AX \registers_14[[23__867  (.D(\registers[14] [27]), .CK(clk_c), 
            .Q(\registers[14] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[23__867 .GSR = "DISABLED";
    FD1S3AX \registers_14[[22__868  (.D(\registers[14] [26]), .CK(clk_c), 
            .Q(\registers[14] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[22__868 .GSR = "DISABLED";
    FD1S3AX \registers_14[[21__869  (.D(\registers[14] [25]), .CK(clk_c), 
            .Q(\registers[14] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[21__869 .GSR = "DISABLED";
    FD1S3AX \registers_14[[20__870  (.D(\registers[14] [24]), .CK(clk_c), 
            .Q(\registers[14] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[20__870 .GSR = "DISABLED";
    FD1S3AX \registers_14[[19__871  (.D(\registers[14] [23]), .CK(clk_c), 
            .Q(\registers[14] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[19__871 .GSR = "DISABLED";
    FD1S3AX \registers_14[[18__872  (.D(\registers[14] [22]), .CK(clk_c), 
            .Q(\registers[14] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[18__872 .GSR = "DISABLED";
    FD1S3AX \registers_14[[17__873  (.D(\registers[14] [21]), .CK(clk_c), 
            .Q(\registers[14] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[17__873 .GSR = "DISABLED";
    FD1S3AX \registers_14[[16__874  (.D(\registers[14] [20]), .CK(clk_c), 
            .Q(\registers[14] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[16__874 .GSR = "DISABLED";
    FD1S3AX \registers_14[[15__875  (.D(\registers[14] [19]), .CK(clk_c), 
            .Q(\registers[14] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[15__875 .GSR = "DISABLED";
    FD1S3AX \registers_14[[14__876  (.D(\registers[14] [18]), .CK(clk_c), 
            .Q(\registers[14] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[14__876 .GSR = "DISABLED";
    FD1S3AX \registers_14[[13__877  (.D(\registers[14] [17]), .CK(clk_c), 
            .Q(\registers[14] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[13__877 .GSR = "DISABLED";
    FD1S3AX \registers_14[[12__878  (.D(\registers[14] [16]), .CK(clk_c), 
            .Q(\registers[14] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[12__878 .GSR = "DISABLED";
    FD1S3AX \registers_14[[11__879  (.D(\registers[14] [15]), .CK(clk_c), 
            .Q(\registers[14] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[11__879 .GSR = "DISABLED";
    FD1S3AX \registers_14[[10__880  (.D(\registers[14] [14]), .CK(clk_c), 
            .Q(\registers[14] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[10__880 .GSR = "DISABLED";
    FD1S3AX \registers_14[[9__881  (.D(\registers[14] [13]), .CK(clk_c), 
            .Q(\registers[14] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[9__881 .GSR = "DISABLED";
    FD1S3AX \registers_14[[8__882  (.D(\registers[14] [12]), .CK(clk_c), 
            .Q(\registers[14] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[8__882 .GSR = "DISABLED";
    FD1S3AX \registers_14[[7__883  (.D(\registers[14] [11]), .CK(clk_c), 
            .Q(\registers[14] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[7__883 .GSR = "DISABLED";
    FD1S3AX \registers_14[[6__884  (.D(\registers[14] [10]), .CK(clk_c), 
            .Q(\registers[14] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[6__884 .GSR = "DISABLED";
    FD1S3AX \registers_14[[5__885  (.D(\registers[14] [9]), .CK(clk_c), 
            .Q(\registers[14] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[5__885 .GSR = "DISABLED";
    FD1S3AX \registers_14[[4__886  (.D(\registers[14] [8]), .CK(clk_c), 
            .Q(\registers[14] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[4__886 .GSR = "DISABLED";
    FD1S3AX \registers_15[[3__887  (.D(registers_15__3__N_1825), .CK(clk_c), 
            .Q(\registers[15] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[3__887 .GSR = "DISABLED";
    FD1S3AX \registers_15[[2__888  (.D(registers_15__2__N_1828), .CK(clk_c), 
            .Q(\registers[15] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[2__888 .GSR = "DISABLED";
    FD1S3AX \registers_15[[1__889  (.D(registers_15__1__N_1829), .CK(clk_c), 
            .Q(\registers[15] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[1__889 .GSR = "DISABLED";
    FD1S3AX \registers_15[[0__890  (.D(registers_15__0__N_1830), .CK(clk_c), 
            .Q(\registers[15] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[0__890 .GSR = "DISABLED";
    FD1S3AX \registers_15[[31__891  (.D(\registers[15] [3]), .CK(clk_c), 
            .Q(\registers[15] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[31__891 .GSR = "DISABLED";
    FD1S3AX \registers_15[[30__892  (.D(\registers[15] [2]), .CK(clk_c), 
            .Q(\registers[15] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[30__892 .GSR = "DISABLED";
    FD1S3AX \registers_15[[29__893  (.D(\registers[15] [1]), .CK(clk_c), 
            .Q(\registers[15] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[29__893 .GSR = "DISABLED";
    FD1S3AX \registers_15[[28__894  (.D(\registers[15] [0]), .CK(clk_c), 
            .Q(\registers[15] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[28__894 .GSR = "DISABLED";
    FD1S3AX \registers_15[[27__895  (.D(\registers[15] [31]), .CK(clk_c), 
            .Q(\registers[15] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[27__895 .GSR = "DISABLED";
    FD1S3AX \registers_15[[26__896  (.D(\registers[15] [30]), .CK(clk_c), 
            .Q(\registers[15] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[26__896 .GSR = "DISABLED";
    FD1S3AX \registers_15[[25__897  (.D(\registers[15] [29]), .CK(clk_c), 
            .Q(\registers[15] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[25__897 .GSR = "DISABLED";
    FD1S3AX \registers_15[[24__898  (.D(\registers[15] [28]), .CK(clk_c), 
            .Q(\registers[15] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[24__898 .GSR = "DISABLED";
    FD1S3AX \registers_15[[23__899  (.D(\registers[15] [27]), .CK(clk_c), 
            .Q(\registers[15] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[23__899 .GSR = "DISABLED";
    FD1S3AX \registers_15[[22__900  (.D(\registers[15] [26]), .CK(clk_c), 
            .Q(\registers[15] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[22__900 .GSR = "DISABLED";
    FD1S3AX \registers_15[[21__901  (.D(\registers[15] [25]), .CK(clk_c), 
            .Q(\registers[15] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[21__901 .GSR = "DISABLED";
    FD1S3AX \registers_15[[20__902  (.D(\registers[15] [24]), .CK(clk_c), 
            .Q(\registers[15] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[20__902 .GSR = "DISABLED";
    FD1S3AX \registers_15[[19__903  (.D(\registers[15] [23]), .CK(clk_c), 
            .Q(\registers[15] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[19__903 .GSR = "DISABLED";
    FD1S3AX \registers_15[[18__904  (.D(\registers[15] [22]), .CK(clk_c), 
            .Q(\registers[15] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[18__904 .GSR = "DISABLED";
    FD1S3AX \registers_15[[17__905  (.D(\registers[15] [21]), .CK(clk_c), 
            .Q(\registers[15] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[17__905 .GSR = "DISABLED";
    FD1S3AX \registers_15[[16__906  (.D(\registers[15] [20]), .CK(clk_c), 
            .Q(\registers[15] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[16__906 .GSR = "DISABLED";
    FD1S3AX \registers_15[[15__907  (.D(\registers[15] [19]), .CK(clk_c), 
            .Q(\registers[15] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[15__907 .GSR = "DISABLED";
    FD1S3AX \registers_15[[14__908  (.D(\registers[15] [18]), .CK(clk_c), 
            .Q(\registers[15] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[14__908 .GSR = "DISABLED";
    FD1S3AX \registers_15[[13__909  (.D(\registers[15] [17]), .CK(clk_c), 
            .Q(\registers[15] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[13__909 .GSR = "DISABLED";
    FD1S3AX \registers_15[[12__910  (.D(\registers[15] [16]), .CK(clk_c), 
            .Q(\registers[15] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[12__910 .GSR = "DISABLED";
    FD1S3AX \registers_15[[11__911  (.D(\registers[15] [15]), .CK(clk_c), 
            .Q(\registers[15] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[11__911 .GSR = "DISABLED";
    FD1S3AX \registers_15[[10__912  (.D(\registers[15] [14]), .CK(clk_c), 
            .Q(\registers[15] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[10__912 .GSR = "DISABLED";
    FD1S3AX \registers_15[[9__913  (.D(\registers[15] [13]), .CK(clk_c), 
            .Q(\registers[15] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[9__913 .GSR = "DISABLED";
    FD1S3AX \registers_15[[8__914  (.D(\registers[15] [12]), .CK(clk_c), 
            .Q(\registers[15] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[8__914 .GSR = "DISABLED";
    FD1S3AX \registers_15[[7__915  (.D(\registers[15] [11]), .CK(clk_c), 
            .Q(\registers[15] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[7__915 .GSR = "DISABLED";
    FD1S3AX \registers_15[[6__916  (.D(\registers[15] [10]), .CK(clk_c), 
            .Q(\registers[15] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[6__916 .GSR = "DISABLED";
    FD1S3AX \registers_15[[5__917  (.D(\registers[15] [9]), .CK(clk_c), 
            .Q(\registers[15] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[5__917 .GSR = "DISABLED";
    FD1S3AX \registers_15[[4__918  (.D(\registers[15] [8]), .CK(clk_c), 
            .Q(\registers[15] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[4__918 .GSR = "DISABLED";
    FD1S3AX \registers_1[[3__503  (.D(registers_1__3__N_1753), .CK(clk_c), 
            .Q(\registers[1] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[3__503 .GSR = "DISABLED";
    LUT4 i22824_3_lut (.A(\registers[14] [6]), .B(\registers[15] [6]), .C(rs2[0]), 
         .Z(n25167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22824_3_lut.init = 16'hcaca;
    LUT4 i22823_3_lut (.A(\registers[12] [6]), .B(\registers[13] [6]), .C(rs2[0]), 
         .Z(n25166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22823_3_lut.init = 16'hcaca;
    LUT4 i22822_3_lut (.A(\registers[10] [6]), .B(\registers[11] [6]), .C(rs2[0]), 
         .Z(n25165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22822_3_lut.init = 16'hcaca;
    LUT4 i22821_3_lut (.A(\registers[8] [6]), .B(\registers[9] [6]), .C(rs2[0]), 
         .Z(n25164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22821_3_lut.init = 16'hcaca;
    LUT4 i22820_3_lut (.A(\registers[6] [6]), .B(\registers[7] [6]), .C(rs2[0]), 
         .Z(n25163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22820_3_lut.init = 16'hcaca;
    LUT4 i22819_3_lut (.A(\registers[5] [6]), .B(rs2[0]), .Z(n25162)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22819_3_lut.init = 16'h8888;
    LUT4 rs1_3__I_0_Mux_1_i12_3_lut (.A(\registers[14] [5]), .B(\registers[15] [5]), 
         .C(rs1[0]), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i12_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i11_3_lut (.A(\registers[12] [5]), .B(\registers[13] [5]), 
         .C(rs1[0]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i11_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i9_3_lut (.A(\registers[10] [5]), .B(\registers[11] [5]), 
         .C(rs1[0]), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i8_3_lut (.A(\registers[8] [5]), .B(\registers[9] [5]), 
         .C(rs1[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i8_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i5_3_lut (.A(\registers[6] [7]), .B(\registers[7] [7]), 
         .C(rs2[0]), .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i5_3_lut (.A(\registers[6] [5]), .B(\registers[7] [5]), 
         .C(rs1[0]), .Z(n5_adj_2600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i12_3_lut (.A(\registers[14] [5]), .B(\registers[15] [5]), 
         .C(rs2[0]), .Z(n12_adj_2601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i12_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i11_3_lut (.A(\registers[12] [5]), .B(\registers[13] [5]), 
         .C(rs2[0]), .Z(n11_adj_2602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i11_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i9_3_lut (.A(\registers[10] [5]), .B(\registers[11] [5]), 
         .C(rs2[0]), .Z(n9_adj_2603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i8_3_lut (.A(\registers[8] [5]), .B(\registers[9] [5]), 
         .C(rs2[0]), .Z(n8_adj_2604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i8_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i5_3_lut (.A(\registers[6] [5]), .B(\registers[7] [5]), 
         .C(rs2[0]), .Z(n5_adj_2605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 registers_15__7__I_0_3_lut_4_lut (.A(n27315), .B(n27116), .C(debug_rd[3]), 
         .D(\registers[15] [7]), .Z(registers_15__3__N_1825)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 rs2_3__I_0_Mux_3_i4_3_lut (.A(\reg_access[4][3] ), .B(\registers[5] [7]), 
         .C(rs2[0]), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i4_3_lut.init = 16'hcaca;
    LUT4 registers_15__6__I_0_3_lut_4_lut (.A(n27315), .B(n27116), .C(debug_rd[2]), 
         .D(\registers[15] [6]), .Z(registers_15__2__N_1828)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i23104_3_lut (.A(n4), .B(n5), .C(rs2[1]), .Z(n25315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23104_3_lut.init = 16'hcaca;
    LUT4 registers_15__5__I_0_3_lut_4_lut (.A(n27315), .B(n27116), .C(debug_rd[1]), 
         .D(\registers[15] [5]), .Z(registers_15__1__N_1829)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_15__4__I_0_3_lut_4_lut (.A(n27315), .B(n27116), .C(debug_rd[0]), 
         .D(\registers[15] [4]), .Z(registers_15__0__N_1830)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__7__I_0_3_lut_4_lut (.A(n27315), .B(n27117), .C(debug_rd[3]), 
         .D(\registers[14] [7]), .Z(registers_14__3__N_1819)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__6__I_0_3_lut_4_lut (.A(n27315), .B(n27117), .C(debug_rd[2]), 
         .D(\registers[14] [6]), .Z(registers_14__2__N_1822)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__5__I_0_3_lut_4_lut (.A(n27315), .B(n27117), .C(debug_rd[1]), 
         .D(\registers[14] [5]), .Z(registers_14__1__N_1823)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__4__I_0_3_lut_4_lut (.A(n27315), .B(n27117), .C(debug_rd[0]), 
         .D(\registers[14] [4]), .Z(registers_14__0__N_1824)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__7__I_0_3_lut_4_lut (.A(n27315), .B(n27118), .C(debug_rd[3]), 
         .D(\registers[13] [7]), .Z(registers_13__3__N_1813)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__6__I_0_3_lut_4_lut (.A(n27315), .B(n27118), .C(debug_rd[2]), 
         .D(\registers[13] [6]), .Z(registers_13__2__N_1816)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 rs1_3__I_0_Mux_3_i5_3_lut (.A(\registers[6] [7]), .B(\registers[7] [7]), 
         .C(rs1[0]), .Z(n5_adj_2606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 i22970_3_lut (.A(n25311), .B(n25312), .C(rs1[3]), .Z(data_rs1[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22970_3_lut.init = 16'hcaca;
    LUT4 registers_13__5__I_0_3_lut_4_lut (.A(n27315), .B(n27118), .C(debug_rd[1]), 
         .D(\registers[13] [5]), .Z(registers_13__1__N_1817)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__4__I_0_3_lut_4_lut (.A(n27315), .B(n27118), .C(debug_rd[0]), 
         .D(\registers[13] [4]), .Z(registers_13__0__N_1818)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__5__I_0_3_lut_4_lut (.A(n27315), .B(n27115), .C(debug_rd[1]), 
         .D(\registers[12] [5]), .Z(registers_12__1__N_1811)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__6__I_0_3_lut_4_lut (.A(n27315), .B(n27115), .C(debug_rd[2]), 
         .D(\registers[12] [6]), .Z(registers_12__2__N_1810)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__7__I_0_3_lut_4_lut (.A(n27315), .B(n27115), .C(debug_rd[3]), 
         .D(\registers[12] [7]), .Z(registers_12__3__N_1807)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__4__I_0_3_lut_4_lut (.A(n27315), .B(n27115), .C(debug_rd[0]), 
         .D(\registers[12] [4]), .Z(registers_12__0__N_1812)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_11__7__I_0_3_lut_4_lut (.A(n27316), .B(n27116), .C(debug_rd[3]), 
         .D(\registers[11] [7]), .Z(registers_11__3__N_1801)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs1_3__I_0_Mux_3_i4_3_lut (.A(\reg_access[4][3] ), .B(\registers[5] [7]), 
         .C(rs1[0]), .Z(n4_adj_2607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i4_3_lut.init = 16'hcaca;
    LUT4 registers_11__6__I_0_3_lut_4_lut (.A(n27316), .B(n27116), .C(debug_rd[2]), 
         .D(\registers[11] [6]), .Z(registers_11__2__N_1804)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__5__I_0_3_lut_4_lut (.A(n27316), .B(n27116), .C(debug_rd[1]), 
         .D(\registers[11] [5]), .Z(registers_11__1__N_1805)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__4__I_0_3_lut_4_lut (.A(n27316), .B(n27116), .C(debug_rd[0]), 
         .D(\registers[11] [4]), .Z(registers_11__0__N_1806)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__7__I_0_3_lut_4_lut (.A(n27316), .B(n27117), .C(debug_rd[3]), 
         .D(\registers[10] [7]), .Z(registers_10__3__N_1795)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 i23106_3_lut (.A(n4_adj_2607), .B(n5_adj_2606), .C(rs1[1]), .Z(n25308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23106_3_lut.init = 16'hcaca;
    LUT4 registers_10__6__I_0_3_lut_4_lut (.A(n27316), .B(n27117), .C(debug_rd[2]), 
         .D(\registers[10] [6]), .Z(registers_10__2__N_1798)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__5__I_0_3_lut_4_lut (.A(n27316), .B(n27117), .C(debug_rd[1]), 
         .D(\registers[10] [5]), .Z(registers_10__1__N_1799)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__4__I_0_3_lut_4_lut (.A(n27316), .B(n27117), .C(debug_rd[0]), 
         .D(\registers[10] [4]), .Z(registers_10__0__N_1800)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__7__I_0_3_lut_4_lut (.A(n27316), .B(n27118), .C(debug_rd[3]), 
         .D(\registers[9] [7]), .Z(registers_9__3__N_1789)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__6__I_0_3_lut_4_lut (.A(n27316), .B(n27118), .C(debug_rd[2]), 
         .D(\registers[9] [6]), .Z(registers_9__2__N_1792)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__5__I_0_3_lut_4_lut (.A(n27316), .B(n27118), .C(debug_rd[1]), 
         .D(\registers[9] [5]), .Z(registers_9__1__N_1793)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__4__I_0_3_lut_4_lut (.A(n27316), .B(n27118), .C(debug_rd[0]), 
         .D(\registers[9] [4]), .Z(registers_9__0__N_1794)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs2_3__I_0_Mux_3_i12_3_lut (.A(\registers[14] [7]), .B(\registers[15] [7]), 
         .C(rs2[0]), .Z(n12_adj_2608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i12_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i11_3_lut (.A(\registers[12] [7]), .B(\registers[13] [7]), 
         .C(rs2[0]), .Z(n11_adj_2609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i9_3_lut (.A(\registers[10] [7]), .B(\registers[11] [7]), 
         .C(rs2[0]), .Z(n9_adj_2610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i8_3_lut (.A(\registers[8] [7]), .B(\registers[9] [7]), 
         .C(rs2[0]), .Z(n8_adj_2611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i12_3_lut (.A(\registers[14] [7]), .B(\registers[15] [7]), 
         .C(rs1[0]), .Z(n12_adj_2612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i12_3_lut.init = 16'hcaca;
    LUT4 registers_8__7__I_0_3_lut_4_lut (.A(n27316), .B(n27115), .C(debug_rd[3]), 
         .D(\registers[8] [7]), .Z(registers_8__3__N_1783)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__6__I_0_3_lut_4_lut (.A(n27316), .B(n27115), .C(debug_rd[2]), 
         .D(\registers[8] [6]), .Z(registers_8__2__N_1786)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__5__I_0_3_lut_4_lut (.A(n27316), .B(n27115), .C(debug_rd[1]), 
         .D(\registers[8] [5]), .Z(registers_8__1__N_1787)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__4__I_0_3_lut_4_lut (.A(n27316), .B(n27115), .C(debug_rd[0]), 
         .D(\registers[8] [4]), .Z(registers_8__0__N_1788)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__7__I_0_3_lut_4_lut (.A(n27317), .B(n27116), .C(debug_rd[3]), 
         .D(\registers[7] [7]), .Z(registers_7__3__N_1777)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__6__I_0_3_lut_4_lut (.A(n27317), .B(n27116), .C(debug_rd[2]), 
         .D(\registers[7] [6]), .Z(registers_7__2__N_1780)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__5__I_0_3_lut_4_lut (.A(n27317), .B(n27116), .C(debug_rd[1]), 
         .D(\registers[7] [5]), .Z(registers_7__1__N_1781)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__4__I_0_3_lut_4_lut (.A(n27317), .B(n27116), .C(debug_rd[0]), 
         .D(\registers[7] [4]), .Z(registers_7__0__N_1782)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__7__I_0_3_lut_4_lut (.A(n27317), .B(n27117), .C(debug_rd[3]), 
         .D(\registers[6] [7]), .Z(registers_6__3__N_1771)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__6__I_0_3_lut_4_lut (.A(n27317), .B(n27117), .C(debug_rd[2]), 
         .D(\registers[6] [6]), .Z(registers_6__2__N_1774)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__5__I_0_3_lut_4_lut (.A(n27317), .B(n27117), .C(debug_rd[1]), 
         .D(\registers[6] [5]), .Z(registers_6__1__N_1775)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__4__I_0_3_lut_4_lut (.A(n27317), .B(n27117), .C(debug_rd[0]), 
         .D(\registers[6] [4]), .Z(registers_6__0__N_1776)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs1_3__I_0_Mux_3_i11_3_lut (.A(\registers[12] [7]), .B(\registers[13] [7]), 
         .C(rs1[0]), .Z(n11_adj_2613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 registers_5__6__I_0_3_lut_4_lut (.A(n27317), .B(n27118), .C(debug_rd[2]), 
         .D(\registers[5] [6]), .Z(registers_5__2__N_1768)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs1_3__I_0_Mux_3_i9_3_lut (.A(\registers[10] [7]), .B(\registers[11] [7]), 
         .C(rs1[0]), .Z(n9_adj_2614)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i8_3_lut (.A(\registers[8] [7]), .B(\registers[9] [7]), 
         .C(rs1[0]), .Z(n8_adj_2615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 registers_5__4__I_0_3_lut_4_lut (.A(n27317), .B(n27118), .C(debug_rd[0]), 
         .D(\registers[5] [4]), .Z(registers_5__0__N_1770)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__4__I_0_3_lut_4_lut.init = 16'hfb40;
    PFUMX i22905 (.BLUT(n25240), .ALUT(n25241), .C0(rs1[1]), .Z(n25248));
    LUT4 registers_5__5__I_0_3_lut_4_lut (.A(n27317), .B(n27118), .C(debug_rd[1]), 
         .D(\registers[5] [5]), .Z(registers_5__1__N_1769)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__7__I_0_3_lut_4_lut (.A(n27317), .B(n27118), .C(debug_rd[3]), 
         .D(\registers[5] [7]), .Z(registers_5__3__N_1765)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_2__6__I_0_3_lut_4_lut (.A(n27117), .B(n27318), .C(debug_rd[2]), 
         .D(\registers[2] [6]), .Z(registers_2__2__N_1762)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__4__I_0_3_lut_4_lut (.A(n27117), .B(n27318), .C(debug_rd[0]), 
         .D(\registers[2] [4]), .Z(registers_2__0__N_1764)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__4__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__5__I_0_3_lut_4_lut (.A(n27117), .B(n27318), .C(debug_rd[1]), 
         .D(\registers[2] [5]), .Z(registers_2__1__N_1763)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__7__I_0_3_lut_4_lut (.A(n27117), .B(n27318), .C(debug_rd[3]), 
         .D(\registers[2] [7]), .Z(registers_2__3__N_1759)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__7__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__5__I_0_3_lut_4_lut (.A(n27118), .B(n27318), .C(debug_rd[1]), 
         .D(\registers[1] [5]), .Z(registers_1__1__N_1757)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__7__I_0_3_lut_4_lut (.A(n27118), .B(n27318), .C(debug_rd[3]), 
         .D(\registers[1] [7]), .Z(registers_1__3__N_1753)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__7__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__4__I_0_3_lut_4_lut (.A(n27118), .B(n27318), .C(debug_rd[0]), 
         .D(\registers[1] [4]), .Z(registers_1__0__N_1758)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__4__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__6__I_0_3_lut_4_lut (.A(n27118), .B(n27318), .C(debug_rd[2]), 
         .D(\registers[1] [6]), .Z(registers_1__2__N_1756)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 i12295_2_lut_rep_690 (.A(rd[2]), .B(rd[3]), .Z(n27315)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12295_2_lut_rep_690.init = 16'h8888;
    LUT4 i22889_3_lut (.A(n25230), .B(n25231), .C(rs1[3]), .Z(data_rs1[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22889_3_lut.init = 16'hcaca;
    LUT4 equal_139_i6_2_lut_rep_691 (.A(rd[2]), .B(rd[3]), .Z(n27316)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam equal_139_i6_2_lut_rep_691.init = 16'hbbbb;
    LUT4 equal_135_i6_2_lut_rep_692 (.A(rd[2]), .B(rd[3]), .Z(n27317)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam equal_135_i6_2_lut_rep_692.init = 16'hdddd;
    LUT4 i12640_2_lut_rep_693 (.A(rd[3]), .B(rd[2]), .Z(n27318)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12640_2_lut_rep_693.init = 16'heeee;
    LUT4 i23543_3_lut (.A(n28571), .B(n28573), .C(\counter_hi[2] ), .Z(\reg_access[4][3] )) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(40[41:55])
    defparam i23543_3_lut.init = 16'h0808;
    LUT4 i22977_3_lut (.A(n25318), .B(n25319), .C(rs2[3]), .Z(data_rs2[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22977_3_lut.init = 16'hcaca;
    LUT4 i22889_3_lut_rep_768 (.A(n25230), .B(n25231), .C(rs1[3]), .Z(n28580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22889_3_lut_rep_768.init = 16'hcaca;
    L6MUX21 i22969 (.D0(n25309), .D1(n25310), .SD(rs1[2]), .Z(n25312));
    L6MUX21 i22976 (.D0(n25316), .D1(n25317), .SD(rs2[2]), .Z(n25319));
    LUT4 i22971_4_lut_4_lut (.A(\registers[2] [7]), .B(rs2[0]), .C(rs2[1]), 
         .D(\registers[1] [7]), .Z(n25314)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i22971_4_lut_4_lut.init = 16'h2c20;
    LUT4 i22964_4_lut_4_lut (.A(\registers[2] [7]), .B(rs1[0]), .C(rs1[1]), 
         .D(\registers[1] [7]), .Z(n25307)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i22964_4_lut_4_lut.init = 16'h2c20;
    LUT4 i1_3_lut_4_lut (.A(n27231), .B(data_rs1[0]), .C(n24605), .D(\mie[12] ), 
         .Z(n928)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut.init = 16'h8f88;
    PFUMX i22807 (.BLUT(n25146), .ALUT(n25147), .C0(rs2[2]), .Z(n25150));
    L6MUX21 i22808 (.D0(n25148), .D1(n25149), .SD(rs2[2]), .Z(n25151));
    PFUMX i22814 (.BLUT(n25153), .ALUT(n25154), .C0(rs1[2]), .Z(n25157));
    L6MUX21 i22815 (.D0(n25155), .D1(n25156), .SD(rs1[2]), .Z(n25158));
    L6MUX21 i22830 (.D0(n25170), .D1(n25171), .SD(rs2[2]), .Z(n25173));
    LUT4 i22898_3_lut (.A(\registers[2] [6]), .B(\reg_access[3][2] ), .C(rs1[0]), 
         .Z(n25241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22898_3_lut.init = 16'hcaca;
    LUT4 i23546_3_lut (.A(\counter_hi[2] ), .B(n28573), .C(n28571), .Z(\reg_access[3][2] )) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(38[47:61])
    defparam i23546_3_lut.init = 16'h0404;
    L6MUX21 i22873 (.D0(n25213), .D1(n25214), .SD(rs2[2]), .Z(n25216));
    LUT4 i22897_3_lut (.A(\registers[1] [6]), .B(rs1[0]), .Z(n25240)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22897_3_lut.init = 16'h8888;
    LUT4 i22816_3_lut (.A(n25157), .B(n25158), .C(rs1[3]), .Z(data_rs1[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22816_3_lut.init = 16'hcaca;
    LUT4 i22816_3_lut_rep_769 (.A(n25157), .B(n25158), .C(rs1[3]), .Z(n28581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22816_3_lut_rep_769.init = 16'hcaca;
    L6MUX21 i22888 (.D0(n25228), .D1(n25229), .SD(rs1[2]), .Z(n25231));
    L6MUX21 i22910 (.D0(n25250), .D1(n25251), .SD(rs1[2]), .Z(n25253));
    PFUMX i22966 (.BLUT(n8_adj_2615), .ALUT(n9_adj_2614), .C0(rs1[1]), 
          .Z(n25309));
    PFUMX i22967 (.BLUT(n11_adj_2613), .ALUT(n12_adj_2612), .C0(rs1[1]), 
          .Z(n25310));
    PFUMX i22973 (.BLUT(n8_adj_2611), .ALUT(n9_adj_2610), .C0(rs2[1]), 
          .Z(n25316));
    PFUMX i22974 (.BLUT(n11_adj_2609), .ALUT(n12_adj_2608), .C0(rs2[1]), 
          .Z(n25317));
    LUT4 i22810_4_lut_4_lut (.A(\registers[2] [5]), .B(rs1[0]), .C(rs1[1]), 
         .D(\registers[1] [5]), .Z(n25153)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i22810_4_lut_4_lut.init = 16'h2c20;
    LUT4 i22803_4_lut_4_lut (.A(\registers[2] [5]), .B(rs2[0]), .C(rs2[1]), 
         .D(\registers[1] [5]), .Z(n25146)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i22803_4_lut_4_lut.init = 16'h2c20;
    LUT4 mux_1554_i1_3_lut_4_lut_4_lut (.A(rd[0]), .B(n27205), .C(n27113), 
         .D(any_additional_mem_ops), .Z(n2356)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam mux_1554_i1_3_lut_4_lut_4_lut.init = 16'h5ccc;
    LUT4 i23039_3_lut_4_lut (.A(\registers[5] [5]), .B(rs2[0]), .C(rs2[1]), 
         .D(n5_adj_2605), .Z(n25147)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i23039_3_lut_4_lut.init = 16'hf808;
    LUT4 i23036_3_lut_4_lut (.A(\registers[5] [5]), .B(rs1[0]), .C(rs1[1]), 
         .D(n5_adj_2600), .Z(n25154)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i23036_3_lut_4_lut.init = 16'hf808;
    PFUMX i22805 (.BLUT(n8_adj_2604), .ALUT(n9_adj_2603), .C0(rs2[1]), 
          .Z(n25148));
    PFUMX i22806 (.BLUT(n11_adj_2602), .ALUT(n12_adj_2601), .C0(rs2[1]), 
          .Z(n25149));
    LUT4 i1_3_lut_4_lut_adj_239 (.A(n27231), .B(data_rs1[0]), .C(n24605), 
         .D(\mie[8] ), .Z(n895)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_239.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_240 (.A(n27231), .B(data_rs1[0]), .C(n24605), 
         .D(\mie[4] ), .Z(n862)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_240.init = 16'h8f88;
    LUT4 i22876_3_lut (.A(\registers[2] [4]), .B(\reg_access[4][3] ), .C(rs1[0]), 
         .Z(n25219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22876_3_lut.init = 16'hcaca;
    PFUMX i22812 (.BLUT(n8), .ALUT(n9), .C0(rs1[1]), .Z(n25155));
    LUT4 i22875_3_lut (.A(\registers[1] [4]), .B(rs1[0]), .Z(n25218)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22875_3_lut.init = 16'h8888;
    PFUMX i22813 (.BLUT(n11), .ALUT(n12), .C0(rs1[1]), .Z(n25156));
    LUT4 i22861_3_lut (.A(\registers[2] [4]), .B(\reg_access[4][3] ), .C(rs2[0]), 
         .Z(n25204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22861_3_lut.init = 16'hcaca;
    LUT4 i22860_3_lut (.A(\registers[1] [4]), .B(rs2[0]), .Z(n25203)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22860_3_lut.init = 16'h8888;
    LUT4 i22818_3_lut (.A(\registers[2] [6]), .B(\reg_access[3][2] ), .C(rs2[0]), 
         .Z(n25161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22818_3_lut.init = 16'hcaca;
    LUT4 i22817_3_lut (.A(\registers[1] [6]), .B(rs2[0]), .Z(n25160)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22817_3_lut.init = 16'h8888;
    PFUMX i22826 (.BLUT(n25162), .ALUT(n25163), .C0(rs2[1]), .Z(n25169));
    LUT4 i22809_3_lut (.A(n25150), .B(n25151), .C(rs2[3]), .Z(data_rs2[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22809_3_lut.init = 16'hcaca;
    PFUMX i22827 (.BLUT(n25164), .ALUT(n25165), .C0(rs2[1]), .Z(n25170));
    PFUMX i22828 (.BLUT(n25166), .ALUT(n25167), .C0(rs2[1]), .Z(n25171));
    PFUMX i22869 (.BLUT(n25205), .ALUT(n25206), .C0(rs2[1]), .Z(n25212));
    PFUMX i22870 (.BLUT(n25207), .ALUT(n25208), .C0(rs2[1]), .Z(n25213));
    PFUMX i22871 (.BLUT(n25209), .ALUT(n25210), .C0(rs2[1]), .Z(n25214));
    PFUMX i22884 (.BLUT(n25220), .ALUT(n25221), .C0(rs1[1]), .Z(n25227));
    PFUMX i22885 (.BLUT(n25222), .ALUT(n25223), .C0(rs1[1]), .Z(n25228));
    L6MUX21 i22831 (.D0(n25172), .D1(n25173), .SD(rs2[3]), .Z(data_rs2[2]));
    L6MUX21 i22874 (.D0(n25215), .D1(n25216), .SD(rs2[3]), .Z(data_rs2[0]));
    L6MUX21 i22911 (.D0(n25252), .D1(n25253), .SD(rs1[3]), .Z(data_rs1[2]));
    PFUMX i22968 (.BLUT(n25307), .ALUT(n25308), .C0(rs1[2]), .Z(n25311));
    PFUMX i22975 (.BLUT(n25314), .ALUT(n25315), .C0(rs2[2]), .Z(n25318));
    PFUMX i22886 (.BLUT(n25224), .ALUT(n25225), .C0(rs1[1]), .Z(n25229));
    L6MUX21 i22829 (.D0(n25168), .D1(n25169), .SD(rs2[2]), .Z(n25172));
    L6MUX21 i22872 (.D0(n25211), .D1(n25212), .SD(rs2[2]), .Z(n25215));
    L6MUX21 i22887 (.D0(n25226), .D1(n25227), .SD(rs1[2]), .Z(n25230));
    L6MUX21 i22909 (.D0(n25248), .D1(n25249), .SD(rs1[2]), .Z(n25252));
    PFUMX i22906 (.BLUT(n25242), .ALUT(n25243), .C0(rs1[1]), .Z(n25249));
    PFUMX i22907 (.BLUT(n25244), .ALUT(n25245), .C0(rs1[1]), .Z(n25250));
    PFUMX i22908 (.BLUT(n25246), .ALUT(n25247), .C0(rs1[1]), .Z(n25251));
    
endmodule
//
// Verilog Description of module tinyqv_counter_U0
//

module tinyqv_counter_U0 (cy, clk_c, n27326, \increment_result_3__N_1925[0] , 
            instrret_count, n27229, n27246) /* synthesis syn_module_defined=1 */ ;
    output cy;
    input clk_c;
    input n27326;
    input \increment_result_3__N_1925[0] ;
    output [3:0]instrret_count;
    input n27229;
    input n27246;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [4:0]increment_result_3__N_1925;
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    
    FD1S3IX cy_51 (.D(increment_result_3__N_1925[4]), .CK(clk_c), .CD(n27326), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3IX register_2__48 (.D(increment_result_3__N_1925[2]), .CK(clk_c), 
            .CD(n27326), .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result_3__N_1925[1]), .CK(clk_c), 
            .CD(n27326), .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(\increment_result_3__N_1925[0] ), .CK(clk_c), 
            .CD(n27326), .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(register[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(register[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(register[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(instrret_count[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(register[10]), .CK(clk_c), .Q(instrret_count[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(register[9]), .CK(clk_c), .Q(instrret_count[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(register[8]), .CK(clk_c), .Q(instrret_count[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result_3__N_1925[3]), .CK(clk_c), 
            .CD(n27326), .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 i4126_2_lut_3_lut_4_lut (.A(instrret_count[1]), .B(n27229), .C(instrret_count[3]), 
         .D(instrret_count[2]), .Z(increment_result_3__N_1925[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4126_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4128_2_lut_3_lut_4_lut (.A(instrret_count[1]), .B(n27229), .C(instrret_count[3]), 
         .D(instrret_count[2]), .Z(increment_result_3__N_1925[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4128_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4112_2_lut_3_lut (.A(instrret_count[0]), .B(n27246), .C(instrret_count[1]), 
         .Z(increment_result_3__N_1925[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4112_2_lut_3_lut.init = 16'h7878;
    LUT4 i4119_2_lut_3_lut_4_lut (.A(instrret_count[0]), .B(n27246), .C(instrret_count[2]), 
         .D(instrret_count[1]), .Z(increment_result_3__N_1925[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4119_2_lut_3_lut_4_lut.init = 16'h78f0;
    
endmodule
//
// Verilog Description of module \tinyqv_counter(OUTPUT_WIDTH=7) 
//

module \tinyqv_counter(OUTPUT_WIDTH=7)  (cy, clk_c, n27326, \increment_result_3__N_1911[1] , 
            \increment_result_3__N_1911[0] , cycle_count_wide, n27228, 
            n27245, n27180) /* synthesis syn_module_defined=1 */ ;
    output cy;
    input clk_c;
    input n27326;
    input \increment_result_3__N_1911[1] ;
    input \increment_result_3__N_1911[0] ;
    output [6:0]cycle_count_wide;
    input n27228;
    input n27245;
    output n27180;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [4:0]increment_result_3__N_1911;
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    
    FD1S3IX cy_51 (.D(increment_result_3__N_1911[4]), .CK(clk_c), .CD(n27326), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3IX register_2__48 (.D(increment_result_3__N_1911[2]), .CK(clk_c), 
            .CD(n27326), .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(\increment_result_3__N_1911[1] ), .CK(clk_c), 
            .CD(n27326), .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(\increment_result_3__N_1911[0] ), .CK(clk_c), 
            .CD(n27326), .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(cycle_count_wide[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(cycle_count_wide[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(cycle_count_wide[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(cycle_count_wide[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(cycle_count_wide[6]), .CK(clk_c), .Q(cycle_count_wide[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(cycle_count_wide[5]), .CK(clk_c), .Q(cycle_count_wide[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(cycle_count_wide[4]), .CK(clk_c), .Q(cycle_count_wide[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result_3__N_1911[3]), .CK(clk_c), 
            .CD(n27326), .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 i4100_2_lut_3_lut_4_lut (.A(cycle_count_wide[1]), .B(n27228), .C(cycle_count_wide[3]), 
         .D(cycle_count_wide[2]), .Z(increment_result_3__N_1911[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4100_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4098_2_lut_3_lut_4_lut (.A(cycle_count_wide[1]), .B(n27228), .C(cycle_count_wide[3]), 
         .D(cycle_count_wide[2]), .Z(increment_result_3__N_1911[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4098_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4093_2_lut_rep_555_3_lut_4_lut (.A(cycle_count_wide[0]), .B(n27245), 
         .C(cycle_count_wide[2]), .D(cycle_count_wide[1]), .Z(n27180)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4093_2_lut_rep_555_3_lut_4_lut.init = 16'h8000;
    LUT4 i4091_2_lut_3_lut_4_lut (.A(cycle_count_wide[0]), .B(n27245), .C(cycle_count_wide[2]), 
         .D(cycle_count_wide[1]), .Z(increment_result_3__N_1911[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4091_2_lut_3_lut_4_lut.init = 16'h78f0;
    
endmodule
//
// Verilog Description of module tinyqv_alu
//

module tinyqv_alu (alu_a_in, n27187, n24124, alu_b_in, \alu_op[2] , 
            n27188, n27252, n27215, n27154, n27181, n23342, n26482, 
            n27267, cy_out, n27266, n26484, n4528, n27270, alu_out) /* synthesis syn_module_defined=1 */ ;
    input [3:0]alu_a_in;
    input n27187;
    input n24124;
    input [3:0]alu_b_in;
    input \alu_op[2] ;
    input n27188;
    input n27252;
    input n27215;
    input n27154;
    input n27181;
    input n23342;
    output n26482;
    input n27267;
    output cy_out;
    input n27266;
    output n26484;
    input [3:0]n4528;
    input n27270;
    output [3:0]alu_out;
    
    
    wire n28561, n27125, n28560, n6, n24499, n24068, n27216, n27134;
    wire [3:0]n4538;
    
    wire n27155, n27120, n27119, n26483, n24026;
    wire [3:0]a_xor_b;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[16:23])
    
    wire n24020, cmp_res_N_1855;
    wire [3:0]n4547;
    
    LUT4 i4687_4_lut_rep_756 (.A(alu_a_in[2]), .B(n28561), .C(n27125), 
         .D(n27187), .Z(n28560)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4687_4_lut_rep_756.init = 16'haaa8;
    LUT4 i4068_2_lut_3_lut_4_lut_4_lut (.A(alu_a_in[2]), .B(n28561), .C(n27125), 
         .D(n27187), .Z(n6)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4068_2_lut_3_lut_4_lut_4_lut.init = 16'hfea8;
    LUT4 i22224_4_lut (.A(alu_a_in[0]), .B(n24124), .C(alu_b_in[0]), .D(\alu_op[2] ), 
         .Z(n24499)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam i22224_4_lut.init = 16'h5a66;
    LUT4 i4059_2_lut_rep_500_3_lut_4_lut_4_lut (.A(alu_a_in[0]), .B(n27188), 
         .C(n27252), .D(n27215), .Z(n27125)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4059_2_lut_rep_500_3_lut_4_lut_4_lut.init = 16'he800;
    LUT4 mux_2762_i2_4_lut (.A(n24068), .B(n27216), .C(\alu_op[2] ), .D(n27134), 
         .Z(n4538[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_2762_i2_4_lut.init = 16'hc5ca;
    LUT4 i4697_4_lut_rep_757 (.A(alu_a_in[1]), .B(n27154), .C(n27155), 
         .D(n27215), .Z(n28561)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4697_4_lut_rep_757.init = 16'haaa8;
    LUT4 i4061_2_lut_rep_495_3_lut_4_lut_4_lut (.A(alu_a_in[1]), .B(n27154), 
         .C(n27155), .D(n27215), .Z(n27120)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4061_2_lut_rep_495_3_lut_4_lut_4_lut.init = 16'hfea8;
    LUT4 n6205_bdd_4_lut (.A(n27119), .B(n28560), .C(n27181), .D(alu_a_in[3]), 
         .Z(n26483)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+(D)))) */ ;
    defparam n6205_bdd_4_lut.init = 16'hf110;
    LUT4 mux_2762_i3_4_lut (.A(n24026), .B(a_xor_b[2]), .C(\alu_op[2] ), 
         .D(n27120), .Z(n4538[2])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_2762_i3_4_lut.init = 16'hc5ca;
    LUT4 mux_2762_i4_4_lut (.A(n24020), .B(a_xor_b[3]), .C(\alu_op[2] ), 
         .D(n6), .Z(n4538[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_2762_i4_4_lut.init = 16'hc5ca;
    LUT4 a_3__I_0_29_i3_2_lut (.A(alu_a_in[2]), .B(alu_b_in[2]), .Z(a_xor_b[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i3_2_lut.init = 16'h6666;
    LUT4 a_3__I_0_29_i4_2_lut (.A(alu_a_in[3]), .B(alu_b_in[3]), .Z(a_xor_b[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i4_2_lut.init = 16'h6666;
    LUT4 i1_4_lut (.A(a_xor_b[2]), .B(a_xor_b[3]), .C(a_xor_b[0]), .D(n23342), 
         .Z(cmp_res_N_1855)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    LUT4 a_3__I_0_29_i1_2_lut (.A(alu_a_in[0]), .B(alu_b_in[0]), .Z(a_xor_b[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i1_2_lut.init = 16'h6666;
    LUT4 alu_op_in_0__bdd_4_lut (.A(n27119), .B(n28560), .C(n27181), .D(alu_a_in[3]), 
         .Z(n26482)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C (D))))) */ ;
    defparam alu_op_in_0__bdd_4_lut.init = 16'h011f;
    LUT4 i1_2_lut_3_lut (.A(alu_b_in[3]), .B(n27267), .C(alu_a_in[3]), 
         .Z(n24020)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut.init = 16'h9696;
    LUT4 i4075_4_lut_4_lut (.A(alu_a_in[3]), .B(n27119), .C(n28560), .D(n27181), 
         .Z(cy_out)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4075_4_lut_4_lut.init = 16'hfea8;
    LUT4 i1_2_lut_3_lut_adj_237 (.A(alu_b_in[2]), .B(n27267), .C(alu_a_in[2]), 
         .Z(n24026)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut_adj_237.init = 16'h9696;
    LUT4 i4702_3_lut_rep_530_4_lut (.A(alu_b_in[0]), .B(n27267), .C(n27252), 
         .D(alu_a_in[0]), .Z(n27155)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i4702_3_lut_rep_530_4_lut.init = 16'hf600;
    LUT4 i4054_2_lut_rep_509_3_lut_3_lut_4_lut (.A(alu_b_in[0]), .B(n27267), 
         .C(n27252), .D(alu_a_in[0]), .Z(n27134)) /* synthesis lut_function=(A (B (C (D))+!B (C+(D)))+!A (B (C+(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i4054_2_lut_rep_509_3_lut_3_lut_4_lut.init = 16'hf660;
    LUT4 i4066_2_lut_rep_494_3_lut_4_lut (.A(n27215), .B(n27134), .C(n27187), 
         .D(n28561), .Z(n27119)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4066_2_lut_rep_494_3_lut_4_lut.init = 16'hf080;
    PFUMX i23980 (.BLUT(cmp_res_N_1855), .ALUT(n26483), .C0(n27266), .Z(n26484));
    PFUMX mux_2767_i4 (.BLUT(n4538[3]), .ALUT(n4528[3]), .C0(n27266), 
          .Z(n4547[3]));
    PFUMX mux_2767_i3 (.BLUT(n4538[2]), .ALUT(n4528[2]), .C0(n27266), 
          .Z(n4547[2]));
    PFUMX mux_2767_i2 (.BLUT(n4538[1]), .ALUT(n4528[1]), .C0(n27266), 
          .Z(n4547[1]));
    PFUMX mux_2767_i1 (.BLUT(n24499), .ALUT(n4528[0]), .C0(n27266), .Z(n4547[0]));
    LUT4 i1_2_lut_3_lut_adj_238 (.A(alu_b_in[1]), .B(n27267), .C(alu_a_in[1]), 
         .Z(n24068)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut_adj_238.init = 16'h9696;
    LUT4 a_3__I_0_29_i2_2_lut_rep_591 (.A(alu_a_in[1]), .B(alu_b_in[1]), 
         .Z(n27216)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i2_2_lut_rep_591.init = 16'h6666;
    LUT4 i12618_2_lut_4_lut (.A(n27270), .B(\alu_op[2] ), .C(n27266), 
         .D(n4547[1]), .Z(alu_out[1])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i12618_2_lut_4_lut.init = 16'hc500;
    LUT4 i12281_2_lut_4_lut (.A(n27270), .B(\alu_op[2] ), .C(n27266), 
         .D(n4547[0]), .Z(alu_out[0])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i12281_2_lut_4_lut.init = 16'hc500;
    LUT4 i12620_2_lut_4_lut (.A(n27270), .B(\alu_op[2] ), .C(n27266), 
         .D(n4547[3]), .Z(alu_out[3])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i12620_2_lut_4_lut.init = 16'hc500;
    LUT4 i12619_2_lut_4_lut (.A(n27270), .B(\alu_op[2] ), .C(n27266), 
         .D(n4547[2]), .Z(alu_out[2])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i12619_2_lut_4_lut.init = 16'hc500;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module sim_qspi_pmod
//

module sim_qspi_pmod (qspi_data_in, qspi_clk_N_56, spi_clk_pos_derived_59, 
            GND_net, VCC_net, qspi_data_in_3__N_1, \addr[14] , \addr_24__N_228[14] , 
            \addr[13] , \addr[12] , \addr[11] , \addr[10] , \addr[9] , 
            \addr[8] , writing, \addr[7] , \addr[6] , \addr[5] , \addr[4] , 
            \addr[3] , \addr[2] , \addr[1] , n24803, \addr[0] , qspi_ram_a_select, 
            \addr_24__N_228[0] , n22999, \writing_N_164[3] , qspi_ram_b_select, 
            \addr_24__N_228[12] , \addr_24__N_228[2] , \addr_24__N_228[1] , 
            \addr_24__N_228[3] , \addr_24__N_228[4] , \addr_24__N_228[5] , 
            \addr_24__N_228[6] , \addr_24__N_228[7] , \addr_24__N_228[8] , 
            \addr_24__N_228[9] , \addr_24__N_228[10] , \addr_24__N_228[13] , 
            \addr_24__N_228[11] , n27335, n24428) /* synthesis syn_module_defined=1 */ ;
    output [3:0]qspi_data_in;
    input qspi_clk_N_56;
    input spi_clk_pos_derived_59;
    input GND_net;
    input VCC_net;
    input [3:0]qspi_data_in_3__N_1;
    output \addr[14] ;
    input \addr_24__N_228[14] ;
    output \addr[13] ;
    output \addr[12] ;
    output \addr[11] ;
    output \addr[10] ;
    output \addr[9] ;
    output \addr[8] ;
    output writing;
    output \addr[7] ;
    output \addr[6] ;
    output \addr[5] ;
    output \addr[4] ;
    output \addr[3] ;
    output \addr[2] ;
    output \addr[1] ;
    input n24803;
    output \addr[0] ;
    input qspi_ram_a_select;
    input \addr_24__N_228[0] ;
    output n22999;
    input \writing_N_164[3] ;
    input qspi_ram_b_select;
    input \addr_24__N_228[12] ;
    input \addr_24__N_228[2] ;
    input \addr_24__N_228[1] ;
    input \addr_24__N_228[3] ;
    input \addr_24__N_228[4] ;
    input \addr_24__N_228[5] ;
    input \addr_24__N_228[6] ;
    input \addr_24__N_228[7] ;
    input \addr_24__N_228[8] ;
    input \addr_24__N_228[9] ;
    input \addr_24__N_228[10] ;
    input \addr_24__N_228[13] ;
    input \addr_24__N_228[11] ;
    output n27335;
    output n24428;
    
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire [3:0]qspi_data_out_3__N_51;
    wire [5:0]start_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(24[15:26])
    wire [5:0]n29;
    
    wire n19915, n19916;
    wire [31:0]cmd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(22[16:19])
    
    wire cmd_31__N_132;
    wire [12:0]n5639;
    wire [24:0]addr_24__N_89;
    wire [3:0]data_buff_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(29[15:27])
    
    wire spi_clk_pos_derived_59_enable_4, qspi_clk_N_56_enable_1;
    wire [11:0]n5655;
    
    wire reading, error_N_160, reading_N_139, n27387, n14418, writing_N_151, 
        n27386, reading_dummy, qspi_clk_N_56_enable_2, reading_dummy_N_262, 
        n19914, qspi_clk_N_56_enable_3, error, qspi_clk_N_56_enable_4, 
        n24805, n24680;
    wire [3:0]qspi_data_out_3__N_253;
    
    wire n24811;
    wire [7:0]ram_b_buff_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(32[16:30])
    
    wire n24673, n24677, n5738, n5746, n5753, n24734, n5742, n5750, 
        n24733, n5739, n5747, n24731, n5743, n5751, n24730, n5740, 
        n5748, n24728, n5744, n5752, n24727, n24793, n24676, n24679, 
        n5737, n5745, n24713, n5741, n5749, n24712, ram_a_buff_out_7__N_127, 
        qspi_clk_N_56_enable_5, n9644, n26618, n26617, n5690;
    wire [7:0]rom_buff_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(30[16:28])
    
    wire n26602, n26601, n27384, n24674, n26605, n26604, n5696, 
        n5704, n5732, n26501, n5716, n5724, n26500, ram_b_buff_out_7__N_131, 
        n27383;
    wire [3:0]qspi_data_out_3__N_257;
    
    wire n24794, addr_24__N_202, addr_24__N_222, addr_24__N_224, addr_24__N_220, 
        addr_24__N_218, addr_24__N_216, addr_24__N_214, addr_24__N_212, 
        addr_24__N_210, addr_24__N_208, addr_24__N_206, addr_24__N_200, 
        addr_24__N_204, n27385, n5698, n5706, n5718, n5726, n5719, 
        n5727, n5699, n5707, n5717, n5725, n5697, n5705, rom_buff_out_7__N_118, 
        n22126, n22125, ram_b_buff_out_7__N_128, n22274, n24304, n24300, 
        n24436, n24344, n24458, n24460;
    
    FD1S3AX qspi_data_out_i0 (.D(qspi_data_out_3__N_51[0]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i0.GSR = "DISABLED";
    FD1S3AX start_count_3235__i5 (.D(n29[5]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235__i5.GSR = "ENABLED";
    FD1S3AX start_count_3235__i4 (.D(n29[4]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235__i4.GSR = "ENABLED";
    FD1S3AX start_count_3235__i3 (.D(n29[3]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235__i3.GSR = "ENABLED";
    FD1S3AX start_count_3235__i2 (.D(n29[2]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235__i2.GSR = "ENABLED";
    FD1S3AX start_count_3235__i1 (.D(n29[1]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235__i1.GSR = "ENABLED";
    FD1S3AX start_count_3235__i0 (.D(n29[0]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235__i0.GSR = "ENABLED";
    CCU2C start_count_3235_add_4_5 (.A0(start_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(start_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19915), .COUT(n19916), .S0(n29[3]), .S1(n29[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235_add_4_5.INIT0 = 16'haaa0;
    defparam start_count_3235_add_4_5.INIT1 = 16'haaa0;
    defparam start_count_3235_add_4_5.INJECT1_0 = "NO";
    defparam start_count_3235_add_4_5.INJECT1_1 = "NO";
    FD1P3AX cmd_i0_i0 (.D(qspi_data_in_3__N_1[0]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i0.GSR = "ENABLED";
    FD1S3AX qspi_data_out_i3 (.D(qspi_data_out_3__N_51[3]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i3.GSR = "DISABLED";
    FD1S3AX qspi_data_out_i2 (.D(qspi_data_out_3__N_51[2]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i2.GSR = "DISABLED";
    FD1S3AX qspi_data_out_i1 (.D(qspi_data_out_3__N_51[1]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i1.GSR = "DISABLED";
    FD1S3AX addr_res1_i0_i0 (.D(addr_24__N_89[1]), .CK(qspi_clk_N_56), .Q(n5639[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i0.GSR = "ENABLED";
    FD1P3AX data_buff_in_i0_i0 (.D(qspi_data_in_3__N_1[0]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i0.GSR = "DISABLED";
    FD1P3AX addr_i14 (.D(\addr_24__N_228[14] ), .SP(qspi_clk_N_56_enable_1), 
            .CK(qspi_clk_N_56), .Q(\addr[14] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i14.GSR = "ENABLED";
    FD1S3AX addr_i13 (.D(addr_24__N_89[13]), .CK(qspi_clk_N_56), .Q(\addr[13] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i13.GSR = "ENABLED";
    FD1S3AX addr_i12 (.D(addr_24__N_89[12]), .CK(qspi_clk_N_56), .Q(\addr[12] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i12.GSR = "ENABLED";
    FD1S3AX addr_i11 (.D(addr_24__N_89[11]), .CK(qspi_clk_N_56), .Q(\addr[11] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i11.GSR = "ENABLED";
    FD1S3AX addr_i10 (.D(addr_24__N_89[10]), .CK(qspi_clk_N_56), .Q(\addr[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i10.GSR = "ENABLED";
    FD1S3AX addr_i9 (.D(addr_24__N_89[9]), .CK(qspi_clk_N_56), .Q(\addr[9] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i9.GSR = "ENABLED";
    FD1S3AX addr_res2_i0_i11 (.D(addr_24__N_89[12]), .CK(qspi_clk_N_56), 
            .Q(n5655[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res2_i0_i11.GSR = "ENABLED";
    FD1S3AX addr_i8 (.D(addr_24__N_89[8]), .CK(qspi_clk_N_56), .Q(\addr[8] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i8.GSR = "ENABLED";
    LUT4 i23560_4_lut_then_3_lut_4_lut (.A(reading), .B(writing), .C(error_N_160), 
         .D(reading_N_139), .Z(n27387)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i23560_4_lut_then_3_lut_4_lut.init = 16'h1110;
    LUT4 i23560_4_lut_else_3_lut_4_lut (.A(reading), .B(writing), .C(n14418), 
         .D(writing_N_151), .Z(n27386)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i23560_4_lut_else_3_lut_4_lut.init = 16'h0100;
    FD1S3AX addr_i7 (.D(addr_24__N_89[7]), .CK(qspi_clk_N_56), .Q(\addr[7] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i7.GSR = "ENABLED";
    FD1S3AX addr_i6 (.D(addr_24__N_89[6]), .CK(qspi_clk_N_56), .Q(\addr[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i6.GSR = "ENABLED";
    FD1S3AX addr_i5 (.D(addr_24__N_89[5]), .CK(qspi_clk_N_56), .Q(\addr[5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i5.GSR = "ENABLED";
    FD1S3AX addr_i4 (.D(addr_24__N_89[4]), .CK(qspi_clk_N_56), .Q(\addr[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i4.GSR = "ENABLED";
    FD1S3AX addr_i3 (.D(addr_24__N_89[3]), .CK(qspi_clk_N_56), .Q(\addr[3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i3.GSR = "ENABLED";
    FD1S3AX addr_i2 (.D(addr_24__N_89[2]), .CK(qspi_clk_N_56), .Q(\addr[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i2.GSR = "ENABLED";
    FD1S3AX addr_i1 (.D(addr_24__N_89[1]), .CK(qspi_clk_N_56), .Q(\addr[1] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i1.GSR = "ENABLED";
    FD1P3AX reading_dummy_116 (.D(reading_dummy_N_262), .SP(qspi_clk_N_56_enable_2), 
            .CK(qspi_clk_N_56), .Q(reading_dummy)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam reading_dummy_116.GSR = "ENABLED";
    CCU2C start_count_3235_add_4_7 (.A0(start_count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19916), .S0(n29[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235_add_4_7.INIT0 = 16'haaa0;
    defparam start_count_3235_add_4_7.INIT1 = 16'h0000;
    defparam start_count_3235_add_4_7.INJECT1_0 = "NO";
    defparam start_count_3235_add_4_7.INJECT1_1 = "NO";
    CCU2C start_count_3235_add_4_3 (.A0(start_count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(start_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n19914), .COUT(n19915), .S0(n29[1]), .S1(n29[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235_add_4_3.INIT0 = 16'haaa0;
    defparam start_count_3235_add_4_3.INIT1 = 16'haaa0;
    defparam start_count_3235_add_4_3.INJECT1_0 = "NO";
    defparam start_count_3235_add_4_3.INJECT1_1 = "NO";
    CCU2C start_count_3235_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n19914), .S1(n29[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3235_add_4_1.INIT0 = 16'h0000;
    defparam start_count_3235_add_4_1.INIT1 = 16'h555f;
    defparam start_count_3235_add_4_1.INJECT1_0 = "NO";
    defparam start_count_3235_add_4_1.INJECT1_1 = "NO";
    FD1P3AX writing_117 (.D(n24803), .SP(qspi_clk_N_56_enable_3), .CK(qspi_clk_N_56), 
            .Q(writing)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam writing_117.GSR = "ENABLED";
    FD1P3AX error_118 (.D(VCC_net), .SP(qspi_clk_N_56_enable_4), .CK(qspi_clk_N_56), 
            .Q(error)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam error_118.GSR = "ENABLED";
    FD1P3AX reading_115 (.D(n24805), .SP(reading_N_139), .CK(qspi_clk_N_56), 
            .Q(reading)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam reading_115.GSR = "ENABLED";
    PFUMX qspi_data_out_3__I_0_i2 (.BLUT(n24680), .ALUT(qspi_data_out_3__N_253[1]), 
          .C0(n24811), .Z(qspi_data_out_3__N_51[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    LUT4 i22330_3_lut (.A(ram_b_buff_out[7]), .B(ram_b_buff_out[3]), .C(\addr[0] ), 
         .Z(n24673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22330_3_lut.init = 16'hcaca;
    PFUMX qspi_data_out_3__I_0_i3 (.BLUT(n24677), .ALUT(qspi_data_out_3__N_253[2]), 
          .C0(n24811), .Z(qspi_data_out_3__N_51[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    LUT4 i22391_3_lut (.A(n5738), .B(n5746), .C(n5753), .Z(n24734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22391_3_lut.init = 16'hcaca;
    LUT4 i22390_3_lut (.A(n5742), .B(n5750), .C(n5753), .Z(n24733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22390_3_lut.init = 16'hcaca;
    LUT4 i22388_3_lut (.A(n5739), .B(n5747), .C(n5753), .Z(n24731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22388_3_lut.init = 16'hcaca;
    LUT4 i22387_3_lut (.A(n5743), .B(n5751), .C(n5753), .Z(n24730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22387_3_lut.init = 16'hcaca;
    LUT4 i22385_3_lut (.A(n5740), .B(n5748), .C(n5753), .Z(n24728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22385_3_lut.init = 16'hcaca;
    LUT4 i22384_3_lut (.A(n5744), .B(n5752), .C(n5753), .Z(n24727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22384_3_lut.init = 16'hcaca;
    LUT4 i22450_3_lut (.A(ram_b_buff_out[4]), .B(ram_b_buff_out[0]), .C(\addr[0] ), 
         .Z(n24793)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22450_3_lut.init = 16'hcaca;
    PFUMX i24341 (.BLUT(n27386), .ALUT(n27387), .C0(reading_dummy), .Z(qspi_clk_N_56_enable_2));
    LUT4 i22333_3_lut (.A(ram_b_buff_out[6]), .B(ram_b_buff_out[2]), .C(\addr[0] ), 
         .Z(n24676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22333_3_lut.init = 16'hcaca;
    LUT4 i22336_3_lut (.A(ram_b_buff_out[5]), .B(ram_b_buff_out[1]), .C(\addr[0] ), 
         .Z(n24679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22336_3_lut.init = 16'hcaca;
    LUT4 i22370_3_lut (.A(n5737), .B(n5745), .C(n5753), .Z(n24713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22370_3_lut.init = 16'hcaca;
    LUT4 i22369_3_lut (.A(n5741), .B(n5749), .C(n5753), .Z(n24712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22369_3_lut.init = 16'hcaca;
    FD1S3AX addr_res3_i0_i1 (.D(addr_24__N_89[2]), .CK(qspi_clk_N_56), .Q(n5639[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i1.GSR = "ENABLED";
    FD1S3AX addr_res3_i0_i2 (.D(addr_24__N_89[3]), .CK(qspi_clk_N_56), .Q(n5639[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i2.GSR = "ENABLED";
    FD1S3AX addr_res3_i0_i3 (.D(addr_24__N_89[4]), .CK(qspi_clk_N_56), .Q(n5639[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i3.GSR = "ENABLED";
    FD1S3AX addr_res3_i0_i4 (.D(addr_24__N_89[5]), .CK(qspi_clk_N_56), .Q(n5639[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i4.GSR = "ENABLED";
    FD1S3AX addr_res3_i0_i5 (.D(addr_24__N_89[6]), .CK(qspi_clk_N_56), .Q(n5639[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i5.GSR = "ENABLED";
    FD1S3AX addr_res3_i0_i6 (.D(addr_24__N_89[7]), .CK(qspi_clk_N_56), .Q(n5639[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i6.GSR = "ENABLED";
    FD1S3AX addr_res3_i0_i7 (.D(addr_24__N_89[8]), .CK(qspi_clk_N_56), .Q(n5639[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i7.GSR = "ENABLED";
    FD1S3AX addr_res3_i0_i8 (.D(addr_24__N_89[9]), .CK(qspi_clk_N_56), .Q(n5639[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i8.GSR = "ENABLED";
    FD1S3AX addr_res3_i0_i9 (.D(addr_24__N_89[10]), .CK(qspi_clk_N_56), 
            .Q(n5639[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i9.GSR = "ENABLED";
    FD1S3AX addr_res3_i0_i10 (.D(addr_24__N_89[11]), .CK(qspi_clk_N_56), 
            .Q(n5639[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res3_i0_i10.GSR = "ENABLED";
    LUT4 i23427_2_lut (.A(\addr[0] ), .B(qspi_ram_a_select), .Z(ram_a_buff_out_7__N_127)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i23427_2_lut.init = 16'h1111;
    FD1P3IX addr_i0 (.D(\addr_24__N_228[0] ), .SP(qspi_clk_N_56_enable_5), 
            .CD(n9644), .CK(qspi_clk_N_56), .Q(\addr[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i0.GSR = "ENABLED";
    PFUMX i24062 (.BLUT(n26618), .ALUT(n26617), .C0(n5690), .Z(rom_buff_out[1]));
    PFUMX i24051 (.BLUT(n26602), .ALUT(n26601), .C0(n5690), .Z(rom_buff_out[3]));
    FD1P3AX cmd_i0_i1 (.D(qspi_data_in_3__N_1[1]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i1.GSR = "ENABLED";
    FD1P3AX cmd_i0_i2 (.D(qspi_data_in_3__N_1[2]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i2.GSR = "ENABLED";
    FD1P3AX cmd_i0_i3 (.D(qspi_data_in_3__N_1[3]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i3.GSR = "ENABLED";
    FD1P3AX cmd_i0_i4 (.D(cmd[0]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i4.GSR = "ENABLED";
    FD1P3AX cmd_i0_i5 (.D(cmd[1]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i5.GSR = "ENABLED";
    FD1P3AX cmd_i0_i6 (.D(cmd[2]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i6.GSR = "ENABLED";
    FD1P3AX cmd_i0_i7 (.D(cmd[3]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i7.GSR = "ENABLED";
    FD1P3AX cmd_i0_i8 (.D(cmd[4]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i8.GSR = "ENABLED";
    FD1P3AX cmd_i0_i9 (.D(cmd[5]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i9.GSR = "ENABLED";
    FD1P3AX cmd_i0_i10 (.D(cmd[6]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i10.GSR = "ENABLED";
    FD1P3AX cmd_i0_i11 (.D(cmd[7]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i11.GSR = "ENABLED";
    FD1P3AX cmd_i0_i12 (.D(cmd[8]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i12.GSR = "ENABLED";
    FD1P3AX cmd_i0_i13 (.D(cmd[9]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i13.GSR = "ENABLED";
    FD1P3AX cmd_i0_i14 (.D(cmd[10]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i14.GSR = "ENABLED";
    FD1P3AX cmd_i0_i15 (.D(cmd[11]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i15.GSR = "ENABLED";
    FD1P3AX cmd_i0_i16 (.D(cmd[12]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i16.GSR = "ENABLED";
    FD1P3AX cmd_i0_i17 (.D(cmd[13]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i17.GSR = "ENABLED";
    FD1P3AX cmd_i0_i18 (.D(cmd[14]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i18.GSR = "ENABLED";
    FD1P3AX cmd_i0_i19 (.D(cmd[15]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i19.GSR = "ENABLED";
    FD1P3AX cmd_i0_i20 (.D(cmd[16]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i20.GSR = "ENABLED";
    FD1P3AX cmd_i0_i21 (.D(cmd[17]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i21.GSR = "ENABLED";
    FD1P3AX cmd_i0_i22 (.D(cmd[18]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i22.GSR = "ENABLED";
    FD1P3AX cmd_i0_i23 (.D(cmd[19]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i23.GSR = "ENABLED";
    FD1P3AX cmd_i0_i24 (.D(cmd[20]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i24.GSR = "ENABLED";
    FD1P3AX cmd_i0_i25 (.D(cmd[21]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i25.GSR = "ENABLED";
    FD1P3AX cmd_i0_i26 (.D(cmd[22]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i26.GSR = "ENABLED";
    FD1P3AX cmd_i0_i27 (.D(cmd[23]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i27.GSR = "ENABLED";
    FD1P3AX cmd_i0_i28 (.D(cmd[24]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i28.GSR = "ENABLED";
    FD1P3AX cmd_i0_i29 (.D(cmd[25]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i29.GSR = "ENABLED";
    FD1P3AX cmd_i0_i30 (.D(cmd[26]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i30.GSR = "ENABLED";
    FD1P3AX cmd_i0_i31 (.D(cmd[27]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i31.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i12 (.D(addr_24__N_89[13]), .CK(qspi_clk_N_56), 
            .Q(n5639[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i12.GSR = "ENABLED";
    LUT4 i1_4_lut_then_4_lut (.A(writing_N_151), .B(cmd[27]), .C(n22999), 
         .D(\writing_N_164[3] ), .Z(n27384)) /* synthesis lut_function=(A (B (C (D))+!B (D))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'ha200;
    PFUMX qspi_data_out_3__I_0_i4 (.BLUT(n24674), .ALUT(qspi_data_out_3__N_253[3]), 
          .C0(n24811), .Z(qspi_data_out_3__N_51[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    PFUMX i24054 (.BLUT(n26605), .ALUT(n26604), .C0(n5690), .Z(rom_buff_out[2]));
    FD1P3AX data_buff_in_i0_i1 (.D(qspi_data_in_3__N_1[1]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i1.GSR = "DISABLED";
    FD1P3AX data_buff_in_i0_i2 (.D(qspi_data_in_3__N_1[2]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i2.GSR = "DISABLED";
    FD1P3AX data_buff_in_i0_i3 (.D(qspi_data_in_3__N_1[3]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i3.GSR = "DISABLED";
    LUT4 n5716_bdd_3_lut (.A(n5696), .B(n5704), .C(n5732), .Z(n26501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n5716_bdd_3_lut.init = 16'hcaca;
    LUT4 n5716_bdd_3_lut_23987 (.A(n5716), .B(n5732), .C(n5724), .Z(n26500)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n5716_bdd_3_lut_23987.init = 16'he2e2;
    LUT4 i23430_2_lut (.A(\addr[0] ), .B(qspi_ram_b_select), .Z(ram_b_buff_out_7__N_131)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i23430_2_lut.init = 16'h1111;
    LUT4 i1_4_lut_else_4_lut (.A(writing_N_151), .B(cmd[27]), .C(n22999), 
         .D(\writing_N_164[3] ), .Z(n27383)) /* synthesis lut_function=(A (B (D)+!B (C (D)))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'ha800;
    LUT4 i22452_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[0]), 
         .C(rom_buff_out[4]), .Z(qspi_data_out_3__N_253[0])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i22452_3_lut_3_lut.init = 16'he4e4;
    LUT4 i22332_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[3]), 
         .C(rom_buff_out[7]), .Z(qspi_data_out_3__N_253[3])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i22332_3_lut_3_lut.init = 16'he4e4;
    LUT4 i22335_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[2]), 
         .C(rom_buff_out[6]), .Z(qspi_data_out_3__N_253[2])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i22335_3_lut_3_lut.init = 16'he4e4;
    LUT4 i22338_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[1]), 
         .C(rom_buff_out[5]), .Z(qspi_data_out_3__N_253[1])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i22338_3_lut_3_lut.init = 16'he4e4;
    LUT4 i23060_3_lut_3_lut (.A(qspi_ram_b_select), .B(n24673), .C(rom_buff_out[3]), 
         .Z(n24674)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i23060_3_lut_3_lut.init = 16'he4e4;
    LUT4 i23048_3_lut_3_lut (.A(qspi_ram_b_select), .B(n24793), .C(rom_buff_out[0]), 
         .Z(n24794)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i23048_3_lut_3_lut.init = 16'he4e4;
    LUT4 i23062_3_lut_3_lut (.A(qspi_ram_b_select), .B(n24676), .C(rom_buff_out[2]), 
         .Z(n24677)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i23062_3_lut_3_lut.init = 16'he4e4;
    LUT4 i23064_3_lut_3_lut (.A(qspi_ram_b_select), .B(n24679), .C(rom_buff_out[1]), 
         .Z(n24680)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i23064_3_lut_3_lut.init = 16'he4e4;
    PFUMX qspi_data_out_3__I_0_i1 (.BLUT(n24794), .ALUT(qspi_data_out_3__N_253[0]), 
          .C0(n24811), .Z(qspi_data_out_3__N_51[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    LUT4 addr_24__I_0_i13_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[12] ), 
         .D(addr_24__N_202), .Z(addr_24__N_89[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i22462_4_lut_3_lut (.A(reading), .B(writing), .C(reading_dummy), 
         .Z(n24805)) /* synthesis lut_function=(A+!(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i22462_4_lut_3_lut.init = 16'hbaba;
    LUT4 addr_24__I_0_i3_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[2] ), 
         .D(addr_24__N_222), .Z(addr_24__N_89[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(reading), .B(writing), .C(writing_N_151), 
         .D(reading_dummy), .Z(qspi_clk_N_56_enable_5)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i1_2_lut_3_lut_4_lut.init = 16'heefe;
    LUT4 i7297_2_lut_3_lut_4_lut (.A(reading), .B(writing), .C(writing_N_151), 
         .D(reading_dummy), .Z(n9644)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i7297_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 addr_24__I_0_i2_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[1] ), 
         .D(addr_24__N_224), .Z(addr_24__N_89[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i4_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[3] ), 
         .D(addr_24__N_220), .Z(addr_24__N_89[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i5_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[4] ), 
         .D(addr_24__N_218), .Z(addr_24__N_89[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i6_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[5] ), 
         .D(addr_24__N_216), .Z(addr_24__N_89[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i7_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[6] ), 
         .D(addr_24__N_214), .Z(addr_24__N_89[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i8_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[7] ), 
         .D(addr_24__N_212), .Z(addr_24__N_89[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i9_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[8] ), 
         .D(addr_24__N_210), .Z(addr_24__N_89[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i10_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[9] ), 
         .D(addr_24__N_208), .Z(addr_24__N_89[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i11_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[10] ), 
         .D(addr_24__N_206), .Z(addr_24__N_89[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i14_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[13] ), 
         .D(addr_24__N_200), .Z(addr_24__N_89[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i12_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[11] ), 
         .D(addr_24__N_204), .Z(addr_24__N_89[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23484_3_lut_rep_710 (.A(\writing_N_164[3] ), .B(qspi_ram_b_select), 
         .C(qspi_ram_a_select), .Z(n27335)) /* synthesis lut_function=(!(A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(34[23:82])
    defparam i23484_3_lut_rep_710.init = 16'h7f7f;
    LUT4 i23480_2_lut_4_lut (.A(\writing_N_164[3] ), .B(qspi_ram_b_select), 
         .C(qspi_ram_a_select), .D(\addr[0] ), .Z(spi_clk_pos_derived_59_enable_4)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(34[23:82])
    defparam i23480_2_lut_4_lut.init = 16'h007f;
    PFUMX i24339 (.BLUT(n27383), .ALUT(n27384), .C0(cmd[24]), .Z(n27385));
    PFUMX i23988 (.BLUT(n26501), .ALUT(n26500), .C0(n5690), .Z(rom_buff_out[0]));
    LUT4 n5718_bdd_3_lut (.A(n5698), .B(n5706), .C(n5732), .Z(n26605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n5718_bdd_3_lut.init = 16'hcaca;
    LUT4 n5718_bdd_3_lut_24053 (.A(n5718), .B(n5732), .C(n5726), .Z(n26604)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n5718_bdd_3_lut_24053.init = 16'he2e2;
    LUT4 n5719_bdd_3_lut_24050 (.A(n5719), .B(n5732), .C(n5727), .Z(n26601)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n5719_bdd_3_lut_24050.init = 16'he2e2;
    LUT4 n5719_bdd_3_lut (.A(n5699), .B(n5707), .C(n5732), .Z(n26602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n5719_bdd_3_lut.init = 16'hcaca;
    LUT4 n5717_bdd_3_lut_24061 (.A(n5717), .B(n5732), .C(n5725), .Z(n26617)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n5717_bdd_3_lut_24061.init = 16'he2e2;
    LUT4 n5717_bdd_3_lut (.A(n5697), .B(n5705), .C(n5732), .Z(n26618)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n5717_bdd_3_lut.init = 16'hcaca;
    LUT4 i23424_2_lut (.A(\addr[0] ), .B(\writing_N_164[3] ), .Z(rom_buff_out_7__N_118)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i23424_2_lut.init = 16'h1111;
    LUT4 i23574_3_lut (.A(reading), .B(writing), .C(error), .Z(cmd_31__N_132)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i23574_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_3_lut_4_lut_adj_228 (.A(writing), .B(\addr[0] ), .C(\addr[12] ), 
         .D(qspi_ram_a_select), .Z(n22126)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(49[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_228.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_229 (.A(writing), .B(\addr[0] ), .C(\addr[12] ), 
         .D(qspi_ram_a_select), .Z(n22125)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(49[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_229.init = 16'h0008;
    LUT4 ram_a_buff_out_7__N_124_I_0_2_lut_3_lut (.A(writing), .B(\addr[0] ), 
         .C(qspi_ram_b_select), .Z(ram_b_buff_out_7__N_128)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(49[14:31])
    defparam ram_a_buff_out_7__N_124_I_0_2_lut_3_lut.init = 16'h0808;
    LUT4 i1_4_lut (.A(start_count[3]), .B(n22274), .C(n24304), .D(\writing_N_164[3] ), 
         .Z(writing_N_151)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h2010;
    LUT4 i1_4_lut_adj_230 (.A(start_count[0]), .B(n24300), .C(start_count[1]), 
         .D(\writing_N_164[3] ), .Z(n24304)) /* synthesis lut_function=(!(A+((C (D)+!C !(D))+!B))) */ ;
    defparam i1_4_lut_adj_230.init = 16'h0440;
    LUT4 i1_3_lut (.A(start_count[2]), .B(error), .C(\writing_N_164[3] ), 
         .Z(n24300)) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(C)))) */ ;
    defparam i1_3_lut.init = 16'h1212;
    LUT4 i20056_2_lut (.A(start_count[5]), .B(start_count[4]), .Z(n22274)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20056_2_lut.init = 16'heeee;
    PFUMX i22371 (.BLUT(n24712), .ALUT(n24713), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[0]));
    PFUMX i22386 (.BLUT(n24727), .ALUT(n24728), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[3]));
    PFUMX i22389 (.BLUT(n24730), .ALUT(n24731), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[2]));
    PFUMX i22392 (.BLUT(n24733), .ALUT(n24734), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[1]));
    LUT4 i23529_3_lut (.A(qspi_ram_a_select), .B(qspi_ram_b_select), .C(\addr[0] ), 
         .Z(n24811)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26] 113[96])
    defparam i23529_3_lut.init = 16'h5d5d;
    LUT4 i23511_4_lut (.A(start_count[2]), .B(start_count[3]), .C(n24436), 
         .D(n22274), .Z(reading_N_139)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(93[21:38])
    defparam i23511_4_lut.init = 16'h0008;
    LUT4 i1_2_lut (.A(start_count[0]), .B(start_count[1]), .Z(n24436)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(93[21:38])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_231 (.A(n24344), .B(n22274), .C(start_count[3]), 
         .D(cmd[3]), .Z(error_N_160)) /* synthesis lut_function=(!(A (B+(C))+!A (B+(C+(D))))) */ ;
    defparam i1_4_lut_adj_231.init = 16'h0203;
    LUT4 i1_3_lut_adj_232 (.A(cmd[1]), .B(cmd[2]), .C(cmd[0]), .Z(n24344)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_3_lut_adj_232.init = 16'hfdfd;
    LUT4 i12117_4_lut (.A(\writing_N_164[3] ), .B(cmd[27]), .C(n22999), 
         .D(cmd[24]), .Z(n14418)) /* synthesis lut_function=(A ((C+!(D))+!B)) */ ;
    defparam i12117_4_lut.init = 16'ha2aa;
    LUT4 i1_4_lut_adj_233 (.A(n24458), .B(cmd[25]), .C(n24460), .D(cmd[26]), 
         .Z(n22999)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_233.init = 16'hfffb;
    LUT4 i1_2_lut_adj_234 (.A(cmd[31]), .B(cmd[30]), .Z(n24458)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_234.init = 16'heeee;
    LUT4 i1_2_lut_adj_235 (.A(cmd[29]), .B(cmd[28]), .Z(n24460)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_235.init = 16'heeee;
    LUT4 reading_I_0_126_2_lut_rep_761 (.A(reading), .B(writing), .Z(qspi_clk_N_56_enable_1)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam reading_I_0_126_2_lut_rep_761.init = 16'heeee;
    LUT4 i7252_2_lut_3_lut (.A(n14418), .B(writing_N_151), .C(reading_dummy), 
         .Z(reading_dummy_N_262)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i7252_2_lut_3_lut.init = 16'h0404;
    LUT4 i2_2_lut_rep_618 (.A(reading_dummy), .B(writing_N_151), .Z(qspi_clk_N_56_enable_3)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i2_2_lut_rep_618.init = 16'h4444;
    LUT4 i4572_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[0]), 
         .D(\addr[1] ), .Z(addr_24__N_224)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4572_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4548_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[12]), 
         .D(\addr[13] ), .Z(addr_24__N_200)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4548_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4550_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[11]), 
         .D(\addr[12] ), .Z(addr_24__N_202)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4550_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4552_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[10]), 
         .D(\addr[11] ), .Z(addr_24__N_204)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4552_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4554_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[9]), 
         .D(\addr[10] ), .Z(addr_24__N_206)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4554_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4556_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[8]), 
         .D(\addr[9] ), .Z(addr_24__N_208)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4556_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4558_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[7]), 
         .D(\addr[8] ), .Z(addr_24__N_210)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4558_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4560_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[6]), 
         .D(\addr[7] ), .Z(addr_24__N_212)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4560_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4562_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[5]), 
         .D(\addr[6] ), .Z(addr_24__N_214)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4562_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4564_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[4]), 
         .D(\addr[5] ), .Z(addr_24__N_216)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4564_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4566_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[3]), 
         .D(\addr[4] ), .Z(addr_24__N_218)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4566_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_adj_236 (.A(cmd[27]), .B(cmd[24]), .C(qspi_clk_N_56_enable_1), 
         .D(\writing_N_164[3] ), .Z(n24428)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_236.init = 16'h0100;
    LUT4 i4568_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[2]), 
         .D(\addr[3] ), .Z(addr_24__N_220)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4568_3_lut_4_lut.init = 16'hfb40;
    LUT4 i4570_3_lut_4_lut (.A(reading_dummy), .B(writing_N_151), .C(cmd[1]), 
         .D(\addr[2] ), .Z(addr_24__N_222)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i4570_3_lut_4_lut.init = 16'hfb40;
    LUT4 i23551_4_lut (.A(n27385), .B(qspi_clk_N_56_enable_1), .C(error_N_160), 
         .D(reading_dummy), .Z(qspi_clk_N_56_enable_4)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i23551_4_lut.init = 16'h3022;
    \BRAM(ADDR_WIDTH=13,INIT_FILE="ledstrip.hex")  rom (.\addr[1] (\addr[1] ), 
            .\addr[2] (\addr[2] ), .\addr[3] (\addr[3] ), .\addr[4] (\addr[4] ), 
            .\addr[5] (\addr[5] ), .\addr[6] (\addr[6] ), .\addr[7] (\addr[7] ), 
            .\addr[8] (\addr[8] ), .\addr[9] (\addr[9] ), .\addr[10] (\addr[10] ), 
            .\addr[11] (\addr[11] ), .n5643(n5639[0]), .n5638(n5639[1]), 
            .n5637(n5639[2]), .n5636(n5639[3]), .n5635(n5639[4]), .n5634(n5639[5]), 
            .n5633(n5639[6]), .n5632(n5639[7]), .n5631(n5639[8]), .n5630(n5639[9]), 
            .n5629(n5639[10]), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .data_buff_in({data_buff_in}), .n5696(n5696), .n5697(n5697), 
            .n5698(n5698), .n5699(n5699), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .GND_net(GND_net), .rom_buff_out_7__N_118(rom_buff_out_7__N_118), 
            .VCC_net(VCC_net), .n5690(n5690), .n5627(n5639[12]), .n5704(n5704), 
            .n5705(n5705), .n5706(n5706), .n5707(n5707), .n5732(n5732), 
            .n5644(n5655[11]), .n5724(n5724), .n5725(n5725), .n5726(n5726), 
            .n5727(n5727), .n5716(n5716), .n5717(n5717), .n5718(n5718), 
            .n5719(n5719), .\rom_buff_out[5] (rom_buff_out[5]), .\rom_buff_out[4] (rom_buff_out[4]), 
            .\rom_buff_out[7] (rom_buff_out[7]), .\rom_buff_out[6] (rom_buff_out[6])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(36[58] 43[6])
    \BRAM(ADDR_WIDTH=11)  ram_b (.\addr[1] (\addr[1] ), .\addr[2] (\addr[2] ), 
            .\addr[3] (\addr[3] ), .\addr[4] (\addr[4] ), .\addr[5] (\addr[5] ), 
            .\addr[6] (\addr[6] ), .\addr[7] (\addr[7] ), .\addr[8] (\addr[8] ), 
            .\addr[9] (\addr[9] ), .\addr[10] (\addr[10] ), .\addr[11] (\addr[11] ), 
            .n5643(n5639[0]), .n5638(n5639[1]), .n5637(n5639[2]), .n5636(n5639[3]), 
            .n5635(n5639[4]), .n5634(n5639[5]), .n5633(n5639[6]), .n5632(n5639[7]), 
            .n5631(n5639[8]), .n5630(n5639[9]), .n5629(n5639[10]), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .data_buff_in({data_buff_in}), .ram_b_buff_out({ram_b_buff_out}), 
            .spi_clk_pos_derived_59(spi_clk_pos_derived_59), .ram_b_buff_out_7__N_128(ram_b_buff_out_7__N_128), 
            .ram_b_buff_out_7__N_131(ram_b_buff_out_7__N_131), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(52[37] 59[6])
    \BRAM(ADDR_WIDTH=12)  ram_a (.\addr[1] (\addr[1] ), .\addr[2] (\addr[2] ), 
            .\addr[3] (\addr[3] ), .\addr[4] (\addr[4] ), .\addr[5] (\addr[5] ), 
            .\addr[6] (\addr[6] ), .\addr[7] (\addr[7] ), .\addr[8] (\addr[8] ), 
            .\addr[9] (\addr[9] ), .\addr[10] (\addr[10] ), .\addr[11] (\addr[11] ), 
            .n5643(n5639[0]), .n5638(n5639[1]), .n5637(n5639[2]), .n5636(n5639[3]), 
            .n5635(n5639[4]), .n5634(n5639[5]), .n5633(n5639[6]), .n5632(n5639[7]), 
            .n5631(n5639[8]), .n5630(n5639[9]), .n5629(n5639[10]), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .data_buff_in({data_buff_in}), .n5745(n5745), .n5746(n5746), 
            .n5747(n5747), .n5748(n5748), .n5749(n5749), .n5750(n5750), 
            .n5751(n5751), .n5752(n5752), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .n22126(n22126), .ram_a_buff_out_7__N_127(ram_a_buff_out_7__N_127), 
            .GND_net(GND_net), .VCC_net(VCC_net), .n5753(n5753), .n5644(n5655[11]), 
            .n5737(n5737), .n5738(n5738), .n5739(n5739), .n5740(n5740), 
            .n5741(n5741), .n5742(n5742), .n5743(n5743), .n5744(n5744), 
            .n22125(n22125)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(44[37] 51[6])
    
endmodule
//
// Verilog Description of module \BRAM(ADDR_WIDTH=13,INIT_FILE="ledstrip.hex") 
//

module \BRAM(ADDR_WIDTH=13,INIT_FILE="ledstrip.hex")  (\addr[1] , \addr[2] , 
            \addr[3] , \addr[4] , \addr[5] , \addr[6] , \addr[7] , 
            \addr[8] , \addr[9] , \addr[10] , \addr[11] , n5643, n5638, 
            n5637, n5636, n5635, n5634, n5633, n5632, n5631, n5630, 
            n5629, qspi_data_in_3__N_1, data_buff_in, n5696, n5697, 
            n5698, n5699, spi_clk_pos_derived_59, GND_net, rom_buff_out_7__N_118, 
            VCC_net, n5690, n5627, n5704, n5705, n5706, n5707, 
            n5732, n5644, n5724, n5725, n5726, n5727, n5716, n5717, 
            n5718, n5719, \rom_buff_out[5] , \rom_buff_out[4] , \rom_buff_out[7] , 
            \rom_buff_out[6] ) /* synthesis syn_module_defined=1 */ ;
    input \addr[1] ;
    input \addr[2] ;
    input \addr[3] ;
    input \addr[4] ;
    input \addr[5] ;
    input \addr[6] ;
    input \addr[7] ;
    input \addr[8] ;
    input \addr[9] ;
    input \addr[10] ;
    input \addr[11] ;
    input n5643;
    input n5638;
    input n5637;
    input n5636;
    input n5635;
    input n5634;
    input n5633;
    input n5632;
    input n5631;
    input n5630;
    input n5629;
    input [3:0]qspi_data_in_3__N_1;
    input [3:0]data_buff_in;
    output n5696;
    output n5697;
    output n5698;
    output n5699;
    input spi_clk_pos_derived_59;
    input GND_net;
    input rom_buff_out_7__N_118;
    input VCC_net;
    output n5690;
    input n5627;
    output n5704;
    output n5705;
    output n5706;
    output n5707;
    output n5732;
    input n5644;
    output n5724;
    output n5725;
    output n5726;
    output n5727;
    output n5716;
    output n5717;
    output n5718;
    output n5719;
    output \rom_buff_out[5] ;
    output \rom_buff_out[4] ;
    output \rom_buff_out[7] ;
    output \rom_buff_out[6] ;
    
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    wire n5700, n5701, n5702, n5703, n5708, n5709, n5710, n5711, 
        n5728, n5729, n5730, n5731, n5720, n5721, n5722, n5723, 
        n24770, n24769, n24767, n24766, n24761, n24760, n24716, 
        n24715;
    
    DP16KD mem0 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n5643), .ADB4(n5638), 
           .ADB5(n5637), .ADB6(n5636), .ADB7(n5635), .ADB8(n5634), .ADB9(n5633), 
           .ADB10(n5632), .ADB11(n5631), .ADB12(n5630), .ADB13(n5629), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n5696), .DOB1(n5697), .DOB2(n5698), 
           .DOB3(n5699), .DOB4(n5700), .DOB5(n5701), .DOB6(n5702), .DOB7(n5703));
    defparam mem0.DATA_WIDTH_A = 9;
    defparam mem0.DATA_WIDTH_B = 9;
    defparam mem0.REGMODE_A = "NOREG";
    defparam mem0.REGMODE_B = "NOREG";
    defparam mem0.RESETMODE = "SYNC";
    defparam mem0.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem0.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem0.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem0.CSDECODE_A = "0b000";
    defparam mem0.CSDECODE_B = "0b000";
    defparam mem0.GSR = "DISABLED";
    defparam mem0.INITVAL_00 = "0x1E8930828C0100410A93004B411A6308AF100025028930682004A731E028008600006F004600006F";
    defparam mem0.INITVAL_01 = "0x00AB701860000EF1F8E10021300200042170100000437080011029300200002B710A821C8B100604";
    defparam mem0.INITVAL_02 = "0x05C1D01A01102131C0511FC231088A108061C0C11EC23060200007314001054BD060451407300004";
    defparam mem0.INITVAL_03 = "0x100E701A01102131C0511FC231088A108061C0C11EC2306020000731C2C11E48306E0210226100A2";
    defparam mem0.INITVAL_04 = "0x000000000000000000000000000000000000000006020000731C2C11E48306E0210226100A200005";
    defparam mem0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_06 = "0x0000000422000000042200000004220000000422000000045400000004D400000002F800000002F8";
    defparam mem0.INITVAL_07 = "0x00000004220000000422000000042200000004220000000422000000042200000004220000000422";
    defparam mem0.INITVAL_08 = "0x10E931800110C131FCE71DAE300EC1000071C0231C80110E93000E61F2631CA0110E131C80110C93";
    defparam mem0.INITVAL_09 = "0x08690076E000E9312CB21800110E1300C91076E000C13134F111C911FEF710C93004F60EA6318241";
    defparam mem0.INITVAL_0A = "0x07A2000E131C60110E93000670FC631C801106131C60110E131FCD7136E31FCC705C2300E1100E91";
    defparam mem0.INITVAL_0B = "0x1802208C0102E2000A930188000A1302261100821FC671D4E300EC100E41000A71E023000070EA03";
    defparam mem0.INITVAL_0C = "0x00423010050CE931BEFD1061C000F70042313EE11FEF500E931C64114E031C60118A03044F518406";
    defparam mem0.INITVAL_0D = "0x088021C4F111023080920041000E93000E71286313EE100E8500EF000E131C60118E83040FD000F7";
    defparam mem0.INITVAL_0E = "0x1C64114C831A6F808E490100000EB71CC3E01EF000E930409D180060760000A13022711008200221";
    defparam mem0.INITVAL_0F = "0x16073000A512AB308A851400107EBD116F81C64114E8300006102231C64114C83114D808A0108E29";
    defparam mem0.INITVAL_10 = "0x06045060730100000A13060200007306A020604516073000A512AB308A85060200007306A0206845";
    defparam mem0.INITVAL_11 = "0x0080518A09102081082A184061802202261100820604516073000A512AB308A85000400006F10082";
    defparam mem0.INITVAL_12 = "0x1C226102040049500A6318001168831503D0022108A290809208802040A108A351FA6D1000805081";
    defparam mem0.INITVAL_13 = "0x0007306A02180A1144231D20110A13060200007306A02180A1144230009500E631DA011089300A05";
    defparam mem0.INITVAL_14 = "0x112881800116A830600616CF308CA11DA0110E13060200007306A0206045060730000800A3706020";
    defparam mem0.INITVAL_15 = "0x1D20110A9310082060061407306045140730000800AB7180B114023000B601C63000E511A6300A85";
    defparam mem0.INITVAL_16 = "0x10063008851D20110A93180811688317EE106006160731FCE601CE31804114E03060061407316EDD";
    defparam mem0.INITVAL_17 = "0x10893060200007306A02004B500A631820112A0318091148231FCB411EA3000A410C630CA8A004B4";
    defparam mem0.INITVAL_18 = "0x08A05060200007306A02000B500A631820112A0318091148231FCA511EA30CA0A1FCA410EE31CA01";
    defparam mem0.INITVAL_19 = "0x10488000D6010631808116C030600706E7308E211D20110A930AA7D060200007306A02180A111223";
    defparam mem0.INITVAL_1A = "0x16C03100820600704073180B114C231CA0110A93100820600704073180D114C23000B610E6300C85";
    defparam mem0.INITVAL_1B = "0x06047160730100000E9314A3E1E0000460307C8000E931008208A051008208A01000D60086318081";
    defparam mem0.INITVAL_1C = "0x1C84114E8306047160730100000E931008206047140731E0A0044231C8C1140231C8B11442312A1A";
    defparam mem0.INITVAL_1D = "0x00490000210C86C0E46F0EE200586F0D86C0CA48000001008210E821C801144231C80114A0318E91";
    defparam mem0.INITVAL_1E = "0x00000000000000001000008200000000021000000000300200004500020000450002000049000200";
    defparam mem0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INIT_DATA = "STATIC";
    FD1P3AX i3589 (.D(n5627), .SP(rom_buff_out_7__N_118), .CK(spi_clk_pos_derived_59), 
            .Q(n5690));
    defparam i3589.GSR = "DISABLED";
    DP16KD mem2 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n5643), .ADB4(n5638), 
           .ADB5(n5637), .ADB6(n5636), .ADB7(n5635), .ADB8(n5634), .ADB9(n5633), 
           .ADB10(n5632), .ADB11(n5631), .ADB12(n5630), .ADB13(n5629), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n5704), .DOB1(n5705), .DOB2(n5706), 
           .DOB3(n5707), .DOB4(n5708), .DOB5(n5709), .DOB6(n5710), .DOB7(n5711));
    defparam mem2.DATA_WIDTH_A = 9;
    defparam mem2.DATA_WIDTH_B = 9;
    defparam mem2.REGMODE_A = "NOREG";
    defparam mem2.REGMODE_B = "NOREG";
    defparam mem2.RESETMODE = "SYNC";
    defparam mem2.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem2.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem2.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem2.CSDECODE_A = "0b000";
    defparam mem2.CSDECODE_B = "0b000";
    defparam mem2.GSR = "DISABLED";
    defparam mem2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INIT_DATA = "STATIC";
    FD1P3AX i3607 (.D(n5644), .SP(rom_buff_out_7__N_118), .CK(spi_clk_pos_derived_59), 
            .Q(n5732));
    defparam i3607.GSR = "DISABLED";
    DP16KD mem3 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n5643), .ADB4(n5638), 
           .ADB5(n5637), .ADB6(n5636), .ADB7(n5635), .ADB8(n5634), .ADB9(n5633), 
           .ADB10(n5632), .ADB11(n5631), .ADB12(n5630), .ADB13(n5629), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n5724), .DOB1(n5725), .DOB2(n5726), 
           .DOB3(n5727), .DOB4(n5728), .DOB5(n5729), .DOB6(n5730), .DOB7(n5731));
    defparam mem3.DATA_WIDTH_A = 9;
    defparam mem3.DATA_WIDTH_B = 9;
    defparam mem3.REGMODE_A = "NOREG";
    defparam mem3.REGMODE_B = "NOREG";
    defparam mem3.RESETMODE = "SYNC";
    defparam mem3.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem3.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem3.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem3.CSDECODE_A = "0b000";
    defparam mem3.CSDECODE_B = "0b000";
    defparam mem3.GSR = "DISABLED";
    defparam mem3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INIT_DATA = "STATIC";
    DP16KD mem1 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n5643), .ADB4(n5638), 
           .ADB5(n5637), .ADB6(n5636), .ADB7(n5635), .ADB8(n5634), .ADB9(n5633), 
           .ADB10(n5632), .ADB11(n5631), .ADB12(n5630), .ADB13(n5629), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n5716), .DOB1(n5717), .DOB2(n5718), 
           .DOB3(n5719), .DOB4(n5720), .DOB5(n5721), .DOB6(n5722), .DOB7(n5723));
    defparam mem1.DATA_WIDTH_A = 9;
    defparam mem1.DATA_WIDTH_B = 9;
    defparam mem1.REGMODE_A = "NOREG";
    defparam mem1.REGMODE_B = "NOREG";
    defparam mem1.RESETMODE = "SYNC";
    defparam mem1.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem1.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem1.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem1.CSDECODE_A = "0b000";
    defparam mem1.CSDECODE_B = "0b000";
    defparam mem1.GSR = "DISABLED";
    defparam mem1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INIT_DATA = "STATIC";
    LUT4 i22427_3_lut (.A(n5722), .B(n5730), .C(n5732), .Z(n24770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22427_3_lut.init = 16'hcaca;
    LUT4 i22426_3_lut (.A(n5702), .B(n5710), .C(n5732), .Z(n24769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22426_3_lut.init = 16'hcaca;
    LUT4 i22424_3_lut (.A(n5723), .B(n5731), .C(n5732), .Z(n24767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22424_3_lut.init = 16'hcaca;
    LUT4 i22423_3_lut (.A(n5703), .B(n5711), .C(n5732), .Z(n24766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22423_3_lut.init = 16'hcaca;
    LUT4 i22418_3_lut (.A(n5720), .B(n5728), .C(n5732), .Z(n24761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22418_3_lut.init = 16'hcaca;
    LUT4 i22417_3_lut (.A(n5700), .B(n5708), .C(n5732), .Z(n24760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22417_3_lut.init = 16'hcaca;
    LUT4 i22373_3_lut (.A(n5721), .B(n5729), .C(n5732), .Z(n24716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22373_3_lut.init = 16'hcaca;
    LUT4 i22372_3_lut (.A(n5701), .B(n5709), .C(n5732), .Z(n24715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22372_3_lut.init = 16'hcaca;
    PFUMX i22374 (.BLUT(n24715), .ALUT(n24716), .C0(n5690), .Z(\rom_buff_out[5] ));
    PFUMX i22419 (.BLUT(n24760), .ALUT(n24761), .C0(n5690), .Z(\rom_buff_out[4] ));
    PFUMX i22425 (.BLUT(n24766), .ALUT(n24767), .C0(n5690), .Z(\rom_buff_out[7] ));
    PFUMX i22428 (.BLUT(n24769), .ALUT(n24770), .C0(n5690), .Z(\rom_buff_out[6] ));
    
endmodule
//
// Verilog Description of module \BRAM(ADDR_WIDTH=11) 
//

module \BRAM(ADDR_WIDTH=11)  (\addr[1] , \addr[2] , \addr[3] , \addr[4] , 
            \addr[5] , \addr[6] , \addr[7] , \addr[8] , \addr[9] , 
            \addr[10] , \addr[11] , n5643, n5638, n5637, n5636, 
            n5635, n5634, n5633, n5632, n5631, n5630, n5629, qspi_data_in_3__N_1, 
            data_buff_in, ram_b_buff_out, spi_clk_pos_derived_59, ram_b_buff_out_7__N_128, 
            ram_b_buff_out_7__N_131, GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input \addr[1] ;
    input \addr[2] ;
    input \addr[3] ;
    input \addr[4] ;
    input \addr[5] ;
    input \addr[6] ;
    input \addr[7] ;
    input \addr[8] ;
    input \addr[9] ;
    input \addr[10] ;
    input \addr[11] ;
    input n5643;
    input n5638;
    input n5637;
    input n5636;
    input n5635;
    input n5634;
    input n5633;
    input n5632;
    input n5631;
    input n5630;
    input n5629;
    input [3:0]qspi_data_in_3__N_1;
    input [3:0]data_buff_in;
    output [7:0]ram_b_buff_out;
    input spi_clk_pos_derived_59;
    input ram_b_buff_out_7__N_128;
    input ram_b_buff_out_7__N_131;
    input GND_net;
    input VCC_net;
    
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    DP16KD mem0 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(ram_b_buff_out_7__N_128), .CSA0(GND_net), .CSA1(GND_net), 
           .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
           .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
           .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), 
           .DIB10(GND_net), .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), 
           .DIB14(GND_net), .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), 
           .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(n5643), 
           .ADB4(n5638), .ADB5(n5637), .ADB6(n5636), .ADB7(n5635), .ADB8(n5634), 
           .ADB9(n5633), .ADB10(n5632), .ADB11(n5631), .ADB12(n5630), 
           .ADB13(n5629), .CEB(ram_b_buff_out_7__N_131), .OCEB(VCC_net), 
           .CLKB(spi_clk_pos_derived_59), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOB0(ram_b_buff_out[0]), 
           .DOB1(ram_b_buff_out[1]), .DOB2(ram_b_buff_out[2]), .DOB3(ram_b_buff_out[3]), 
           .DOB4(ram_b_buff_out[4]), .DOB5(ram_b_buff_out[5]), .DOB6(ram_b_buff_out[6]), 
           .DOB7(ram_b_buff_out[7]));
    defparam mem0.DATA_WIDTH_A = 9;
    defparam mem0.DATA_WIDTH_B = 9;
    defparam mem0.REGMODE_A = "NOREG";
    defparam mem0.REGMODE_B = "NOREG";
    defparam mem0.RESETMODE = "SYNC";
    defparam mem0.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem0.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem0.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem0.CSDECODE_A = "0b000";
    defparam mem0.CSDECODE_B = "0b000";
    defparam mem0.GSR = "DISABLED";
    defparam mem0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INIT_DATA = "STATIC";
    
endmodule
//
// Verilog Description of module \BRAM(ADDR_WIDTH=12) 
//

module \BRAM(ADDR_WIDTH=12)  (\addr[1] , \addr[2] , \addr[3] , \addr[4] , 
            \addr[5] , \addr[6] , \addr[7] , \addr[8] , \addr[9] , 
            \addr[10] , \addr[11] , n5643, n5638, n5637, n5636, 
            n5635, n5634, n5633, n5632, n5631, n5630, n5629, qspi_data_in_3__N_1, 
            data_buff_in, n5745, n5746, n5747, n5748, n5749, n5750, 
            n5751, n5752, spi_clk_pos_derived_59, n22126, ram_a_buff_out_7__N_127, 
            GND_net, VCC_net, n5753, n5644, n5737, n5738, n5739, 
            n5740, n5741, n5742, n5743, n5744, n22125) /* synthesis syn_module_defined=1 */ ;
    input \addr[1] ;
    input \addr[2] ;
    input \addr[3] ;
    input \addr[4] ;
    input \addr[5] ;
    input \addr[6] ;
    input \addr[7] ;
    input \addr[8] ;
    input \addr[9] ;
    input \addr[10] ;
    input \addr[11] ;
    input n5643;
    input n5638;
    input n5637;
    input n5636;
    input n5635;
    input n5634;
    input n5633;
    input n5632;
    input n5631;
    input n5630;
    input n5629;
    input [3:0]qspi_data_in_3__N_1;
    input [3:0]data_buff_in;
    output n5745;
    output n5746;
    output n5747;
    output n5748;
    output n5749;
    output n5750;
    output n5751;
    output n5752;
    input spi_clk_pos_derived_59;
    input n22126;
    input ram_a_buff_out_7__N_127;
    input GND_net;
    input VCC_net;
    output n5753;
    input n5644;
    output n5737;
    output n5738;
    output n5739;
    output n5740;
    output n5741;
    output n5742;
    output n5743;
    output n5744;
    input n22125;
    
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    DP16KD mem1 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(n22126), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n5643), .ADB4(n5638), 
           .ADB5(n5637), .ADB6(n5636), .ADB7(n5635), .ADB8(n5634), .ADB9(n5633), 
           .ADB10(n5632), .ADB11(n5631), .ADB12(n5630), .ADB13(n5629), 
           .CEB(ram_a_buff_out_7__N_127), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n5745), .DOB1(n5746), .DOB2(n5747), 
           .DOB3(n5748), .DOB4(n5749), .DOB5(n5750), .DOB6(n5751), .DOB7(n5752));
    defparam mem1.DATA_WIDTH_A = 9;
    defparam mem1.DATA_WIDTH_B = 9;
    defparam mem1.REGMODE_A = "NOREG";
    defparam mem1.REGMODE_B = "NOREG";
    defparam mem1.RESETMODE = "SYNC";
    defparam mem1.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem1.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem1.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem1.CSDECODE_A = "0b000";
    defparam mem1.CSDECODE_B = "0b000";
    defparam mem1.GSR = "DISABLED";
    defparam mem1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INIT_DATA = "STATIC";
    FD1P3AX i3614 (.D(n5644), .SP(ram_a_buff_out_7__N_127), .CK(spi_clk_pos_derived_59), 
            .Q(n5753));
    defparam i3614.GSR = "DISABLED";
    DP16KD mem0 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(n22125), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n5643), .ADB4(n5638), 
           .ADB5(n5637), .ADB6(n5636), .ADB7(n5635), .ADB8(n5634), .ADB9(n5633), 
           .ADB10(n5632), .ADB11(n5631), .ADB12(n5630), .ADB13(n5629), 
           .CEB(ram_a_buff_out_7__N_127), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n5737), .DOB1(n5738), .DOB2(n5739), 
           .DOB3(n5740), .DOB4(n5741), .DOB5(n5742), .DOB6(n5743), .DOB7(n5744));
    defparam mem0.DATA_WIDTH_A = 9;
    defparam mem0.DATA_WIDTH_B = 9;
    defparam mem0.REGMODE_A = "NOREG";
    defparam mem0.REGMODE_B = "NOREG";
    defparam mem0.RESETMODE = "SYNC";
    defparam mem0.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem0.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem0.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem0.CSDECODE_A = "0b000";
    defparam mem0.CSDECODE_B = "0b000";
    defparam mem0.GSR = "DISABLED";
    defparam mem0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INIT_DATA = "STATIC";
    
endmodule
