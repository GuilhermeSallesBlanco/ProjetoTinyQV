// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Thu Nov 20 15:56:30 2025
//
// Verilog Description of module tinyQV_top
//

module tinyQV_top (clk, rst_n, ui_in, uo_out) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(8[8:18])
    input clk;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    input rst_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(10[20:25])
    input [7:0]ui_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    output [7:0]uo_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_41 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    
    wire GND_net, VCC_net, rst_n_c, ui_in_c_1, ui_in_c_0, uo_out_c_6, 
        uo_out_c_5, uo_out_c_4, uo_out_c_3, uo_out_c_2, rst_reg_n, 
        n3597;
    wire [27:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    wire [31:0]data_to_write;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(56[17:30])
    wire [31:0]data_from_read;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(59[16:30])
    wire [3:0]debug_rd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(75[16:24])
    
    wire debug_uart_txd;
    wire [7:6]gpio_out_sel;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(79[16:28])
    
    wire debug_register_data;
    wire [3:0]debug_rd_r;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(85[15:25])
    
    wire peri_data_ready, read_en;
    wire [7:0]ui_in_sync0;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(101[15:26])
    wire [7:0]ui_in_sync;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(102[15:25])
    wire [7:0]time_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(222[15:25])
    wire [1:0]gpio_out_sel_7__N_9;
    
    wire debug_instr_valid;
    wire [1:0]qv_data_write_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(64[15:30])
    wire [1:0]qv_data_read_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(65[15:29])
    
    wire rst_reg_n_adj_2398, next_bit, uart_txd_N_2327, mem_op_increment_reg_de;
    wire [31:0]imm;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(100[16:19])
    wire [2:1]instr_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(113[15:24])
    
    wire mem_op_increment_reg;
    wire [31:0]pc;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(128[17:19])
    wire [31:0]next_pc_for_core;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(129[17:33])
    wire [4:2]counter_hi;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(139[15:25])
    wire [3:1]instr_write_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(152[15:33])
    wire [3:1]instr_avail_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(156[16:31])
    wire [23:1]early_branch_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[17:34])
    
    wire n6595, n18562, n6837, n47, n26, clk_c_enable_354, n22526, 
        clk_c_enable_27, n22518, n21541;
    wire [22:0]instr_addr_23__N_49;
    
    wire n20901, qspi_write_done, data_stall, n25151, n18561, n14111, 
        continue_txn_N_1862, data_stall_N_1889, n38, n39, n40, n41, 
        n42, n43, n44, n45, clk_c_enable_397, n25463;
    wire [31:0]next_fsm_state_3__N_2230;
    
    wire n2010, n20732, n17512, n17515, n1949, n1032, n2015, n1969, 
        n18560;
    wire [1:0]cycle;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(58[15:20])
    wire [3:0]mul_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(138[16:23])
    
    wire n8527, instr_complete_N_1378, n777, n18546, n18538, n18537, 
        n18545, n18559, n18544, clk_c_enable_208, n22334, n25419, 
        n25154, clk_c_enable_322, n25417, is_writing, is_writing_N_2062, 
        n18558, n23082, n18543, n18571, n18557, n18556, n8457, 
        n1092, n18555, n18542, n18536, n18570, n18541, n18535, 
        n8229, n18569, n18554, n18553, n18540, n18568, n18567, 
        n18552;
    wire [15:0]accum;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(104[22:27])
    wire [19:0]next_accum;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[23:33])
    wire [19:0]d_3__N_1599;
    
    wire n18566, n18551, n8146, n18565, n18532, n25371, n25370, 
        n18530, n20638, n18531, n18526, n18533, n18527, n18525, 
        n25363, n18529, n18528, n18548, n18539, clk_c_enable_206, 
        n18564, n25360, n18563, n18547, n23085, n23084, n25194, 
        n20728, n25321, n25320, n21746, n4, n25299, n20582, n22895, 
        n20097, n25464, n22788, n25276, n25273, n22728, n22726, 
        n20731, n25252, n24185, n25175, n24186;
    
    VHI i2 (.Z(VCC_net));
    INV i23149 (.A(clk_c), .Z(clk_N_41));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    FD1S3AX debug_rd_r_i0 (.D(debug_rd[0]), .CK(clk_c), .Q(debug_rd_r[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(241[12] 243[8])
    defparam debug_rd_r_i0.GSR = "DISABLED";
    FD1S3AX rst_reg_n_52 (.D(rst_n_c), .CK(clk_N_41), .Q(rst_reg_n));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(31[12:46])
    defparam rst_reg_n_52.GSR = "DISABLED";
    \uart_tx(BIT_RATE=1000000,CLK_HZ=14000000)  i_debug_uart_tx (.debug_uart_txd(debug_uart_txd), 
            .clk_c(clk_c), .n17515(n17515), .clk_c_enable_397(clk_c_enable_397), 
            .n25276(n25276), .rst_reg_n(rst_reg_n), .next_bit(next_bit), 
            .uart_txd_N_2327(uart_txd_N_2327), .n25360(n25360), .\data_to_write[7] (data_to_write[7]), 
            .\data_to_write[5] (data_to_write[5]), .\data_to_write[0] (data_to_write[0]), 
            .\data_to_write[6] (data_to_write[6]), .\data_to_write[1] (data_to_write[1]), 
            .\data_to_write[2] (data_to_write[2]), .\data_to_write[3] (data_to_write[3]), 
            .\data_to_write[4] (data_to_write[4])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(213[67] 220[6])
    CCU2C _add_1_4236_add_4_12 (.A0(imm[11]), .B0(pc[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[12]), .B1(pc[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18555), .COUT(n18556), .S0(early_branch_addr[11]), .S1(early_branch_addr[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_4233_add_4_5 (.A0(pc[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[7]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18540), .COUT(n18541), .S0(next_pc_for_core[6]), .S1(next_pc_for_core[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_5.INJECT1_1 = "NO";
    FD1S3IX time_count_3135__i0 (.D(n45), .CK(clk_c), .CD(n777), .Q(time_count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135__i0.GSR = "DISABLED";
    CCU2C _add_1_4236_add_4_10 (.A0(imm[9]), .B0(pc[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[10]), .B1(pc[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18554), .COUT(n18555), .S0(early_branch_addr[9]), .S1(early_branch_addr[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_4 (.A0(accum[2]), .B0(d_3__N_1599[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[3]), .B1(d_3__N_1599[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18525), .COUT(n18526), .S0(mul_out[2]), 
          .S1(mul_out[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_4.INJECT1_1 = "NO";
    FD1P3AX gpio_out_sel_i7 (.D(gpio_out_sel_7__N_9[1]), .SP(clk_c_enable_322), 
            .CK(clk_c), .Q(gpio_out_sel[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(204[12] 211[8])
    defparam gpio_out_sel_i7.GSR = "DISABLED";
    OB uo_out_pad_4 (.I(uo_out_c_4), .O(uo_out[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    LUT4 i3245_4_lut_then_3_lut (.A(n25273), .B(counter_hi[4]), .C(counter_hi[3]), 
         .Z(n25464)) /* synthesis lut_function=(A+!((C)+!B)) */ ;
    defparam i3245_4_lut_then_3_lut.init = 16'haeae;
    LUT4 i3245_4_lut_else_3_lut (.A(n25273), .B(counter_hi[4]), .C(counter_hi[3]), 
         .D(counter_hi[2]), .Z(n25463)) /* synthesis lut_function=(A+!((C+!(D))+!B)) */ ;
    defparam i3245_4_lut_else_3_lut.init = 16'haeaa;
    FD1S3AX ui_in_sync_i2 (.D(ui_in_sync0[1]), .CK(clk_c), .Q(ui_in_sync[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i2.GSR = "DISABLED";
    LUT4 gnd_bdd_2_lut_21962 (.A(n24185), .B(rst_reg_n_adj_2398), .Z(n24186)) /* synthesis lut_function=(A (B)) */ ;
    defparam gnd_bdd_2_lut_21962.init = 16'h8888;
    LUT4 i20992_2_lut_rep_458_4_lut (.A(pc[2]), .B(n25363), .C(debug_instr_valid), 
         .D(n3597), .Z(n25194)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i20992_2_lut_rep_458_4_lut.init = 16'h0035;
    IB ui_in_pad_0 (.I(ui_in[0]), .O(ui_in_c_0));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_1 (.I(ui_in[1]), .O(ui_in_c_1));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB rst_n_pad (.I(rst_n), .O(rst_n_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(10[20:25])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    OB uo_out_pad_0 (.I(GND_net), .O(uo_out[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_1 (.I(GND_net), .O(uo_out[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_2 (.I(uo_out_c_2), .O(uo_out[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_3 (.I(uo_out_c_3), .O(uo_out[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    LUT4 i11899_2_lut_rep_585_3_lut_4_lut (.A(n25370), .B(n17512), .C(qspi_write_done), 
         .D(n25371), .Z(n25321)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11899_2_lut_rep_585_3_lut_4_lut.init = 16'hfffe;
    LUT4 i4425_2_lut_rep_584_3_lut_4_lut (.A(n25370), .B(n17512), .C(qspi_write_done), 
         .D(n25371), .Z(n25320)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;
    defparam i4425_2_lut_rep_584_3_lut_4_lut.init = 16'hfff1;
    FD1S3AX ui_in_sync0_i2 (.D(ui_in_c_1), .CK(clk_c), .Q(ui_in_sync0[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i2.GSR = "DISABLED";
    OB uo_out_pad_5 (.I(uo_out_c_5), .O(uo_out[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    FD1S3AX ui_in_sync0_i1 (.D(ui_in_c_0), .CK(clk_c), .Q(ui_in_sync0[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i1.GSR = "DISABLED";
    CCU2C _add_1_4236_add_4_8 (.A0(imm[7]), .B0(pc[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[8]), .B1(pc[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18553), .COUT(n18554), .S0(early_branch_addr[7]), .S1(early_branch_addr[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_8.INJECT1_1 = "NO";
    LUT4 i11667_4_lut (.A(n25360), .B(data_from_read[2]), .C(n25299), 
         .D(addr[4]), .Z(data_from_read[0])) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i11667_4_lut.init = 16'heccc;
    LUT4 i11948_3_lut (.A(gpio_out_sel[6]), .B(data_from_read[2]), .C(n8229), 
         .Z(data_from_read[6])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i11948_3_lut.init = 16'hecec;
    FD1P3AX debug_register_data_57 (.D(n6837), .SP(clk_c_enable_208), .CK(clk_c), 
            .Q(debug_register_data));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(234[12] 239[8])
    defparam debug_register_data_57.GSR = "DISABLED";
    OB uo_out_pad_6 (.I(uo_out_c_6), .O(uo_out[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    FD1S3AX debug_rd_r_i3 (.D(debug_rd[3]), .CK(clk_c), .Q(debug_rd_r[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(241[12] 243[8])
    defparam debug_rd_r_i3.GSR = "DISABLED";
    FD1S3AX debug_rd_r_i2 (.D(debug_rd[2]), .CK(clk_c), .Q(debug_rd_r[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(241[12] 243[8])
    defparam debug_rd_r_i2.GSR = "DISABLED";
    FD1S3AX debug_rd_r_i1 (.D(debug_rd[1]), .CK(clk_c), .Q(debug_rd_r[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(241[12] 243[8])
    defparam debug_rd_r_i1.GSR = "DISABLED";
    OB uo_out_pad_7 (.I(GND_net), .O(uo_out[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    LUT4 i22_4_lut (.A(n20901), .B(n8457), .C(n47), .D(n20728), .Z(data_from_read[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i22_4_lut.init = 16'hcacf;
    LUT4 i18748_2_lut (.A(addr[5]), .B(addr[4]), .Z(n20901)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i18748_2_lut.init = 16'h2222;
    CCU2C _add_1_4233_add_4_3 (.A0(pc[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[5]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18539), .COUT(n18540), .S0(next_pc_for_core[4]), .S1(next_pc_for_core[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_20 (.A0(d_3__N_1599[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_3__N_1599[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18533), .S0(next_accum[18]), .S1(next_accum[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_add_4_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_add_4_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_18 (.A0(d_3__N_1599[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_3__N_1599[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18532), .COUT(n18533), .S0(next_accum[16]), 
          .S1(next_accum[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_add_4_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_add_4_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_18.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n22526), .B(n8457), .C(n22518), .D(addr[8]), .Z(n47)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_464 (.A(addr[7]), .B(addr[9]), .C(addr[6]), .D(addr[10]), 
         .Z(n22526)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_4_lut_adj_464.init = 16'hfffe;
    LUT4 i1_2_lut (.A(addr[0]), .B(addr[1]), .Z(n22518)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i1_2_lut.init = 16'heeee;
    FD1S3IX time_count_3135__i1 (.D(n44), .CK(clk_c), .CD(n777), .Q(time_count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135__i1.GSR = "DISABLED";
    VLO i1 (.Z(GND_net));
    LUT4 i11445_2_lut (.A(debug_rd_r[0]), .B(debug_register_data), .Z(uo_out_c_2)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(154[24:73])
    defparam i11445_2_lut.init = 16'h8888;
    FD1S3IX time_count_3135__i2 (.D(n43), .CK(clk_c), .CD(n777), .Q(time_count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135__i2.GSR = "DISABLED";
    FD1S3IX time_count_3135__i3 (.D(n42), .CK(clk_c), .CD(n777), .Q(time_count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135__i3.GSR = "DISABLED";
    FD1S3IX time_count_3135__i4 (.D(n41), .CK(clk_c), .CD(n777), .Q(time_count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135__i4.GSR = "DISABLED";
    FD1S3IX time_count_3135__i5 (.D(n40), .CK(clk_c), .CD(n777), .Q(time_count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135__i5.GSR = "DISABLED";
    FD1S3IX time_count_3135__i6 (.D(n39), .CK(clk_c), .CD(n777), .Q(time_count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135__i6.GSR = "DISABLED";
    FD1S3IX time_count_3135__i7 (.D(n38), .CK(clk_c), .CD(n777), .Q(time_count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135__i7.GSR = "DISABLED";
    LUT4 i1270_4_lut (.A(pc[2]), .B(n2010), .C(debug_instr_valid), .D(pc[1]), 
         .Z(n1969)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i1270_4_lut.init = 16'hcac0;
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i1275_4_lut (.A(pc[2]), .B(n2015), .C(debug_instr_valid), .D(pc[1]), 
         .Z(n1949)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i1275_4_lut.init = 16'hc5c0;
    LUT4 rst_reg_n_bdd_4_lut (.A(cycle[0]), .B(n14111), .C(clk_c_enable_206), 
         .D(instr_complete_N_1378), .Z(n24185)) /* synthesis lut_function=(!(A (B (C))+!A (((D)+!C)+!B))) */ ;
    defparam rst_reg_n_bdd_4_lut.init = 16'h2a6a;
    FD1P3IX gpio_out_sel_i6 (.D(data_to_write[6]), .SP(clk_c_enable_322), 
            .CD(n20097), .CK(clk_c), .Q(gpio_out_sel[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(204[12] 211[8])
    defparam gpio_out_sel_i6.GSR = "DISABLED";
    FD1S3AX ui_in_sync_i1 (.D(ui_in_sync0[0]), .CK(clk_c), .Q(next_fsm_state_3__N_2230[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i1.GSR = "DISABLED";
    LUT4 i1_3_lut (.A(addr[2]), .B(n47), .C(addr[4]), .Z(n20638)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut.init = 16'h1010;
    LUT4 i222_2_lut_rep_516_4_lut (.A(n25299), .B(n20638), .C(n20582), 
         .D(n25360), .Z(n25252)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(183[13:50])
    defparam i222_2_lut_rep_516_4_lut.init = 16'h0080;
    CCU2C _add_1_4233_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[3]), .B1(n25419), .C1(instr_len[2]), 
          .D1(pc[2]), .COUT(n18539), .S1(next_pc_for_core[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_4233_add_4_1.INIT1 = 16'h566a;
    defparam _add_1_4233_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_22 (.A0(pc[23]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18571), .S0(instr_addr_23__N_49[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_22.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_22.INIT1 = 16'h0000;
    defparam _add_1_4241_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_22.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_20 (.A0(pc[21]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[22]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18570), .COUT(n18571));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_20.INJECT1_1 = "NO";
    CCU2C time_count_3135_add_4_9 (.A0(time_count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18538), .S0(n38));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135_add_4_9.INIT0 = 16'haaa0;
    defparam time_count_3135_add_4_9.INIT1 = 16'h0000;
    defparam time_count_3135_add_4_9.INJECT1_0 = "NO";
    defparam time_count_3135_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_4236_add_4_6 (.A0(imm[5]), .B0(pc[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[6]), .B1(pc[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18552), .COUT(n18553), .S0(early_branch_addr[5]), .S1(early_branch_addr[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_6.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_465 (.A(qv_data_write_n[0]), .B(n20731), .C(qv_data_read_n[0]), 
         .Z(n20732)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_adj_465.init = 16'hecec;
    GSR GSR_INST (.GSR(rst_reg_n));
    CCU2C _add_1_4241_add_4_18 (.A0(pc[19]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[20]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18569), .COUT(n18570));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_16 (.A0(pc[17]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[18]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18568), .COUT(n18569));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_16.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_16.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_14 (.A0(pc[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[16]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18567), .COUT(n18568));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_14.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_14.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_4236_add_4_4 (.A0(imm[3]), .B0(pc[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[4]), .B1(pc[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18551), .COUT(n18552), .S0(early_branch_addr[3]), .S1(early_branch_addr[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_4.INJECT1_1 = "NO";
    CCU2C time_count_3135_add_4_7 (.A0(time_count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18537), .COUT(n18538), .S0(n40), .S1(n39));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135_add_4_7.INIT0 = 16'haaa0;
    defparam time_count_3135_add_4_7.INIT1 = 16'haaa0;
    defparam time_count_3135_add_4_7.INJECT1_0 = "NO";
    defparam time_count_3135_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_12 (.A0(pc[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[14]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18566), .COUT(n18567));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_12.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_12.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_4236_add_4_2 (.A0(imm[1]), .B0(pc[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[2]), .B1(pc[2]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n18551), .S1(early_branch_addr[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_4236_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_10 (.A0(pc[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[12]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18565), .COUT(n18566));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_10.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_10.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_4233_add_4_21 (.A0(pc[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[23]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18548), .S0(next_pc_for_core[22]), .S1(next_pc_for_core[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_21.INJECT1_1 = "NO";
    CCU2C time_count_3135_add_4_5 (.A0(time_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18536), .COUT(n18537), .S0(n42), .S1(n41));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135_add_4_5.INIT0 = 16'haaa0;
    defparam time_count_3135_add_4_5.INIT1 = 16'haaa0;
    defparam time_count_3135_add_4_5.INJECT1_0 = "NO";
    defparam time_count_3135_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_16 (.A0(accum[14]), .B0(d_3__N_1599[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[15]), .B1(d_3__N_1599[15]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18531), .COUT(n18532), .S0(next_accum[14]), 
          .S1(next_accum[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_16.INJECT1_1 = "NO";
    CCU2C time_count_3135_add_4_3 (.A0(time_count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18535), .COUT(n18536), .S0(n44), .S1(n43));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135_add_4_3.INIT0 = 16'haaa0;
    defparam time_count_3135_add_4_3.INIT1 = 16'haaa0;
    defparam time_count_3135_add_4_3.INJECT1_0 = "NO";
    defparam time_count_3135_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_6 (.A0(accum[4]), .B0(d_3__N_1599[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[5]), .B1(d_3__N_1599[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18526), .COUT(n18527), .S0(next_accum[4]), 
          .S1(next_accum[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_8 (.A0(pc[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[10]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18564), .COUT(n18565));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_8.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_8.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_4233_add_4_19 (.A0(pc[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[21]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18547), .COUT(n18548), .S0(next_pc_for_core[20]), .S1(next_pc_for_core[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_19.INJECT1_1 = "NO";
    LUT4 i20807_4_lut (.A(is_writing), .B(is_writing_N_2062), .C(n6595), 
         .D(n25151), .Z(n23082)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i20807_4_lut.init = 16'hcaaa;
    CCU2C _add_1_4233_add_4_17 (.A0(pc[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[19]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18546), .COUT(n18547), .S0(next_pc_for_core[18]), .S1(next_pc_for_core[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_17.INJECT1_1 = "NO";
    CCU2C time_count_3135_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n18535), .S1(n45));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[32:46])
    defparam time_count_3135_add_4_1.INIT0 = 16'h0000;
    defparam time_count_3135_add_4_1.INIT1 = 16'h555f;
    defparam time_count_3135_add_4_1.INJECT1_0 = "NO";
    defparam time_count_3135_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_6 (.A0(pc[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18563), .COUT(n18564));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_6.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_6.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_4233_add_4_15 (.A0(pc[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18545), .COUT(n18546), .S0(next_pc_for_core[16]), .S1(next_pc_for_core[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_4 (.A0(pc[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18562), .COUT(n18563));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_4.INIT0 = 16'haaa0;
    defparam _add_1_4241_add_4_4.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_4241_add_4_2 (.A0(instr_write_offset[3]), .B0(pc[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n18562));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_4241_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_4241_add_4_2.INIT1 = 16'haaa0;
    defparam _add_1_4241_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_4241_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_4236_add_4_24 (.A0(imm[23]), .B0(pc[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n18561), .S0(early_branch_addr[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_24.INIT1 = 16'h0000;
    defparam _add_1_4236_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_4233_add_4_13 (.A0(pc[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[15]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18544), .COUT(n18545), .S0(next_pc_for_core[14]), .S1(next_pc_for_core[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_4233_add_4_11 (.A0(pc[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[13]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18543), .COUT(n18544), .S0(next_pc_for_core[12]), .S1(next_pc_for_core[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_14 (.A0(accum[12]), .B0(d_3__N_1599[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[13]), .B1(d_3__N_1599[13]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18530), .COUT(n18531), .S0(next_accum[12]), 
          .S1(next_accum[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_2 (.A0(accum[0]), .B0(d_3__N_1599[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[1]), .B1(d_3__N_1599[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n18525), .S1(mul_out[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_add_4_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_10 (.A0(accum[8]), .B0(d_3__N_1599[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[9]), .B1(d_3__N_1599[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18528), .COUT(n18529), .S0(next_accum[8]), 
          .S1(next_accum[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_8 (.A0(accum[6]), .B0(d_3__N_1599[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[7]), .B1(d_3__N_1599[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18527), .COUT(n18528), .S0(next_accum[6]), 
          .S1(next_accum[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_12 (.A0(accum[10]), .B0(d_3__N_1599[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[11]), .B1(d_3__N_1599[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n18529), .COUT(n18530), .S0(next_accum[10]), 
          .S1(next_accum[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_4233_add_4_9 (.A0(pc[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[11]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18542), .COUT(n18543), .S0(next_pc_for_core[10]), .S1(next_pc_for_core[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_4236_add_4_22 (.A0(imm[21]), .B0(pc[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[22]), .B1(pc[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18560), .COUT(n18561), .S0(early_branch_addr[21]), .S1(early_branch_addr[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_22.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_681 (.A(addr[4]), .B(addr[5]), .Z(n25417)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_681.init = 16'heeee;
    CCU2C _add_1_4236_add_4_20 (.A0(imm[19]), .B0(pc[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[20]), .B1(pc[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18559), .COUT(n18560), .S0(early_branch_addr[19]), .S1(early_branch_addr[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_20.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(addr[4]), .B(addr[5]), .C(n47), .D(n8457), 
         .Z(n8229)) /* synthesis lut_function=(A (D)+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff01;
    CCU2C _add_1_4236_add_4_18 (.A0(imm[17]), .B0(pc[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[18]), .B1(pc[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18558), .COUT(n18559), .S0(early_branch_addr[17]), .S1(early_branch_addr[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_18.INJECT1_1 = "NO";
    LUT4 i21720_2_lut (.A(n8527), .B(rst_reg_n), .Z(n777)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i21720_2_lut.init = 16'h7777;
    LUT4 i1_4_lut_adj_466 (.A(n22728), .B(n22895), .C(time_count[0]), 
         .D(n22726), .Z(n8527)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_466.init = 16'hffbf;
    LUT4 i1_3_lut_adj_467 (.A(time_count[4]), .B(time_count[7]), .C(time_count[6]), 
         .Z(n22728)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_467.init = 16'hfefe;
    LUT4 i20681_2_lut (.A(time_count[2]), .B(time_count[3]), .Z(n22895)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20681_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_468 (.A(time_count[5]), .B(time_count[1]), .Z(n22726)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_468.init = 16'heeee;
    CCU2C _add_1_4233_add_4_7 (.A0(pc[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[9]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18541), .COUT(n18542), .S0(next_pc_for_core[8]), .S1(next_pc_for_core[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_4233_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_4233_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_4233_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_4233_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_4236_add_4_16 (.A0(imm[15]), .B0(pc[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[16]), .B1(pc[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18557), .COUT(n18558), .S0(early_branch_addr[15]), .S1(early_branch_addr[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_4236_add_4_14 (.A0(imm[13]), .B0(pc[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[14]), .B1(pc[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n18556), .COUT(n18557), .S0(early_branch_addr[13]), .S1(early_branch_addr[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_4236_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_4236_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_4236_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_4236_add_4_14.INJECT1_1 = "NO";
    LUT4 mux_33_i2_3_lut (.A(ui_in_c_0), .B(data_to_write[7]), .C(n4), 
         .Z(gpio_out_sel_7__N_9[1])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(209[13:93])
    defparam mux_33_i2_3_lut.init = 16'hc5c5;
    LUT4 i1_4_lut_adj_469 (.A(n20582), .B(n47), .C(n25417), .D(addr[2]), 
         .Z(n4)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_469.init = 16'h0200;
    LUT4 i11447_2_lut (.A(debug_rd_r[2]), .B(debug_register_data), .Z(uo_out_c_4)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(156[24:73])
    defparam i11447_2_lut.init = 16'h8888;
    LUT4 i3254_4_lut (.A(n21746), .B(n25154), .C(n26), .D(n1032), .Z(clk_c_enable_354)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C))) */ ;
    defparam i3254_4_lut.init = 16'hfcdc;
    LUT4 i11446_2_lut (.A(debug_rd_r[1]), .B(debug_register_data), .Z(uo_out_c_3)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(155[24:73])
    defparam i11446_2_lut.init = 16'h8888;
    LUT4 i21765_2_lut_rep_563 (.A(n47), .B(addr[5]), .Z(n25299)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21765_2_lut_rep_563.init = 16'h1111;
    LUT4 i1_3_lut_rep_540_4_lut (.A(n47), .B(addr[5]), .C(n20582), .D(n20638), 
         .Z(n25276)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_rep_540_4_lut.init = 16'h1000;
    LUT4 i11448_2_lut (.A(debug_rd_r[3]), .B(debug_register_data), .Z(uo_out_c_5)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(157[24:73])
    defparam i11448_2_lut.init = 16'h8888;
    \peripherals_min(CLOCK_MHZ=14)  i_peripherals (.peri_data_ready(peri_data_ready), 
            .clk_c(clk_c), .n17515(n17515), .read_en(read_en)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(161[46] 180[6])
    LUT4 i20810_3_lut (.A(data_stall), .B(data_stall_N_1889), .C(continue_txn_N_1862), 
         .Z(n23085)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam i20810_3_lut.init = 16'hcece;
    LUT4 i1_2_lut_adj_470 (.A(addr[3]), .B(addr[5]), .Z(n22788)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(64[15:30])
    defparam i1_2_lut_adj_470.init = 16'h4444;
    LUT4 i4622_3_lut (.A(ui_in_c_1), .B(data_to_write[0]), .C(rst_reg_n), 
         .Z(n6837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(234[12] 239[8])
    defparam i4622_3_lut.init = 16'hcaca;
    LUT4 i11450_2_lut (.A(debug_uart_txd), .B(gpio_out_sel[6]), .Z(uo_out_c_6)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(158[24:70])
    defparam i11450_2_lut.init = 16'h2222;
    LUT4 i20809_4_lut (.A(mem_op_increment_reg), .B(mem_op_increment_reg_de), 
         .C(n22334), .D(n25175), .Z(n23084)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i20809_4_lut.init = 16'hcaaa;
    LUT4 i21835_2_lut (.A(rst_reg_n), .B(n4), .Z(n20097)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21835_2_lut.init = 16'h1111;
    tinyQV i_tinyqv (.rst_reg_n_adj_10(rst_reg_n_adj_2398), .clk_c(clk_c), 
           .rst_reg_n(rst_reg_n), .peri_data_ready(peri_data_ready), .n25370(n25370), 
           .n8457(n8457), .n47(n47), .n20728(n20728), .\addr[2] (addr[2]), 
           .\addr[3] (addr[3]), .counter_hi({counter_hi}), .n17512(n17512), 
           .n20731(n20731), .n20732(n20732), .qspi_write_done(qspi_write_done), 
           .data_stall_N_1889(data_stall_N_1889), .data_stall(data_stall), 
           .n17515(n17515), .n25321(n25321), .is_writing_N_2062(is_writing_N_2062), 
           .n23085(n23085), .n25151(n25151), .data_to_write({Open_0, Open_1, 
           Open_2, Open_3, Open_4, Open_5, Open_6, Open_7, Open_8, 
           Open_9, Open_10, Open_11, Open_12, Open_13, Open_14, 
           Open_15, Open_16, Open_17, Open_18, Open_19, Open_20, 
           Open_21, Open_22, Open_23, Open_24, Open_25, Open_26, 
           Open_27, Open_28, Open_29, Open_30, data_to_write[0]}), 
           .is_writing(is_writing), .\data_to_write[7] (data_to_write[7]), 
           .\data_to_write[6] (data_to_write[6]), .\data_to_write[5] (data_to_write[5]), 
           .\data_to_write[4] (data_to_write[4]), .\data_to_write[3] (data_to_write[3]), 
           .\data_to_write[2] (data_to_write[2]), .\data_to_write[1] (data_to_write[1]), 
           .continue_txn_N_1862(continue_txn_N_1862), .n25320(n25320), .n25371(n25371), 
           .n1032(n1032), .n25154(n25154), .n23082(n23082), .n21746(n21746), 
           .clk_c_enable_354(clk_c_enable_354), .n6595(n6595), .next_bit(next_bit), 
           .n25252(n25252), .uart_txd_N_2327(uart_txd_N_2327), .clk_c_enable_397(clk_c_enable_397), 
           .n22788(n22788), .n20638(n20638), .clk_c_enable_208(clk_c_enable_208), 
           .n4(n4), .clk_c_enable_322(clk_c_enable_322), .n26(n26), .\pc[10] (pc[10]), 
           .\pc[11] (pc[11]), .\qv_data_read_n[0] (qv_data_read_n[0]), .\pc[12] (pc[12]), 
           .VCC_net(VCC_net), .debug_instr_valid(debug_instr_valid), .\pc[13] (pc[13]), 
           .\instr_len[2] (instr_len[2]), .\pc[14] (pc[14]), .\pc[1] (pc[1]), 
           .\addr[0] (addr[0]), .\pc[2] (pc[2]), .\pc[3] (pc[3]), .\pc[4] (pc[4]), 
           .\pc[5] (pc[5]), .\pc[6] (pc[6]), .\pc[7] (pc[7]), .\instr_write_offset[3] (instr_write_offset[3]), 
           .n25175(n25175), .n2015(n2015), .n2010(n2010), .\data_from_read[2] (data_from_read[2]), 
           .n8229(n8229), .\gpio_out_sel[7] (gpio_out_sel[7]), .n1949(n1949), 
           .n1969(n1969), .instr_complete_N_1378(instr_complete_N_1378), 
           .n21541(n21541), .n8146(n8146), .n3597(n3597), .\pc[15] (pc[15]), 
           .\qv_data_write_n[0] (qv_data_write_n[0]), .\pc[16] (pc[16]), 
           .\pc[17] (pc[17]), .\next_pc_for_core[3] (next_pc_for_core[3]), 
           .\next_pc_for_core[7] (next_pc_for_core[7]), .\pc[18] (pc[18]), 
           .\imm[19] (imm[19]), .\imm[23] (imm[23]), .\imm[11] (imm[11]), 
           .\imm[15] (imm[15]), .\imm[3] (imm[3]), .\imm[7] (imm[7]), 
           .\imm[18] (imm[18]), .\imm[22] (imm[22]), .n25363(n25363), 
           .\imm[10] (imm[10]), .\imm[14] (imm[14]), .\imm[2] (imm[2]), 
           .\imm[6] (imm[6]), .\imm[17] (imm[17]), .\imm[21] (imm[21]), 
           .\imm[9] (imm[9]), .\imm[13] (imm[13]), .\imm[1] (imm[1]), 
           .\imm[5] (imm[5]), .mem_op_increment_reg(mem_op_increment_reg), 
           .n23084(n23084), .\imm[16] (imm[16]), .\imm[20] (imm[20]), 
           .\imm[8] (imm[8]), .\imm[12] (imm[12]), .\imm[4] (imm[4]), 
           .\next_pc_for_core[4] (next_pc_for_core[4]), .\pc[9] (pc[9]), 
           .\next_pc_for_core[9] (next_pc_for_core[9]), .\next_pc_for_core[13] (next_pc_for_core[13]), 
           .\pc[19] (pc[19]), .\addr[4] (addr[4]), .\addr[5] (addr[5]), 
           .\pc[20] (pc[20]), .\pc[8] (pc[8]), .\instr_avail_len[3] (instr_avail_len[3]), 
           .\next_pc_for_core[8] (next_pc_for_core[8]), .\next_pc_for_core[12] (next_pc_for_core[12]), 
           .\addr[1] (addr[1]), .\addr[6] (addr[6]), .\addr[7] (addr[7]), 
           .\addr[8] (addr[8]), .\addr[9] (addr[9]), .\addr[10] (addr[10]), 
           .n25194(n25194), .clk_c_enable_206(clk_c_enable_206), .\next_pc_for_core[5] (next_pc_for_core[5]), 
           .\next_pc_for_core[6] (next_pc_for_core[6]), .\next_pc_for_core[10] (next_pc_for_core[10]), 
           .\next_pc_for_core[11] (next_pc_for_core[11]), .n25417(n25417), 
           .\next_pc_for_core[14] (next_pc_for_core[14]), .\next_pc_for_core[15] (next_pc_for_core[15]), 
           .\next_pc_for_core[16] (next_pc_for_core[16]), .\next_pc_for_core[17] (next_pc_for_core[17]), 
           .\next_pc_for_core[18] (next_pc_for_core[18]), .\next_pc_for_core[19] (next_pc_for_core[19]), 
           .\next_pc_for_core[20] (next_pc_for_core[20]), .\next_pc_for_core[21] (next_pc_for_core[21]), 
           .\next_pc_for_core[22] (next_pc_for_core[22]), .\pc[21] (pc[21]), 
           .\pc[22] (pc[22]), .\pc[23] (pc[23]), .\next_pc_for_core[23] (next_pc_for_core[23]), 
           .n25419(n25419), .n20582(n20582), .read_en(read_en), .\instr_addr_23__N_49[22] (instr_addr_23__N_49[22]), 
           .\early_branch_addr[23] (early_branch_addr[23]), .\early_branch_addr[5] (early_branch_addr[5]), 
           .\early_branch_addr[4] (early_branch_addr[4]), .\early_branch_addr[2] (early_branch_addr[2]), 
           .\early_branch_addr[6] (early_branch_addr[6]), .\early_branch_addr[3] (early_branch_addr[3]), 
           .\early_branch_addr[7] (early_branch_addr[7]), .\early_branch_addr[8] (early_branch_addr[8]), 
           .\early_branch_addr[9] (early_branch_addr[9]), .\early_branch_addr[10] (early_branch_addr[10]), 
           .\early_branch_addr[11] (early_branch_addr[11]), .\early_branch_addr[12] (early_branch_addr[12]), 
           .\early_branch_addr[13] (early_branch_addr[13]), .\early_branch_addr[14] (early_branch_addr[14]), 
           .\early_branch_addr[15] (early_branch_addr[15]), .\early_branch_addr[16] (early_branch_addr[16]), 
           .\early_branch_addr[17] (early_branch_addr[17]), .\early_branch_addr[18] (early_branch_addr[18]), 
           .\early_branch_addr[19] (early_branch_addr[19]), .\early_branch_addr[20] (early_branch_addr[20]), 
           .\early_branch_addr[21] (early_branch_addr[21]), .\early_branch_addr[22] (early_branch_addr[22]), 
           .n8527(n8527), .n22334(n22334), .\data_from_read[6] (data_from_read[6]), 
           .\data_from_read[0] (data_from_read[0]), .mem_op_increment_reg_de(mem_op_increment_reg_de), 
           .n25273(n25273), .clk_c_enable_27(clk_c_enable_27), .\next_fsm_state_3__N_2230[3] (next_fsm_state_3__N_2230[3]), 
           .\cycle[0] (cycle[0]), .\ui_in_sync[1] (ui_in_sync[1]), .n1092(n1092), 
           .debug_rd({debug_rd}), .accum({accum}), .d_3__N_1599({d_3__N_1599}), 
           .\mul_out[1] (mul_out[1]), .\mul_out[3] (mul_out[3]), .n14111(n14111), 
           .n24186(n24186), .\mul_out[2] (mul_out[2]), .\next_accum[6] (next_accum[6]), 
           .\next_accum[7] (next_accum[7]), .\next_accum[8] (next_accum[8]), 
           .\next_accum[9] (next_accum[9]), .\next_accum[10] (next_accum[10]), 
           .\next_accum[11] (next_accum[11]), .\next_accum[12] (next_accum[12]), 
           .\next_accum[13] (next_accum[13]), .\next_accum[14] (next_accum[14]), 
           .\next_accum[15] (next_accum[15]), .GND_net(GND_net), .\next_accum[16] (next_accum[16]), 
           .\next_accum[17] (next_accum[17]), .\next_accum[18] (next_accum[18]), 
           .\next_accum[19] (next_accum[19]), .\next_accum[5] (next_accum[5]), 
           .\next_accum[4] (next_accum[4])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(111[12] 150[6])
    PFUMX mux_3157_i3 (.BLUT(n8146), .ALUT(n21541), .C0(debug_instr_valid), 
          .Z(instr_avail_len[3]));
    PFUMX i22539 (.BLUT(n25463), .ALUT(n25464), .C0(n1092), .Z(clk_c_enable_27));
    
endmodule
//
// Verilog Description of module \uart_tx(BIT_RATE=1000000,CLK_HZ=14000000) 
//

module \uart_tx(BIT_RATE=1000000,CLK_HZ=14000000)  (debug_uart_txd, clk_c, 
            n17515, clk_c_enable_397, n25276, rst_reg_n, next_bit, 
            uart_txd_N_2327, n25360, \data_to_write[7] , \data_to_write[5] , 
            \data_to_write[0] , \data_to_write[6] , \data_to_write[1] , 
            \data_to_write[2] , \data_to_write[3] , \data_to_write[4] ) /* synthesis syn_module_defined=1 */ ;
    output debug_uart_txd;
    input clk_c;
    input n17515;
    input clk_c_enable_397;
    input n25276;
    input rst_reg_n;
    output next_bit;
    output uart_txd_N_2327;
    output n25360;
    input \data_to_write[7] ;
    input \data_to_write[5] ;
    input \data_to_write[0] ;
    input \data_to_write[6] ;
    input \data_to_write[1] ;
    input \data_to_write[2] ;
    input \data_to_write[3] ;
    input \data_to_write[4] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire uart_txd_N_2325;
    wire [7:0]data_to_send;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(51[24:36])
    wire [7:0]data_to_send_7__N_2305;
    wire [4:0]cycle_counter;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(55[25:38])
    
    wire n25332;
    wire [4:0]n18;
    
    wire n21431;
    wire [3:0]fsm_state;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(59[11:20])
    
    wire clk_c_enable_108, n25242, n25462, clk_c_enable_175;
    wire [4:0]n50;
    
    wire n24202, n25391, n25416, n6894, n22810;
    wire [3:0]n122;
    
    wire n24203;
    
    FD1S3JX txd_reg_46 (.D(uart_txd_N_2325), .CK(clk_c), .PD(n17515), 
            .Q(debug_uart_txd)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(135[8] 145[4])
    defparam txd_reg_46.GSR = "DISABLED";
    FD1P3IX data_to_send__i5 (.D(data_to_send_7__N_2305[5]), .SP(clk_c_enable_397), 
            .CD(n17515), .CK(clk_c), .Q(data_to_send[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i5.GSR = "DISABLED";
    FD1S3IX cycle_counter__i0 (.D(n18[0]), .CK(clk_c), .CD(n25332), .Q(cycle_counter[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i0.GSR = "DISABLED";
    FD1P3IX data_to_send__i6 (.D(data_to_send_7__N_2305[6]), .SP(clk_c_enable_397), 
            .CD(n17515), .CK(clk_c), .Q(data_to_send[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i6.GSR = "DISABLED";
    FD1P3AX data_to_send__i7 (.D(n21431), .SP(clk_c_enable_397), .CK(clk_c), 
            .Q(data_to_send[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i7.GSR = "DISABLED";
    FD1P3IX fsm_state__i0 (.D(n25462), .SP(clk_c_enable_108), .CD(n25242), 
            .CK(clk_c), .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam fsm_state__i0.GSR = "DISABLED";
    FD1P3IX cycle_counter__i4 (.D(n50[4]), .SP(clk_c_enable_175), .CD(n25332), 
            .CK(clk_c), .Q(cycle_counter[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i4.GSR = "DISABLED";
    LUT4 fsm_state_3__bdd_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(fsm_state[0]), .Z(n24202)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B (C (D))))) */ ;
    defparam fsm_state_3__bdd_4_lut.init = 16'h6aa2;
    LUT4 fsm_state_0__bdd_4_lut (.A(fsm_state[0]), .B(fsm_state[2]), .C(fsm_state[1]), 
         .D(fsm_state[3]), .Z(n25462)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;
    defparam fsm_state_0__bdd_4_lut.init = 16'h4555;
    FD1P3IX cycle_counter__i3 (.D(n50[3]), .SP(clk_c_enable_175), .CD(n25332), 
            .CK(clk_c), .Q(cycle_counter[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i3.GSR = "DISABLED";
    FD1P3IX cycle_counter__i2 (.D(n50[2]), .SP(clk_c_enable_175), .CD(n25332), 
            .CK(clk_c), .Q(cycle_counter[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i2.GSR = "DISABLED";
    FD1P3IX cycle_counter__i1 (.D(n50[1]), .SP(clk_c_enable_175), .CD(n25332), 
            .CK(clk_c), .Q(cycle_counter[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(111[8] 119[4])
    defparam cycle_counter__i1.GSR = "DISABLED";
    LUT4 i3490_3_lut_4_lut (.A(cycle_counter[2]), .B(n25391), .C(cycle_counter[3]), 
         .D(cycle_counter[4]), .Z(n50[4])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3490_3_lut_4_lut.init = 16'h7f80;
    LUT4 i21789_3_lut_rep_506_4_lut (.A(fsm_state[0]), .B(n25416), .C(n25276), 
         .D(rst_reg_n), .Z(n25242)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam i21789_3_lut_rep_506_4_lut.init = 16'h01ff;
    LUT4 i4679_2_lut_4_lut_2_lut_3_lut (.A(fsm_state[0]), .B(n25416), .C(rst_reg_n), 
         .Z(n6894)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam i4679_2_lut_4_lut_2_lut_3_lut.init = 16'h1f1f;
    LUT4 i3162_2_lut_rep_581_3_lut_4_lut (.A(fsm_state[0]), .B(n25416), 
         .C(rst_reg_n), .D(next_bit), .Z(clk_c_enable_175)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam i3162_2_lut_rep_581_3_lut_4_lut.init = 16'hffef;
    FD1P3IX data_to_send__i0 (.D(data_to_send_7__N_2305[0]), .SP(clk_c_enable_397), 
            .CD(n17515), .CK(clk_c), .Q(data_to_send[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i0.GSR = "DISABLED";
    LUT4 i11465_4_lut (.A(data_to_send[0]), .B(fsm_state[0]), .C(uart_txd_N_2327), 
         .D(n25416), .Z(uart_txd_N_2325)) /* synthesis lut_function=(A ((D)+!B)+!A !(B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(140[14] 144[8])
    defparam i11465_4_lut.init = 16'haf23;
    LUT4 i21729_4_lut (.A(cycle_counter[0]), .B(cycle_counter[2]), .C(cycle_counter[3]), 
         .D(n22810), .Z(next_bit)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(74[21:71])
    defparam i21729_4_lut.init = 16'h0080;
    FD1P3IX data_to_send__i1 (.D(data_to_send_7__N_2305[1]), .SP(clk_c_enable_397), 
            .CD(n17515), .CK(clk_c), .Q(data_to_send[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i1.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(cycle_counter[1]), .B(cycle_counter[4]), .Z(n22810)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3IX fsm_state__i1 (.D(n122[1]), .SP(next_bit), .CD(n6894), .CK(clk_c), 
            .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam fsm_state__i1.GSR = "DISABLED";
    FD1P3IX fsm_state__i2 (.D(n24203), .SP(next_bit), .CD(n6894), .CK(clk_c), 
            .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1P3IX fsm_state__i3 (.D(n24202), .SP(next_bit), .CD(n6894), .CK(clk_c), 
            .Q(fsm_state[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(124[8] 130[4])
    defparam fsm_state__i3.GSR = "DISABLED";
    FD1P3IX data_to_send__i2 (.D(data_to_send_7__N_2305[2]), .SP(clk_c_enable_397), 
            .CD(n17515), .CK(clk_c), .Q(data_to_send[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i2.GSR = "DISABLED";
    FD1P3IX data_to_send__i3 (.D(data_to_send_7__N_2305[3]), .SP(clk_c_enable_397), 
            .CD(n17515), .CK(clk_c), .Q(data_to_send[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i3.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n25360), .B(n25276), .C(\data_to_write[7] ), 
         .D(rst_reg_n), .Z(n21431)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam i1_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_3_lut_4_lut_adj_463 (.A(n25360), .B(n25276), .C(next_bit), 
         .D(n25242), .Z(clk_c_enable_108)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam i1_3_lut_4_lut_adj_463.init = 16'hfff4;
    LUT4 mux_13_i6_3_lut_4_lut (.A(n25360), .B(n25276), .C(\data_to_write[5] ), 
         .D(data_to_send[6]), .Z(data_to_send_7__N_2305[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i1_3_lut_4_lut (.A(n25360), .B(n25276), .C(\data_to_write[0] ), 
         .D(data_to_send[1]), .Z(data_to_send_7__N_2305[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i7_3_lut_4_lut (.A(n25360), .B(n25276), .C(\data_to_write[6] ), 
         .D(data_to_send[7]), .Z(data_to_send_7__N_2305[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i2_3_lut_4_lut (.A(n25360), .B(n25276), .C(\data_to_write[1] ), 
         .D(data_to_send[2]), .Z(data_to_send_7__N_2305[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i3_3_lut_4_lut (.A(n25360), .B(n25276), .C(\data_to_write[2] ), 
         .D(data_to_send[3]), .Z(data_to_send_7__N_2305[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i4_3_lut_4_lut (.A(n25360), .B(n25276), .C(\data_to_write[3] ), 
         .D(data_to_send[4]), .Z(data_to_send_7__N_2305[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i5_3_lut_4_lut (.A(n25360), .B(n25276), .C(\data_to_write[4] ), 
         .D(data_to_send[5]), .Z(data_to_send_7__N_2305[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(101[17:52])
    defparam mux_13_i5_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX data_to_send__i4 (.D(data_to_send_7__N_2305[4]), .SP(clk_c_enable_397), 
            .CD(n17515), .CK(clk_c), .Q(data_to_send[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=67, LSE_RCOL=6, LSE_LLINE=213, LSE_RLINE=220 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(98[8] 106[4])
    defparam data_to_send__i4.GSR = "DISABLED";
    LUT4 i3471_2_lut_rep_655 (.A(cycle_counter[1]), .B(cycle_counter[0]), 
         .Z(n25391)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3471_2_lut_rep_655.init = 16'h8888;
    LUT4 i3483_2_lut_3_lut_4_lut (.A(cycle_counter[1]), .B(cycle_counter[0]), 
         .C(cycle_counter[3]), .D(cycle_counter[2]), .Z(n50[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3483_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i3476_2_lut_3_lut (.A(cycle_counter[1]), .B(cycle_counter[0]), 
         .C(cycle_counter[2]), .Z(n50[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3476_2_lut_3_lut.init = 16'h7878;
    LUT4 i11532_3_lut_3_lut_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(fsm_state[0]), .Z(n122[1])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(D)))) */ ;
    defparam i11532_3_lut_3_lut_4_lut.init = 16'h33c4;
    LUT4 i1_3_lut_rep_680 (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[3]), 
         .Z(n25416)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(84[17:37])
    defparam i1_3_lut_rep_680.init = 16'hfefe;
    LUT4 uart_txd_I_202_4_lut_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(fsm_state[3]), .Z(uart_txd_N_2327)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(84[17:37])
    defparam uart_txd_I_202_4_lut_3_lut.init = 16'h1e1e;
    LUT4 i1_2_lut_rep_624_4_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[3]), 
         .D(fsm_state[0]), .Z(n25360)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(84[17:37])
    defparam i1_2_lut_rep_624_4_lut.init = 16'hfffe;
    LUT4 i3469_2_lut (.A(cycle_counter[1]), .B(cycle_counter[0]), .Z(n50[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(117[26:46])
    defparam i3469_2_lut.init = 16'h6666;
    LUT4 fsm_state_2__bdd_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(fsm_state[0]), 
         .Z(n24203)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam fsm_state_2__bdd_3_lut.init = 16'h6a6a;
    LUT4 i21791_2_lut_rep_596 (.A(next_bit), .B(rst_reg_n), .Z(n25332)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i21791_2_lut_rep_596.init = 16'hbbbb;
    LUT4 i4294_2_lut_3_lut_4_lut (.A(next_bit), .B(rst_reg_n), .C(cycle_counter[0]), 
         .D(n25360), .Z(n18[0])) /* synthesis lut_function=(!(A (C)+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam i4294_2_lut_3_lut_4_lut.init = 16'h0f4b;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \peripherals_min(CLOCK_MHZ=14) 
//

module \peripherals_min(CLOCK_MHZ=14)  (peri_data_ready, clk_c, n17515, 
            read_en) /* synthesis syn_module_defined=1 */ ;
    output peri_data_ready;
    input clk_c;
    input n17515;
    input read_en;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    FD1S3DX data_ready_51 (.D(read_en), .CK(clk_c), .CD(n17515), .Q(peri_data_ready)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(139[13:35])
    defparam data_ready_51.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module tinyQV
//

module tinyQV (rst_reg_n_adj_10, clk_c, rst_reg_n, peri_data_ready, 
            n25370, n8457, n47, n20728, \addr[2] , \addr[3] , counter_hi, 
            n17512, n20731, n20732, qspi_write_done, data_stall_N_1889, 
            data_stall, n17515, n25321, is_writing_N_2062, n23085, 
            n25151, data_to_write, is_writing, \data_to_write[7] , \data_to_write[6] , 
            \data_to_write[5] , \data_to_write[4] , \data_to_write[3] , 
            \data_to_write[2] , \data_to_write[1] , continue_txn_N_1862, 
            n25320, n25371, n1032, n25154, n23082, n21746, clk_c_enable_354, 
            n6595, next_bit, n25252, uart_txd_N_2327, clk_c_enable_397, 
            n22788, n20638, clk_c_enable_208, n4, clk_c_enable_322, 
            n26, \pc[10] , \pc[11] , \qv_data_read_n[0] , \pc[12] , 
            VCC_net, debug_instr_valid, \pc[13] , \instr_len[2] , \pc[14] , 
            \pc[1] , \addr[0] , \pc[2] , \pc[3] , \pc[4] , \pc[5] , 
            \pc[6] , \pc[7] , \instr_write_offset[3] , n25175, n2015, 
            n2010, \data_from_read[2] , n8229, \gpio_out_sel[7] , n1949, 
            n1969, instr_complete_N_1378, n21541, n8146, n3597, \pc[15] , 
            \qv_data_write_n[0] , \pc[16] , \pc[17] , \next_pc_for_core[3] , 
            \next_pc_for_core[7] , \pc[18] , \imm[19] , \imm[23] , \imm[11] , 
            \imm[15] , \imm[3] , \imm[7] , \imm[18] , \imm[22] , n25363, 
            \imm[10] , \imm[14] , \imm[2] , \imm[6] , \imm[17] , \imm[21] , 
            \imm[9] , \imm[13] , \imm[1] , \imm[5] , mem_op_increment_reg, 
            n23084, \imm[16] , \imm[20] , \imm[8] , \imm[12] , \imm[4] , 
            \next_pc_for_core[4] , \pc[9] , \next_pc_for_core[9] , \next_pc_for_core[13] , 
            \pc[19] , \addr[4] , \addr[5] , \pc[20] , \pc[8] , \instr_avail_len[3] , 
            \next_pc_for_core[8] , \next_pc_for_core[12] , \addr[1] , 
            \addr[6] , \addr[7] , \addr[8] , \addr[9] , \addr[10] , 
            n25194, clk_c_enable_206, \next_pc_for_core[5] , \next_pc_for_core[6] , 
            \next_pc_for_core[10] , \next_pc_for_core[11] , n25417, \next_pc_for_core[14] , 
            \next_pc_for_core[15] , \next_pc_for_core[16] , \next_pc_for_core[17] , 
            \next_pc_for_core[18] , \next_pc_for_core[19] , \next_pc_for_core[20] , 
            \next_pc_for_core[21] , \next_pc_for_core[22] , \pc[21] , 
            \pc[22] , \pc[23] , \next_pc_for_core[23] , n25419, n20582, 
            read_en, \instr_addr_23__N_49[22] , \early_branch_addr[23] , 
            \early_branch_addr[5] , \early_branch_addr[4] , \early_branch_addr[2] , 
            \early_branch_addr[6] , \early_branch_addr[3] , \early_branch_addr[7] , 
            \early_branch_addr[8] , \early_branch_addr[9] , \early_branch_addr[10] , 
            \early_branch_addr[11] , \early_branch_addr[12] , \early_branch_addr[13] , 
            \early_branch_addr[14] , \early_branch_addr[15] , \early_branch_addr[16] , 
            \early_branch_addr[17] , \early_branch_addr[18] , \early_branch_addr[19] , 
            \early_branch_addr[20] , \early_branch_addr[21] , \early_branch_addr[22] , 
            n8527, n22334, \data_from_read[6] , \data_from_read[0] , 
            mem_op_increment_reg_de, n25273, clk_c_enable_27, \next_fsm_state_3__N_2230[3] , 
            \cycle[0] , \ui_in_sync[1] , n1092, debug_rd, accum, d_3__N_1599, 
            \mul_out[1] , \mul_out[3] , n14111, n24186, \mul_out[2] , 
            \next_accum[6] , \next_accum[7] , \next_accum[8] , \next_accum[9] , 
            \next_accum[10] , \next_accum[11] , \next_accum[12] , \next_accum[13] , 
            \next_accum[14] , \next_accum[15] , GND_net, \next_accum[16] , 
            \next_accum[17] , \next_accum[18] , \next_accum[19] , \next_accum[5] , 
            \next_accum[4] ) /* synthesis syn_module_defined=1 */ ;
    output rst_reg_n_adj_10;
    input clk_c;
    input rst_reg_n;
    input peri_data_ready;
    output n25370;
    output n8457;
    input n47;
    output n20728;
    output \addr[2] ;
    output \addr[3] ;
    output [4:2]counter_hi;
    output n17512;
    output n20731;
    input n20732;
    output qspi_write_done;
    output data_stall_N_1889;
    output data_stall;
    output n17515;
    input n25321;
    output is_writing_N_2062;
    input n23085;
    output n25151;
    output [31:0]data_to_write;
    output is_writing;
    output \data_to_write[7] ;
    output \data_to_write[6] ;
    output \data_to_write[5] ;
    output \data_to_write[4] ;
    output \data_to_write[3] ;
    output \data_to_write[2] ;
    output \data_to_write[1] ;
    output continue_txn_N_1862;
    input n25320;
    output n25371;
    output n1032;
    output n25154;
    input n23082;
    output n21746;
    input clk_c_enable_354;
    output n6595;
    input next_bit;
    input n25252;
    input uart_txd_N_2327;
    output clk_c_enable_397;
    input n22788;
    input n20638;
    output clk_c_enable_208;
    input n4;
    output clk_c_enable_322;
    output n26;
    output \pc[10] ;
    output \pc[11] ;
    output \qv_data_read_n[0] ;
    output \pc[12] ;
    input VCC_net;
    output debug_instr_valid;
    output \pc[13] ;
    output \instr_len[2] ;
    output \pc[14] ;
    output \pc[1] ;
    output \addr[0] ;
    output \pc[2] ;
    output \pc[3] ;
    output \pc[4] ;
    output \pc[5] ;
    output \pc[6] ;
    output \pc[7] ;
    output \instr_write_offset[3] ;
    output n25175;
    output n2015;
    output n2010;
    input \data_from_read[2] ;
    input n8229;
    input \gpio_out_sel[7] ;
    input n1949;
    input n1969;
    output instr_complete_N_1378;
    output n21541;
    output n8146;
    output n3597;
    output \pc[15] ;
    output \qv_data_write_n[0] ;
    output \pc[16] ;
    output \pc[17] ;
    input \next_pc_for_core[3] ;
    input \next_pc_for_core[7] ;
    output \pc[18] ;
    output \imm[19] ;
    output \imm[23] ;
    output \imm[11] ;
    output \imm[15] ;
    output \imm[3] ;
    output \imm[7] ;
    output \imm[18] ;
    output \imm[22] ;
    output n25363;
    output \imm[10] ;
    output \imm[14] ;
    output \imm[2] ;
    output \imm[6] ;
    output \imm[17] ;
    output \imm[21] ;
    output \imm[9] ;
    output \imm[13] ;
    output \imm[1] ;
    output \imm[5] ;
    output mem_op_increment_reg;
    input n23084;
    output \imm[16] ;
    output \imm[20] ;
    output \imm[8] ;
    output \imm[12] ;
    output \imm[4] ;
    input \next_pc_for_core[4] ;
    output \pc[9] ;
    input \next_pc_for_core[9] ;
    input \next_pc_for_core[13] ;
    output \pc[19] ;
    output \addr[4] ;
    output \addr[5] ;
    output \pc[20] ;
    output \pc[8] ;
    input \instr_avail_len[3] ;
    input \next_pc_for_core[8] ;
    input \next_pc_for_core[12] ;
    output \addr[1] ;
    output \addr[6] ;
    output \addr[7] ;
    output \addr[8] ;
    output \addr[9] ;
    output \addr[10] ;
    input n25194;
    output clk_c_enable_206;
    input \next_pc_for_core[5] ;
    input \next_pc_for_core[6] ;
    input \next_pc_for_core[10] ;
    input \next_pc_for_core[11] ;
    input n25417;
    input \next_pc_for_core[14] ;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[16] ;
    input \next_pc_for_core[17] ;
    input \next_pc_for_core[18] ;
    input \next_pc_for_core[19] ;
    input \next_pc_for_core[20] ;
    input \next_pc_for_core[21] ;
    input \next_pc_for_core[22] ;
    output \pc[21] ;
    output \pc[22] ;
    output \pc[23] ;
    input \next_pc_for_core[23] ;
    output n25419;
    output n20582;
    output read_en;
    input \instr_addr_23__N_49[22] ;
    input \early_branch_addr[23] ;
    input \early_branch_addr[5] ;
    input \early_branch_addr[4] ;
    input \early_branch_addr[2] ;
    input \early_branch_addr[6] ;
    input \early_branch_addr[3] ;
    input \early_branch_addr[7] ;
    input \early_branch_addr[8] ;
    input \early_branch_addr[9] ;
    input \early_branch_addr[10] ;
    input \early_branch_addr[11] ;
    input \early_branch_addr[12] ;
    input \early_branch_addr[13] ;
    input \early_branch_addr[14] ;
    input \early_branch_addr[15] ;
    input \early_branch_addr[16] ;
    input \early_branch_addr[17] ;
    input \early_branch_addr[18] ;
    input \early_branch_addr[19] ;
    input \early_branch_addr[20] ;
    input \early_branch_addr[21] ;
    input \early_branch_addr[22] ;
    input n8527;
    output n22334;
    input \data_from_read[6] ;
    input \data_from_read[0] ;
    output mem_op_increment_reg_de;
    output n25273;
    input clk_c_enable_27;
    input \next_fsm_state_3__N_2230[3] ;
    output \cycle[0] ;
    input \ui_in_sync[1] ;
    output n1092;
    output [3:0]debug_rd;
    output [15:0]accum;
    output [19:0]d_3__N_1599;
    input \mul_out[1] ;
    input \mul_out[3] ;
    output n14111;
    input n24186;
    input \mul_out[2] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input GND_net;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[5] ;
    input \next_accum[4] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire mem_data_ready, n12, n10, n22566, n22550;
    wire [27:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    
    wire n22552, n25431, n22542, n22538, n22548, n22530, n26612, 
        n25337, n25432, n25334, n25342, n25340, instr_fetch_stopped;
    wire [1:0]data_txn_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(49[15:27])
    
    wire instr_active, start_instr;
    wire [15:0]instr_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(61[15:25])
    wire [31:0]qspi_data_buf;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(58[16:29])
    wire [31:0]mem_data_from_read;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(74[15:33])
    
    wire instr_fetch_running_N_676, n25161, debug_stall_txn, debug_data_continue, 
        qspi_data_ready;
    wire [23:1]instr_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(56[15:25])
    wire [24:0]addr_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(57[17:24])
    
    wire n22873;
    wire [3:1]next_instr_write_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[16:39])
    
    wire n25253, n23038, n23037, n24929, n24935, n24998, instr_fetch_running, 
        n25336, n25324, n21800, n25163, n25403, n25272, n1, n25361;
    wire [31:0]data_to_write_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(56[17:30])
    
    wire n25304;
    wire [1:0]txn_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(56[16:23])
    
    wire spi_ram_b_select_N_2044;
    wire [1:0]qv_data_read_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(65[15:29])
    wire [1:0]qv_data_write_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(64[15:30])
    
    FD1S3AX rst_reg_n_16 (.D(rst_reg_n), .CK(clk_c), .Q(rst_reg_n_adj_10)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=111, LSE_RLINE=150 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(92[10:43])
    defparam rst_reg_n_16.GSR = "DISABLED";
    LUT4 i25_4_lut (.A(mem_data_ready), .B(peri_data_ready), .C(n25370), 
         .D(n12), .Z(n10)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C)+!B !((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(77[26:62])
    defparam i25_4_lut.init = 16'h3505;
    LUT4 i26_4_lut (.A(n22566), .B(n8457), .C(n47), .D(n20728), .Z(n12)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(77[26:62])
    defparam i26_4_lut.init = 16'h3a30;
    LUT4 i1_4_lut (.A(n22550), .B(addr[27]), .C(n22552), .D(n25431), 
         .Z(n8457)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i1_4_lut_adj_457 (.A(addr[18]), .B(n22542), .C(n22538), .D(addr[21]), 
         .Z(n22550)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_4_lut_adj_457.init = 16'hfffe;
    LUT4 i1_4_lut_adj_458 (.A(addr[17]), .B(n22548), .C(n22530), .D(addr[20]), 
         .Z(n22552)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_4_lut_adj_458.init = 16'hfffe;
    LUT4 i1_2_lut (.A(addr[24]), .B(addr[23]), .Z(n22542)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_459 (.A(addr[14]), .B(addr[19]), .Z(n22538)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_adj_459.init = 16'heeee;
    LUT4 i1_4_lut_adj_460 (.A(addr[12]), .B(addr[13]), .C(addr[15]), .D(addr[11]), 
         .Z(n22548)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_4_lut_adj_460.init = 16'hfffe;
    LUT4 i1_2_lut_adj_461 (.A(addr[16]), .B(addr[22]), .Z(n22530)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_adj_461.init = 16'heeee;
    LUT4 i1_2_lut_adj_462 (.A(\addr[2] ), .B(\addr[3] ), .Z(n20728)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(77[26:62])
    defparam i1_2_lut_adj_462.init = 16'h8888;
    FD1S3AX rst_reg_n_16_rep_712 (.D(rst_reg_n), .CK(clk_c), .Q(n26612)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=111, LSE_RLINE=150 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(92[10:43])
    defparam rst_reg_n_16_rep_712.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_695 (.A(addr[26]), .B(addr[25]), .Z(n25431)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_rep_695.init = 16'heeee;
    LUT4 i21934_2_lut_rep_601_3_lut_4_lut (.A(addr[26]), .B(addr[25]), .C(counter_hi[3]), 
         .D(addr[27]), .Z(n25337)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i21934_2_lut_rep_601_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_rep_598_3_lut_4_lut (.A(addr[26]), .B(addr[25]), .C(n25432), 
         .D(addr[27]), .Z(n25334)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_rep_598_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i11755_2_lut_rep_606_3_lut_4_lut (.A(addr[26]), .B(addr[25]), .C(n25432), 
         .D(addr[27]), .Z(n25342)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i11755_2_lut_rep_606_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_604_3_lut_4_lut (.A(addr[26]), .B(addr[25]), .C(n17512), 
         .D(addr[27]), .Z(n25340)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_rep_604_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_634_3_lut (.A(addr[26]), .B(addr[25]), .C(addr[27]), 
         .Z(n25370)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_rep_634_3_lut.init = 16'hfefe;
    tinyqv_mem_ctrl mem (.clk_c(clk_c), .instr_fetch_stopped(instr_fetch_stopped), 
            .data_txn_len({data_txn_len}), .n20731(n20731), .n20732(n20732), 
            .qspi_write_done(qspi_write_done), .instr_active(instr_active), 
            .start_instr(start_instr), .instr_data({instr_data}), .data_stall_N_1889(data_stall_N_1889), 
            .\qspi_data_buf[29] (qspi_data_buf[29]), .\qspi_data_buf[25] (qspi_data_buf[25]), 
            .\mem_data_from_read[23] (mem_data_from_read[23]), .\mem_data_from_read[22] (mem_data_from_read[22]), 
            .\mem_data_from_read[21] (mem_data_from_read[21]), .\mem_data_from_read[20] (mem_data_from_read[20]), 
            .\mem_data_from_read[19] (mem_data_from_read[19]), .\mem_data_from_read[18] (mem_data_from_read[18]), 
            .\mem_data_from_read[17] (mem_data_from_read[17]), .\mem_data_from_read[16] (mem_data_from_read[16]), 
            .\qspi_data_buf[14] (qspi_data_buf[14]), .\qspi_data_buf[12] (qspi_data_buf[12]), 
            .\qspi_data_buf[10] (qspi_data_buf[10]), .\qspi_data_buf[8] (qspi_data_buf[8]), 
            .instr_fetch_running_N_676(instr_fetch_running_N_676), .n25161(n25161), 
            .data_stall(data_stall), .debug_stall_txn(debug_stall_txn), 
            .n17515(n17515), .debug_data_continue(debug_data_continue), 
            .mem_data_ready(mem_data_ready), .\mem_data_from_read[31] (mem_data_from_read[31]), 
            .\mem_data_from_read[27] (mem_data_from_read[27]), .\mem_data_from_read[30] (mem_data_from_read[30]), 
            .\mem_data_from_read[26] (mem_data_from_read[26]), .qspi_data_ready(qspi_data_ready), 
            .\mem_data_from_read[28] (mem_data_from_read[28]), .\mem_data_from_read[24] (mem_data_from_read[24]), 
            .\addr[24] (addr[24]), .\instr_addr[23] (instr_addr[23]), .\addr[23] (addr[23]), 
            .\addr_in[23] (addr_in[23]), .n22873(n22873), .\next_instr_write_offset[3] (next_instr_write_offset[3]), 
            .n25253(n25253), .\mem_data_from_read[13] (mem_data_from_read[13]), 
            .n23038(n23038), .n23037(n23037), .\mem_data_from_read[9] (mem_data_from_read[9]), 
            .n24929(n24929), .n24935(n24935), .n24998(n24998), .\mem_data_from_read[3] (mem_data_from_read[3]), 
            .\mem_data_from_read[4] (mem_data_from_read[4]), .\mem_data_from_read[6] (mem_data_from_read[6]), 
            .\mem_data_from_read[1] (mem_data_from_read[1]), .\mem_data_from_read[5] (mem_data_from_read[5]), 
            .n25321(n25321), .is_writing_N_2062(is_writing_N_2062), .instr_fetch_running(instr_fetch_running), 
            .n25336(n25336), .rst_reg_n(rst_reg_n), .n23085(n23085), .n25432(n25432), 
            .n25370(n25370), .n25324(n25324), .n21800(n21800), .n25163(n25163), 
            .n25151(n25151), .data_to_write({data_to_write_c[31:8], \data_to_write[7] , 
            \data_to_write[6] , \data_to_write[5] , \data_to_write[4] , 
            \data_to_write[3] , \data_to_write[2] , \data_to_write[1] , 
            data_to_write[0]}), .n25403(n25403), .is_writing(is_writing), 
            .n25272(n25272), .n1(n1), .n25361(n25361), .continue_txn_N_1862(continue_txn_N_1862), 
            .n25342(n25342), .n25340(n25340), .n25320(n25320), .n17512(n17512), 
            .n25304(n25304), .n25371(n25371), .\txn_len[1] (txn_len[1]), 
            .n1032(n1032), .n25154(n25154), .spi_ram_b_select_N_2044(spi_ram_b_select_N_2044), 
            .n23082(n23082), .n21746(n21746), .clk_c_enable_354(clk_c_enable_354), 
            .n6595(n6595), .next_bit(next_bit), .n25252(n25252), .uart_txd_N_2327(uart_txd_N_2327), 
            .clk_c_enable_397(clk_c_enable_397), .n22788(n22788), .n20638(n20638), 
            .n25334(n25334), .clk_c_enable_208(clk_c_enable_208), .n4(n4), 
            .clk_c_enable_322(clk_c_enable_322), .\qv_data_read_n[1] (qv_data_read_n[1]), 
            .\qv_data_write_n[1] (qv_data_write_n[1]), .n26(n26)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(132[19] 164[6])
    tinyqv_cpu cpu (.clk_c(clk_c), .instr_data({instr_data}), .\pc[10] (\pc[10] ), 
            .\pc[11] (\pc[11] ), .qv_data_read_n({qv_data_read_n[1], \qv_data_read_n[0] }), 
            .\pc[12] (\pc[12] ), .VCC_net(VCC_net), .debug_instr_valid(debug_instr_valid), 
            .n25370(n25370), .n24935(n24935), .\mem_data_from_read[4] (mem_data_from_read[4]), 
            .counter_hi({counter_hi}), .\pc[13] (\pc[13] ), .n24929(n24929), 
            .\mem_data_from_read[6] (mem_data_from_read[6]), .\instr_len[2] (\instr_len[2] ), 
            .instr_fetch_running(instr_fetch_running), .\pc[14] (\pc[14] ), 
            .\pc[1] (\pc[1] ), .addr({addr[27:11], \addr[10] , \addr[9] , 
            \addr[8] , \addr[7] , \addr[6] , \addr[5] , \addr[4] , 
            \addr[3] , \addr[2] , \addr[1] , \addr[0] }), .\pc[2] (\pc[2] ), 
            .\pc[3] (\pc[3] ), .\pc[4] (\pc[4] ), .\pc[5] (\pc[5] ), .\pc[6] (\pc[6] ), 
            .\pc[7] (\pc[7] ), .\instr_write_offset[3] (\instr_write_offset[3] ), 
            .\next_instr_write_offset[3] (next_instr_write_offset[3]), .rst_reg_n(rst_reg_n_adj_10), 
            .n25175(n25175), .n2015(n2015), .n2010(n2010), .\data_from_read[2] (\data_from_read[2] ), 
            .n8229(n8229), .\gpio_out_sel[7] (\gpio_out_sel[7] ), .n1949(n1949), 
            .n1969(n1969), .n26612(n26612), .instr_complete_N_1378(instr_complete_N_1378), 
            .n21541(n21541), .n8146(n8146), .\qspi_data_buf[25] (qspi_data_buf[25]), 
            .\qspi_data_buf[29] (qspi_data_buf[29]), .qspi_data_ready(qspi_data_ready), 
            .n25361(n25361), .\mem_data_from_read[17] (mem_data_from_read[17]), 
            .\mem_data_from_read[21] (mem_data_from_read[21]), .debug_data_continue(debug_data_continue), 
            .n3597(n3597), .data_to_write({data_to_write_c[31:8], \data_to_write[7] , 
            \data_to_write[6] , \data_to_write[5] , \data_to_write[4] , 
            \data_to_write[3] , \data_to_write[2] , \data_to_write[1] , 
            data_to_write[0]}), .\pc[15] (\pc[15] ), .qv_data_write_n({qv_data_write_n[1], 
            \qv_data_write_n[0] }), .\pc[16] (\pc[16] ), .\mem_data_from_read[27] (mem_data_from_read[27]), 
            .\mem_data_from_read[31] (mem_data_from_read[31]), .\pc[17] (\pc[17] ), 
            .instr_fetch_running_N_676(instr_fetch_running_N_676), .debug_stall_txn(debug_stall_txn), 
            .n21800(n21800), .\next_pc_for_core[3] (\next_pc_for_core[3] ), 
            .\next_pc_for_core[7] (\next_pc_for_core[7] ), .\pc[18] (\pc[18] ), 
            .\imm[19] (\imm[19] ), .\imm[23] (\imm[23] ), .n17512(n17512), 
            .\imm[11] (\imm[11] ), .\imm[15] (\imm[15] ), .\imm[3] (\imm[3] ), 
            .\imm[7] (\imm[7] ), .\imm[18] (\imm[18] ), .\imm[22] (\imm[22] ), 
            .n25363(n25363), .\imm[10] (\imm[10] ), .\imm[14] (\imm[14] ), 
            .\imm[2] (\imm[2] ), .\imm[6] (\imm[6] ), .\imm[17] (\imm[17] ), 
            .\imm[21] (\imm[21] ), .\imm[9] (\imm[9] ), .\imm[13] (\imm[13] ), 
            .\imm[1] (\imm[1] ), .\imm[5] (\imm[5] ), .mem_op_increment_reg(mem_op_increment_reg), 
            .n23084(n23084), .\imm[16] (\imm[16] ), .\imm[20] (\imm[20] ), 
            .\imm[8] (\imm[8] ), .\imm[12] (\imm[12] ), .\imm[4] (\imm[4] ), 
            .\next_pc_for_core[4] (\next_pc_for_core[4] ), .\pc[9] (\pc[9] ), 
            .\next_pc_for_core[9] (\next_pc_for_core[9] ), .\next_pc_for_core[13] (\next_pc_for_core[13] ), 
            .\pc[19] (\pc[19] ), .n10(n10), .n22566(n22566), .\pc[20] (\pc[20] ), 
            .\pc[8] (\pc[8] ), .n25163(n25163), .n25161(n25161), .\instr_avail_len[3] (\instr_avail_len[3] ), 
            .\next_pc_for_core[8] (\next_pc_for_core[8] ), .\next_pc_for_core[12] (\next_pc_for_core[12] ), 
            .n25194(n25194), .n25336(n25336), .clk_c_enable_206(clk_c_enable_206), 
            .\next_pc_for_core[5] (\next_pc_for_core[5] ), .\next_pc_for_core[6] (\next_pc_for_core[6] ), 
            .\next_pc_for_core[10] (\next_pc_for_core[10] ), .\next_pc_for_core[11] (\next_pc_for_core[11] ), 
            .n25417(n25417), .\next_pc_for_core[14] (\next_pc_for_core[14] ), 
            .\next_pc_for_core[15] (\next_pc_for_core[15] ), .\next_pc_for_core[16] (\next_pc_for_core[16] ), 
            .\next_pc_for_core[17] (\next_pc_for_core[17] ), .\next_pc_for_core[18] (\next_pc_for_core[18] ), 
            .\next_pc_for_core[19] (\next_pc_for_core[19] ), .\next_pc_for_core[20] (\next_pc_for_core[20] ), 
            .\next_pc_for_core[21] (\next_pc_for_core[21] ), .\next_pc_for_core[22] (\next_pc_for_core[22] ), 
            .data_txn_len({data_txn_len}), .\qspi_data_buf[14] (qspi_data_buf[14]), 
            .n25253(n25253), .\pc[21] (\pc[21] ), .\pc[22] (\pc[22] ), 
            .\pc[23] (\pc[23] ), .\next_pc_for_core[23] (\next_pc_for_core[23] ), 
            .\qspi_data_buf[10] (qspi_data_buf[10]), .n25419(n25419), .\mem_data_from_read[19] (mem_data_from_read[19]), 
            .\mem_data_from_read[23] (mem_data_from_read[23]), .n25431(n25431), 
            .n25432(n25432), .n25324(n25324), .n20582(n20582), .\mem_data_from_read[16] (mem_data_from_read[16]), 
            .\mem_data_from_read[20] (mem_data_from_read[20]), .\mem_data_from_read[18] (mem_data_from_read[18]), 
            .\mem_data_from_read[22] (mem_data_from_read[22]), .\mem_data_from_read[3] (mem_data_from_read[3]), 
            .read_en(read_en), .\qspi_data_buf[12] (qspi_data_buf[12]), 
            .\instr_addr_23__N_49[22] (\instr_addr_23__N_49[22] ), .\early_branch_addr[23] (\early_branch_addr[23] ), 
            .\instr_addr[23] (instr_addr[23]), .instr_fetch_stopped(instr_fetch_stopped), 
            .\early_branch_addr[5] (\early_branch_addr[5] ), .\early_branch_addr[4] (\early_branch_addr[4] ), 
            .\early_branch_addr[2] (\early_branch_addr[2] ), .\early_branch_addr[6] (\early_branch_addr[6] ), 
            .\early_branch_addr[3] (\early_branch_addr[3] ), .\early_branch_addr[7] (\early_branch_addr[7] ), 
            .\early_branch_addr[8] (\early_branch_addr[8] ), .\early_branch_addr[9] (\early_branch_addr[9] ), 
            .\early_branch_addr[10] (\early_branch_addr[10] ), .\early_branch_addr[11] (\early_branch_addr[11] ), 
            .\early_branch_addr[12] (\early_branch_addr[12] ), .\early_branch_addr[13] (\early_branch_addr[13] ), 
            .\early_branch_addr[14] (\early_branch_addr[14] ), .\early_branch_addr[15] (\early_branch_addr[15] ), 
            .\early_branch_addr[16] (\early_branch_addr[16] ), .\early_branch_addr[17] (\early_branch_addr[17] ), 
            .\early_branch_addr[18] (\early_branch_addr[18] ), .\early_branch_addr[19] (\early_branch_addr[19] ), 
            .\early_branch_addr[20] (\early_branch_addr[20] ), .\early_branch_addr[21] (\early_branch_addr[21] ), 
            .\early_branch_addr[22] (\early_branch_addr[22] ), .\qspi_data_buf[8] (qspi_data_buf[8]), 
            .n25304(n25304), .instr_active(instr_active), .\txn_len[1] (txn_len[1]), 
            .n8527(n8527), .n25403(n25403), .\addr_in[23] (addr_in[23]), 
            .spi_ram_b_select_N_2044(spi_ram_b_select_N_2044), .n23037(n23037), 
            .n23038(n23038), .n1(n1), .n22873(n22873), .\mem_data_from_read[1] (mem_data_from_read[1]), 
            .\mem_data_from_read[5] (mem_data_from_read[5]), .\mem_data_from_read[9] (mem_data_from_read[9]), 
            .\mem_data_from_read[13] (mem_data_from_read[13]), .n25272(n25272), 
            .n22334(n22334), .n25337(n25337), .\mem_data_from_read[24] (mem_data_from_read[24]), 
            .\mem_data_from_read[28] (mem_data_from_read[28]), .\mem_data_from_read[26] (mem_data_from_read[26]), 
            .\mem_data_from_read[30] (mem_data_from_read[30]), .mem_data_ready(mem_data_ready), 
            .\data_from_read[6] (\data_from_read[6] ), .\data_from_read[0] (\data_from_read[0] ), 
            .start_instr(start_instr), .n24998(n24998), .mem_op_increment_reg_de(mem_op_increment_reg_de), 
            .n25273(n25273), .clk_c_enable_27(clk_c_enable_27), .\next_fsm_state_3__N_2230[3] (\next_fsm_state_3__N_2230[3] ), 
            .\cycle[0] (\cycle[0] ), .\ui_in_sync[1] (\ui_in_sync[1] ), 
            .n1092(n1092), .debug_rd({debug_rd}), .accum({accum}), .d_3__N_1599({d_3__N_1599}), 
            .\mul_out[1] (\mul_out[1] ), .\mul_out[3] (\mul_out[3] ), .n14111(n14111), 
            .n24186(n24186), .\mul_out[2] (\mul_out[2] ), .\next_accum[6] (\next_accum[6] ), 
            .\next_accum[7] (\next_accum[7] ), .\next_accum[8] (\next_accum[8] ), 
            .\next_accum[9] (\next_accum[9] ), .\next_accum[10] (\next_accum[10] ), 
            .\next_accum[11] (\next_accum[11] ), .\next_accum[12] (\next_accum[12] ), 
            .\next_accum[13] (\next_accum[13] ), .\next_accum[14] (\next_accum[14] ), 
            .\next_accum[15] (\next_accum[15] ), .GND_net(GND_net), .\next_accum[16] (\next_accum[16] ), 
            .\next_accum[17] (\next_accum[17] ), .\next_accum[18] (\next_accum[18] ), 
            .\next_accum[19] (\next_accum[19] ), .\next_accum[5] (\next_accum[5] ), 
            .\next_accum[4] (\next_accum[4] )) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(94[14] 130[6])
    
endmodule
//
// Verilog Description of module tinyqv_mem_ctrl
//

module tinyqv_mem_ctrl (clk_c, instr_fetch_stopped, data_txn_len, n20731, 
            n20732, qspi_write_done, instr_active, start_instr, instr_data, 
            data_stall_N_1889, \qspi_data_buf[29] , \qspi_data_buf[25] , 
            \mem_data_from_read[23] , \mem_data_from_read[22] , \mem_data_from_read[21] , 
            \mem_data_from_read[20] , \mem_data_from_read[19] , \mem_data_from_read[18] , 
            \mem_data_from_read[17] , \mem_data_from_read[16] , \qspi_data_buf[14] , 
            \qspi_data_buf[12] , \qspi_data_buf[10] , \qspi_data_buf[8] , 
            instr_fetch_running_N_676, n25161, data_stall, debug_stall_txn, 
            n17515, debug_data_continue, mem_data_ready, \mem_data_from_read[31] , 
            \mem_data_from_read[27] , \mem_data_from_read[30] , \mem_data_from_read[26] , 
            qspi_data_ready, \mem_data_from_read[28] , \mem_data_from_read[24] , 
            \addr[24] , \instr_addr[23] , \addr[23] , \addr_in[23] , 
            n22873, \next_instr_write_offset[3] , n25253, \mem_data_from_read[13] , 
            n23038, n23037, \mem_data_from_read[9] , n24929, n24935, 
            n24998, \mem_data_from_read[3] , \mem_data_from_read[4] , 
            \mem_data_from_read[6] , \mem_data_from_read[1] , \mem_data_from_read[5] , 
            n25321, is_writing_N_2062, instr_fetch_running, n25336, 
            rst_reg_n, n23085, n25432, n25370, n25324, n21800, n25163, 
            n25151, data_to_write, n25403, is_writing, n25272, n1, 
            n25361, continue_txn_N_1862, n25342, n25340, n25320, n17512, 
            n25304, n25371, \txn_len[1] , n1032, n25154, spi_ram_b_select_N_2044, 
            n23082, n21746, clk_c_enable_354, n6595, next_bit, n25252, 
            uart_txd_N_2327, clk_c_enable_397, n22788, n20638, n25334, 
            clk_c_enable_208, n4, clk_c_enable_322, \qv_data_read_n[1] , 
            \qv_data_write_n[1] , n26) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output instr_fetch_stopped;
    output [1:0]data_txn_len;
    output n20731;
    input n20732;
    output qspi_write_done;
    output instr_active;
    input start_instr;
    output [15:0]instr_data;
    output data_stall_N_1889;
    output \qspi_data_buf[29] ;
    output \qspi_data_buf[25] ;
    output \mem_data_from_read[23] ;
    output \mem_data_from_read[22] ;
    output \mem_data_from_read[21] ;
    output \mem_data_from_read[20] ;
    output \mem_data_from_read[19] ;
    output \mem_data_from_read[18] ;
    output \mem_data_from_read[17] ;
    output \mem_data_from_read[16] ;
    output \qspi_data_buf[14] ;
    output \qspi_data_buf[12] ;
    output \qspi_data_buf[10] ;
    output \qspi_data_buf[8] ;
    output instr_fetch_running_N_676;
    input n25161;
    output data_stall;
    output debug_stall_txn;
    output n17515;
    input debug_data_continue;
    output mem_data_ready;
    output \mem_data_from_read[31] ;
    output \mem_data_from_read[27] ;
    output \mem_data_from_read[30] ;
    output \mem_data_from_read[26] ;
    output qspi_data_ready;
    output \mem_data_from_read[28] ;
    output \mem_data_from_read[24] ;
    input \addr[24] ;
    input \instr_addr[23] ;
    input \addr[23] ;
    output \addr_in[23] ;
    input n22873;
    input \next_instr_write_offset[3] ;
    output n25253;
    output \mem_data_from_read[13] ;
    output n23038;
    output n23037;
    output \mem_data_from_read[9] ;
    output n24929;
    output n24935;
    output n24998;
    output \mem_data_from_read[3] ;
    output \mem_data_from_read[4] ;
    output \mem_data_from_read[6] ;
    output \mem_data_from_read[1] ;
    output \mem_data_from_read[5] ;
    input n25321;
    output is_writing_N_2062;
    input instr_fetch_running;
    output n25336;
    input rst_reg_n;
    input n23085;
    input n25432;
    input n25370;
    input n25324;
    input n21800;
    input n25163;
    output n25151;
    input [31:0]data_to_write;
    output n25403;
    output is_writing;
    input n25272;
    input n1;
    output n25361;
    output continue_txn_N_1862;
    input n25342;
    input n25340;
    input n25320;
    input n17512;
    output n25304;
    output n25371;
    input \txn_len[1] ;
    output n1032;
    output n25154;
    input spi_ram_b_select_N_2044;
    input n23082;
    output n21746;
    input clk_c_enable_354;
    output n6595;
    input next_bit;
    input n25252;
    input uart_txd_N_2327;
    output clk_c_enable_397;
    input n22788;
    input n20638;
    input n25334;
    output clk_c_enable_208;
    input n4;
    output clk_c_enable_322;
    input \qv_data_read_n[1] ;
    input \qv_data_write_n[1] ;
    output n26;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [1:0]qspi_data_byte_idx;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(59[15:33])
    
    wire clk_c_enable_26, qspi_data_byte_idx_1__N_1756;
    wire [1:0]n174;
    
    wire n9, n6611, debug_stop_txn_N_1850, clk_c_enable_43, n9278, 
        data_ready_N_1840, clk_c_enable_52, instr_active_N_1837, clk_c_enable_157;
    wire [31:0]instr_data_7__N_1700;
    
    wire n8138, data_ready_N_1839, n2;
    wire [1:0]write_qspi_data_byte_idx_1__N_1752;
    wire [31:0]qspi_data_buf;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(58[16:29])
    
    wire clk_c_enable_134, clk_c_enable_142, clk_c_enable_150, n8460;
    wire [2:0]fsm_state;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(82[15:24])
    
    wire n25471, n25174, n25384, n1002, n25172, n25355, n25353, 
        n19413;
    wire [1:0]read_cycles_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(105[15:32])
    
    wire n25170, n5, n57;
    wire [1:0]n333;
    
    wire continue_txn, clk_c_enable_193, debug_stop_txn_N_1851, n24335, 
        n25275, clk_c_enable_103, n18783, n25150, n25414, n36, n21878, 
        n20682, n25302, n5278, n25423, debug_stop_txn_N_1873, n21854, 
        n25392, n8888, n25393, spi_ram_a_select_N_2040, n25325, spi_clk_pos, 
        stop_txn_now_N_2094, n4_c, n25364, n25286, n23026, n23016, 
        n23013, n23014, n23019, n23020, n23022, n23031, n23029, 
        n23032, n23035, n24195, n23023, n23034, n23025, n23028;
    wire [1:0]write_qspi_data_byte_idx;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[16:40])
    
    wire n25159;
    wire [24:0]addr_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(57[17:24])
    wire [1:0]txn_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(56[16:23])
    
    wire n25470, n25472;
    
    FD1P3IX qspi_data_byte_idx__i1 (.D(n174[1]), .SP(clk_c_enable_26), .CD(qspi_data_byte_idx_1__N_1756), 
            .CK(clk_c), .Q(qspi_data_byte_idx[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam qspi_data_byte_idx__i1.GSR = "DISABLED";
    FD1P3IX qspi_data_byte_idx__i0 (.D(n9), .SP(clk_c_enable_26), .CD(qspi_data_byte_idx_1__N_1756), 
            .CK(clk_c), .Q(qspi_data_byte_idx[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam qspi_data_byte_idx__i0.GSR = "DISABLED";
    FD1S3IX instr_fetch_stopped_182 (.D(debug_stop_txn_N_1850), .CK(clk_c), 
            .CD(n6611), .Q(instr_fetch_stopped)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam instr_fetch_stopped_182.GSR = "DISABLED";
    FD1P3AX data_txn_len_i0_i1 (.D(n20731), .SP(clk_c_enable_43), .CK(clk_c), 
            .Q(data_txn_len[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(177[12] 183[8])
    defparam data_txn_len_i0_i1.GSR = "DISABLED";
    FD1P3AX data_txn_len_i0_i0 (.D(n20732), .SP(clk_c_enable_43), .CK(clk_c), 
            .Q(data_txn_len[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(177[12] 183[8])
    defparam data_txn_len_i0_i0.GSR = "DISABLED";
    FD1S3IX qspi_write_done_185 (.D(data_ready_N_1840), .CK(clk_c), .CD(n9278), 
            .Q(qspi_write_done)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(173[12] 175[8])
    defparam qspi_write_done_185.GSR = "DISABLED";
    FD1P3IX instr_active_180 (.D(start_instr), .SP(clk_c_enable_52), .CD(instr_active_N_1837), 
            .CK(clk_c), .Q(instr_active)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(103[12] 109[8])
    defparam instr_active_180.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i1 (.D(instr_data_7__N_1700[0]), .SP(clk_c_enable_157), 
            .CK(clk_c), .Q(instr_data[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i1.GSR = "DISABLED";
    LUT4 continue_txn_I_164_4_lut (.A(n8138), .B(data_ready_N_1839), .C(n2), 
         .D(write_qspi_data_byte_idx_1__N_1752[0]), .Z(data_stall_N_1889)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(190[21] 191[76])
    defparam continue_txn_I_164_4_lut.init = 16'hcecc;
    FD1P3AX qspi_data_buf_i32 (.D(instr_data_7__N_1700[31]), .SP(clk_c_enable_134), 
            .CK(clk_c), .Q(qspi_data_buf[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i32.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i31 (.D(instr_data_7__N_1700[30]), .SP(clk_c_enable_134), 
            .CK(clk_c), .Q(qspi_data_buf[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i31.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i30 (.D(instr_data_7__N_1700[29]), .SP(clk_c_enable_134), 
            .CK(clk_c), .Q(\qspi_data_buf[29] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i30.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i29 (.D(instr_data_7__N_1700[28]), .SP(clk_c_enable_134), 
            .CK(clk_c), .Q(qspi_data_buf[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i29.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i28 (.D(instr_data_7__N_1700[27]), .SP(clk_c_enable_134), 
            .CK(clk_c), .Q(qspi_data_buf[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i28.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i27 (.D(instr_data_7__N_1700[26]), .SP(clk_c_enable_134), 
            .CK(clk_c), .Q(qspi_data_buf[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i27.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i26 (.D(instr_data_7__N_1700[25]), .SP(clk_c_enable_134), 
            .CK(clk_c), .Q(\qspi_data_buf[25] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i26.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i25 (.D(instr_data_7__N_1700[24]), .SP(clk_c_enable_134), 
            .CK(clk_c), .Q(qspi_data_buf[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i25.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i24 (.D(instr_data_7__N_1700[23]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(\mem_data_from_read[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i24.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i23 (.D(instr_data_7__N_1700[22]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(\mem_data_from_read[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i23.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i22 (.D(instr_data_7__N_1700[21]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(\mem_data_from_read[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i22.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i21 (.D(instr_data_7__N_1700[20]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(\mem_data_from_read[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i21.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i20 (.D(instr_data_7__N_1700[19]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(\mem_data_from_read[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i20.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i19 (.D(instr_data_7__N_1700[18]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(\mem_data_from_read[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i19.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i18 (.D(instr_data_7__N_1700[17]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(\mem_data_from_read[17] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i18.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i17 (.D(instr_data_7__N_1700[16]), .SP(clk_c_enable_142), 
            .CK(clk_c), .Q(\mem_data_from_read[16] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i17.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i16 (.D(instr_data_7__N_1700[15]), .SP(clk_c_enable_150), 
            .CK(clk_c), .Q(qspi_data_buf[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i16.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i15 (.D(instr_data_7__N_1700[14]), .SP(clk_c_enable_150), 
            .CK(clk_c), .Q(\qspi_data_buf[14] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i15.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i14 (.D(instr_data_7__N_1700[13]), .SP(clk_c_enable_150), 
            .CK(clk_c), .Q(qspi_data_buf[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i14.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i13 (.D(instr_data_7__N_1700[12]), .SP(clk_c_enable_150), 
            .CK(clk_c), .Q(\qspi_data_buf[12] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i13.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i12 (.D(instr_data_7__N_1700[11]), .SP(clk_c_enable_150), 
            .CK(clk_c), .Q(qspi_data_buf[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i12.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i11 (.D(instr_data_7__N_1700[10]), .SP(clk_c_enable_150), 
            .CK(clk_c), .Q(\qspi_data_buf[10] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i11.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i10 (.D(instr_data_7__N_1700[9]), .SP(clk_c_enable_150), 
            .CK(clk_c), .Q(qspi_data_buf[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i10.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i9 (.D(instr_data_7__N_1700[8]), .SP(clk_c_enable_150), 
            .CK(clk_c), .Q(\qspi_data_buf[8] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i9.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i8 (.D(instr_data_7__N_1700[7]), .SP(clk_c_enable_157), 
            .CK(clk_c), .Q(instr_data[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i8.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i7 (.D(instr_data_7__N_1700[6]), .SP(clk_c_enable_157), 
            .CK(clk_c), .Q(instr_data[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i7.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i6 (.D(instr_data_7__N_1700[5]), .SP(clk_c_enable_157), 
            .CK(clk_c), .Q(instr_data[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i6.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i5 (.D(instr_data_7__N_1700[4]), .SP(clk_c_enable_157), 
            .CK(clk_c), .Q(instr_data[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i5.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i4 (.D(instr_data_7__N_1700[3]), .SP(clk_c_enable_157), 
            .CK(clk_c), .Q(instr_data[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i4.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i3 (.D(instr_data_7__N_1700[2]), .SP(clk_c_enable_157), 
            .CK(clk_c), .Q(instr_data[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i3.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i2 (.D(instr_data_7__N_1700[1]), .SP(clk_c_enable_157), 
            .CK(clk_c), .Q(instr_data[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i2.GSR = "DISABLED";
    FD1S3IX instr_fetch_started_181 (.D(n25161), .CK(clk_c), .CD(n8460), 
            .Q(instr_fetch_running_N_676)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam instr_fetch_started_181.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(qspi_data_byte_idx[0]), .B(data_txn_len[0]), .Z(n8138)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i1_2_lut.init = 16'h6666;
    LUT4 continue_txn_I_165_i2_3_lut (.A(qspi_data_byte_idx[1]), .B(data_txn_len[1]), 
         .C(qspi_data_byte_idx[0]), .Z(n2)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(190[39:81])
    defparam continue_txn_I_165_i2_3_lut.init = 16'h9696;
    LUT4 n24336_bdd_3_lut_rep_432_4_lut_then_4_lut (.A(data_stall), .B(debug_stall_txn), 
         .C(fsm_state[2]), .D(fsm_state[1]), .Z(n25471)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam n24336_bdd_3_lut_rep_432_4_lut_then_4_lut.init = 16'he0ef;
    LUT4 i1_2_lut_rep_438 (.A(data_stall), .B(debug_stall_txn), .Z(n25174)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_438.init = 16'heeee;
    LUT4 i6899_3_lut_rep_436_4_lut (.A(data_stall), .B(debug_stall_txn), 
         .C(n25384), .D(n1002), .Z(n25172)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i6899_3_lut_rep_436_4_lut.init = 16'hefe0;
    LUT4 i22_3_lut_4_lut (.A(data_stall), .B(debug_stall_txn), .C(n25355), 
         .D(n25353), .Z(n19413)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam i22_3_lut_4_lut.init = 16'hf101;
    LUT4 i1_2_lut_rep_434_3_lut (.A(data_stall), .B(debug_stall_txn), .C(read_cycles_count[1]), 
         .Z(n25170)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_434_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(data_stall), .B(debug_stall_txn), .C(n5), 
         .D(read_cycles_count[1]), .Z(n57)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_106_i2_3_lut_4_lut (.A(data_stall), .B(debug_stall_txn), .C(n25384), 
         .D(n1002), .Z(n333[1])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_106_i2_3_lut_4_lut.init = 16'hefe0;
    FD1P3IX continue_txn_187 (.D(debug_data_continue), .SP(clk_c_enable_193), 
            .CD(n17515), .CK(clk_c), .Q(continue_txn)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam continue_txn_187.GSR = "DISABLED";
    LUT4 qspi_data_buf_31__I_0_189_3_lut (.A(qspi_data_buf[31]), .B(instr_data[15]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[31] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_31__I_0_189_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_27__I_0_3_lut (.A(qspi_data_buf[27]), .B(instr_data[11]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[27] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_27__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_30__I_0_3_lut (.A(qspi_data_buf[30]), .B(instr_data[14]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[30] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_30__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_26__I_0_3_lut (.A(qspi_data_buf[26]), .B(instr_data[10]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[26] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_26__I_0_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_4_lut (.A(continue_txn), .B(data_ready_N_1840), 
         .C(write_qspi_data_byte_idx_1__N_1752[0]), .D(qspi_data_ready), 
         .Z(debug_stop_txn_N_1851)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[102:115])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 qspi_data_buf_28__I_0_3_lut (.A(qspi_data_buf[28]), .B(instr_data[12]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[28] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_28__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_24__I_0_3_lut (.A(qspi_data_buf[24]), .B(instr_data[8]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_24__I_0_3_lut.init = 16'hcaca;
    LUT4 n57_bdd_2_lut_3_lut (.A(instr_active), .B(start_instr), .C(\addr[24] ), 
         .Z(n24335)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam n57_bdd_2_lut_3_lut.init = 16'hefef;
    LUT4 mux_2710_i1_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr[23] ), 
         .D(\addr[23] ), .Z(\addr_in[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam mux_2710_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_414_3_lut_4_lut (.A(n25275), .B(start_instr), .C(clk_c_enable_103), 
         .D(n18783), .Z(n25150)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i1_2_lut_rep_414_3_lut_4_lut.init = 16'hd000;
    LUT4 i1_4_lut (.A(qspi_data_ready), .B(n22873), .C(n25414), .D(\next_instr_write_offset[3] ), 
         .Z(n36)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(39[23:37])
    defparam i1_4_lut.init = 16'h3b0a;
    LUT4 qspi_data_buf_15__I_0_i6_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), 
         .C(instr_data[13]), .D(qspi_data_buf[13]), .Z(\mem_data_from_read[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam qspi_data_buf_15__I_0_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 i20763_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), .C(instr_data[15]), 
         .D(qspi_data_buf[15]), .Z(n23038)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i20763_3_lut_4_lut.init = 16'hf780;
    LUT4 i20762_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), .C(instr_data[11]), 
         .D(qspi_data_buf[11]), .Z(n23037)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i20762_3_lut_4_lut.init = 16'hf780;
    LUT4 qspi_data_buf_15__I_0_i2_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), 
         .C(instr_data[9]), .D(qspi_data_buf[9]), .Z(\mem_data_from_read[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam qspi_data_buf_15__I_0_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mem_data_from_read_6__bdd_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), 
         .C(instr_data[10]), .D(instr_data[2]), .Z(n24929)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mem_data_from_read_6__bdd_3_lut_4_lut.init = 16'hfb40;
    LUT4 mem_data_from_read_4__bdd_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), 
         .C(instr_data[8]), .D(instr_data[0]), .Z(n24935)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mem_data_from_read_4__bdd_3_lut_4_lut.init = 16'hfb40;
    LUT4 n4956_bdd_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), .C(instr_data[15]), 
         .D(instr_data[7]), .Z(n24998)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam n4956_bdd_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i4_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), 
         .C(instr_data[11]), .D(instr_data[3]), .Z(\mem_data_from_read[3] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i5_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), 
         .C(instr_data[12]), .D(instr_data[4]), .Z(\mem_data_from_read[4] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i7_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), 
         .C(instr_data[14]), .D(instr_data[6]), .Z(\mem_data_from_read[6] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i2_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), 
         .C(instr_data[9]), .D(instr_data[1]), .Z(\mem_data_from_read[1] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i6_3_lut_4_lut (.A(data_txn_len[0]), .B(n25253), 
         .C(instr_data[13]), .D(instr_data[5]), .Z(\mem_data_from_read[5] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_3_lut (.A(start_instr), .B(n25321), .C(n21878), .Z(is_writing_N_2062)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_4_lut_3_lut.init = 16'h4040;
    LUT4 data_ready_I_0_206_4_lut (.A(instr_active), .B(n20682), .C(n25302), 
         .D(data_ready_N_1839), .Z(mem_data_ready)) /* synthesis lut_function=(!(A+!(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[25:190])
    defparam data_ready_I_0_206_4_lut.init = 16'h5545;
    LUT4 qspi_data_ready_I_0_202_2_lut (.A(qspi_data_ready), .B(data_ready_N_1840), 
         .Z(data_ready_N_1839)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[43:98])
    defparam qspi_data_ready_I_0_202_2_lut.init = 16'h8888;
    LUT4 i21709_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(data_txn_len[0]), .D(data_txn_len[1]), .Z(data_ready_N_1840)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[64:98])
    defparam i21709_4_lut.init = 16'h8421;
    LUT4 i1_3_lut_rep_600_4_lut (.A(instr_active), .B(n25414), .C(instr_fetch_running), 
         .D(qspi_data_ready), .Z(n25336)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(103[12] 109[8])
    defparam i1_3_lut_rep_600_4_lut.init = 16'h2000;
    FD1P3IX data_stall_188 (.D(n23085), .SP(rst_reg_n), .CD(n5278), .CK(clk_c), 
            .Q(data_stall)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam data_stall_188.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_445 (.A(n25423), .B(data_stall), .C(n25432), 
         .D(n25370), .Z(n20682)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i1_2_lut_3_lut_4_lut_adj_445.init = 16'h0004;
    LUT4 i11496_4_lut (.A(n25324), .B(n21800), .C(n36), .D(n25163), 
         .Z(debug_stop_txn_N_1873)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[26] 86[20])
    defparam i11496_4_lut.init = 16'heca0;
    LUT4 i1_2_lut_rep_415_3_lut_4_lut (.A(n25321), .B(n25302), .C(n18783), 
         .D(start_instr), .Z(n25151)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_rep_415_3_lut_4_lut.init = 16'hf070;
    LUT4 i21898_4_lut (.A(qspi_data_byte_idx[0]), .B(n21854), .C(start_instr), 
         .D(instr_active), .Z(n9)) /* synthesis lut_function=(!(A+!((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(155[17] 157[20])
    defparam i21898_4_lut.init = 16'h5551;
    LUT4 i1_3_lut (.A(data_txn_len[0]), .B(data_txn_len[1]), .C(qspi_data_byte_idx[1]), 
         .Z(n21854)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C)))) */ ;
    defparam i1_3_lut.init = 16'h4141;
    LUT4 i1_2_lut_rep_517 (.A(mem_data_ready), .B(data_txn_len[1]), .Z(n25253)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_517.init = 16'h2222;
    LUT4 i52_2_lut_rep_656 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n25392)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i52_2_lut_rep_656.init = 16'hbbbb;
    LUT4 i1_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(qspi_data_ready), .D(n8888), .Z(clk_c_enable_142)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (D)+!B !(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h4f00;
    LUT4 i12097_2_lut_rep_657 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n25393)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12097_2_lut_rep_657.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_446 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(qspi_data_ready), .D(n8888), .Z(clk_c_enable_134)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i1_3_lut_4_lut_adj_446.init = 16'h8f00;
    LUT4 instr_data_7__I_148_i1_3_lut (.A(data_to_write[0]), .B(instr_data[8]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1700[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_148_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_447 (.A(instr_active), .B(\addr[24] ), .Z(n21878)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_447.init = 16'h4444;
    LUT4 i1_2_lut_rep_667 (.A(\addr[24] ), .B(instr_active), .Z(n25403)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_2_lut_rep_667.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_adj_448 (.A(\addr[24] ), .B(instr_active), .C(\addr_in[23] ), 
         .D(start_instr), .Z(spi_ram_a_select_N_2040)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_3_lut_4_lut_adj_448.init = 16'hfffd;
    LUT4 i1_4_lut_adj_449 (.A(n25325), .B(debug_stop_txn_N_1850), .C(is_writing), 
         .D(spi_clk_pos), .Z(stop_txn_now_N_2094)) /* synthesis lut_function=(A (B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(91[18] 99[12])
    defparam i1_4_lut_adj_449.init = 16'h8808;
    PFUMX debug_stop_txn_I_157 (.BLUT(debug_stop_txn_N_1851), .ALUT(debug_stop_txn_N_1873), 
          .C0(instr_active), .Z(debug_stop_txn_N_1850)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;
    LUT4 i1_4_lut_adj_450 (.A(n25272), .B(\next_instr_write_offset[3] ), 
         .C(n1), .D(n4_c), .Z(debug_stall_txn)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_450.init = 16'h0400;
    LUT4 qspi_data_byte_idx_1__I_0_197_i3_2_lut_rep_678 (.A(qspi_data_byte_idx[0]), 
         .B(qspi_data_byte_idx[1]), .Z(n25414)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam qspi_data_byte_idx_1__I_0_197_i3_2_lut_rep_678.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_451 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(qspi_data_ready), .D(instr_active), .Z(n4_c)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam i1_2_lut_3_lut_4_lut_adj_451.init = 16'h0200;
    LUT4 i21780_2_lut_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n8888), .D(qspi_data_ready), .Z(clk_c_enable_150)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam i21780_2_lut_3_lut_4_lut.init = 16'h20f0;
    LUT4 i1_2_lut_rep_625_3_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(instr_active), .Z(n25361)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam i1_2_lut_rep_625_3_lut.init = 16'h2020;
    LUT4 qspi_data_byte_idx_1__I_0_i3_2_lut_rep_687 (.A(qspi_data_byte_idx[0]), 
         .B(qspi_data_byte_idx[1]), .Z(n25423)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[144:171])
    defparam qspi_data_byte_idx_1__I_0_i3_2_lut_rep_687.init = 16'heeee;
    LUT4 i6931_3_lut (.A(data_to_write[31]), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6931_3_lut.init = 16'hcaca;
    LUT4 i6933_3_lut (.A(data_to_write[30]), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6933_3_lut.init = 16'hcaca;
    LUT4 i6935_3_lut (.A(data_to_write[29]), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6935_3_lut.init = 16'hcaca;
    LUT4 i6937_3_lut (.A(data_to_write[28]), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6937_3_lut.init = 16'hcaca;
    LUT4 i6939_3_lut (.A(data_to_write[27]), .B(instr_data[11]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6939_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_628_3_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(data_stall), .Z(n25364)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[144:171])
    defparam i1_2_lut_rep_628_3_lut.init = 16'h1010;
    LUT4 i1_3_lut_4_lut_adj_452 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(qspi_data_ready), .D(n8888), .Z(clk_c_enable_157)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[144:171])
    defparam i1_3_lut_4_lut_adj_452.init = 16'h1f00;
    LUT4 i10102_4_lut (.A(data_to_write[26]), .B(instr_data[10]), .C(qspi_data_ready), 
         .D(n25393), .Z(instr_data_7__N_1700[26])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i10102_4_lut.init = 16'hca0a;
    LUT4 i10104_4_lut (.A(data_to_write[25]), .B(instr_data[9]), .C(qspi_data_ready), 
         .D(n25393), .Z(instr_data_7__N_1700[25])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i10104_4_lut.init = 16'hca0a;
    LUT4 i10091_4_lut (.A(data_to_write[24]), .B(instr_data[8]), .C(qspi_data_ready), 
         .D(n25393), .Z(instr_data_7__N_1700[24])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i10091_4_lut.init = 16'hca0a;
    LUT4 i6941_3_lut (.A(data_to_write[23]), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6941_3_lut.init = 16'hcaca;
    LUT4 i6943_3_lut (.A(data_to_write[22]), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6943_3_lut.init = 16'hcaca;
    LUT4 i6945_3_lut (.A(data_to_write[21]), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6945_3_lut.init = 16'hcaca;
    LUT4 i6947_3_lut (.A(data_to_write[20]), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6947_3_lut.init = 16'hcaca;
    LUT4 i6949_3_lut (.A(data_to_write[19]), .B(instr_data[11]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6949_3_lut.init = 16'hcaca;
    LUT4 i10100_4_lut (.A(data_to_write[18]), .B(instr_data[10]), .C(qspi_data_ready), 
         .D(n25392), .Z(instr_data_7__N_1700[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i10100_4_lut.init = 16'h0aca;
    LUT4 i10098_4_lut (.A(data_to_write[17]), .B(instr_data[9]), .C(qspi_data_ready), 
         .D(n25392), .Z(instr_data_7__N_1700[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i10098_4_lut.init = 16'h0aca;
    LUT4 i10096_4_lut (.A(data_to_write[16]), .B(instr_data[8]), .C(qspi_data_ready), 
         .D(n25392), .Z(instr_data_7__N_1700[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i10096_4_lut.init = 16'h0aca;
    LUT4 i6951_3_lut (.A(data_to_write[15]), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6951_3_lut.init = 16'hcaca;
    LUT4 i6953_3_lut (.A(data_to_write[14]), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6953_3_lut.init = 16'hcaca;
    LUT4 i6955_3_lut (.A(data_to_write[13]), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6955_3_lut.init = 16'hcaca;
    LUT4 i6957_3_lut (.A(data_to_write[12]), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6957_3_lut.init = 16'hcaca;
    LUT4 i6959_3_lut (.A(data_to_write[11]), .B(instr_data[11]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6959_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_148_i11_4_lut (.A(data_to_write[10]), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n25414), .Z(instr_data_7__N_1700[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_148_i11_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_148_i10_4_lut (.A(data_to_write[9]), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n25414), .Z(instr_data_7__N_1700[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_148_i10_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_148_i9_4_lut (.A(data_to_write[8]), .B(instr_data[8]), 
         .C(qspi_data_ready), .D(n25414), .Z(instr_data_7__N_1700[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_148_i9_4_lut.init = 16'h0aca;
    LUT4 i6961_3_lut (.A(data_to_write[7]), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6961_3_lut.init = 16'hcaca;
    LUT4 i6963_3_lut (.A(data_to_write[6]), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6963_3_lut.init = 16'hcaca;
    LUT4 i6965_3_lut (.A(data_to_write[5]), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6965_3_lut.init = 16'hcaca;
    LUT4 i6967_3_lut (.A(data_to_write[4]), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1700[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i6967_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_148_i4_4_lut (.A(data_to_write[3]), .B(instr_data[11]), 
         .C(qspi_data_ready), .D(n25423), .Z(instr_data_7__N_1700[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_148_i4_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_148_i3_4_lut (.A(data_to_write[2]), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n25423), .Z(instr_data_7__N_1700[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_148_i3_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_148_i2_4_lut (.A(data_to_write[1]), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n25423), .Z(instr_data_7__N_1700[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_148_i2_4_lut.init = 16'h0aca;
    LUT4 i1_3_lut_4_lut_adj_453 (.A(qspi_data_ready), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(start_instr), .D(n25286), .Z(clk_c_enable_26)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[26:60])
    defparam i1_3_lut_4_lut_adj_453.init = 16'hfeff;
    LUT4 i20751_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[28]), .D(\mem_data_from_read[20] ), .Z(n23026)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20751_3_lut_4_lut.init = 16'hf960;
    LUT4 i20741_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[9]), .D(instr_data[1]), .Z(n23016)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20741_3_lut_4_lut.init = 16'hf960;
    LUT4 i20738_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(\qspi_data_buf[8] ), .D(instr_data[0]), .Z(n23013)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20738_3_lut_4_lut.init = 16'hf960;
    LUT4 i20739_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[24]), .D(\mem_data_from_read[16] ), .Z(n23014)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20739_3_lut_4_lut.init = 16'hf960;
    LUT4 i20744_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(\qspi_data_buf[10] ), .D(instr_data[2]), .Z(n23019)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20744_3_lut_4_lut.init = 16'hf960;
    LUT4 i20745_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[26]), .D(\mem_data_from_read[18] ), .Z(n23020)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20745_3_lut_4_lut.init = 16'hf960;
    LUT4 i20747_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[11]), .D(instr_data[3]), .Z(n23022)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20747_3_lut_4_lut.init = 16'hf960;
    LUT4 i20756_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(\qspi_data_buf[14] ), .D(instr_data[6]), .Z(n23031)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20756_3_lut_4_lut.init = 16'hf960;
    LUT4 i20754_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(\qspi_data_buf[29] ), .D(\mem_data_from_read[21] ), .Z(n23029)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20754_3_lut_4_lut.init = 16'hf960;
    LUT4 i20757_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[30]), .D(\mem_data_from_read[22] ), .Z(n23032)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20757_3_lut_4_lut.init = 16'hf960;
    LUT4 i20760_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[31]), .D(\mem_data_from_read[23] ), .Z(n23035)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20760_3_lut_4_lut.init = 16'hf960;
    LUT4 n14378_bdd_3_lut_22107_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(\qspi_data_buf[25] ), .D(\mem_data_from_read[17] ), .Z(n24195)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n14378_bdd_3_lut_22107_4_lut.init = 16'hf960;
    LUT4 i4434_4_lut (.A(n25275), .B(continue_txn_N_1862), .C(continue_txn), 
         .D(data_stall_N_1889), .Z(clk_c_enable_193)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(198[22] 203[16])
    defparam i4434_4_lut.init = 16'h05c5;
    LUT4 i20748_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[27]), .D(\mem_data_from_read[19] ), .Z(n23023)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20748_3_lut_4_lut.init = 16'hf960;
    LUT4 i20759_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[15]), .D(instr_data[7]), .Z(n23034)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20759_3_lut_4_lut.init = 16'hf960;
    LUT4 i20750_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(\qspi_data_buf[12] ), .D(instr_data[4]), .Z(n23025)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20750_3_lut_4_lut.init = 16'hf960;
    LUT4 i20753_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_1752[0]), 
         .C(qspi_data_buf[13]), .D(instr_data[5]), .Z(n23028)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i20753_3_lut_4_lut.init = 16'hf960;
    LUT4 i1_4_lut_adj_454 (.A(mem_data_ready), .B(n25364), .C(n25342), 
         .D(n25340), .Z(continue_txn_N_1862)) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C (D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i1_4_lut_adj_454.init = 16'h0c4c;
    LUT4 i3618_3_lut (.A(qspi_data_byte_idx[1]), .B(qspi_data_byte_idx[0]), 
         .C(write_qspi_data_byte_idx_1__N_1752[0]), .Z(write_qspi_data_byte_idx[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i3618_3_lut.init = 16'h6a6a;
    LUT4 i2_2_lut_4_lut (.A(n25321), .B(n25302), .C(rst_reg_n), .D(start_instr), 
         .Z(qspi_data_byte_idx_1__N_1756)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i2_2_lut_4_lut.init = 16'hff7f;
    LUT4 i21794_2_lut_3_lut_4_lut (.A(n25342), .B(n25320), .C(rst_reg_n), 
         .D(n25321), .Z(clk_c_enable_43)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(71[15:31])
    defparam i21794_2_lut_3_lut_4_lut.init = 16'h1fff;
    LUT4 i1_2_lut_rep_423_3_lut_4_lut (.A(n25342), .B(n25320), .C(start_instr), 
         .D(n25321), .Z(n25159)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(71[15:31])
    defparam i1_2_lut_rep_423_3_lut_4_lut.init = 16'hf1ff;
    LUT4 i1_3_lut_rep_550_4_lut (.A(n25342), .B(n25320), .C(rst_reg_n), 
         .D(n25321), .Z(n25286)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(71[15:31])
    defparam i1_3_lut_rep_550_4_lut.init = 16'he000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_455 (.A(n25325), .B(n25324), .C(n21878), 
         .D(n25161), .Z(addr_in[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(95[18] 98[33])
    defparam i1_2_lut_3_lut_4_lut_adj_455.init = 16'he0f0;
    LUT4 i3287_2_lut (.A(continue_txn), .B(rst_reg_n), .Z(n5278)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i3287_2_lut.init = 16'h4444;
    LUT4 i2_2_lut_rep_568_4_lut (.A(n25370), .B(n17512), .C(n25432), .D(n25325), 
         .Z(n25304)) /* synthesis lut_function=(A (D)+!A (((D)+!C)+!B)) */ ;
    defparam i2_2_lut_rep_568_4_lut.init = 16'hff15;
    LUT4 i1_2_lut_rep_566_3_lut_4_lut (.A(n25371), .B(qspi_write_done), 
         .C(n25342), .D(n25340), .Z(n25302)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(75[13:41])
    defparam i1_2_lut_rep_566_3_lut_4_lut.init = 16'hfeff;
    LUT4 i12122_2_lut_rep_539_3_lut_4_lut_3_lut_4_lut (.A(n25371), .B(qspi_write_done), 
         .C(n25342), .D(n25340), .Z(n25275)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(75[13:41])
    defparam i12122_2_lut_rep_539_3_lut_4_lut_3_lut_4_lut.init = 16'hfeee;
    LUT4 i11602_4_lut (.A(qspi_data_byte_idx[1]), .B(txn_len[0]), .C(qspi_data_byte_idx[0]), 
         .D(\txn_len[1] ), .Z(n174[1])) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(155[17] 157[20])
    defparam i11602_4_lut.init = 16'h581a;
    LUT4 i1_3_lut_adj_456 (.A(instr_active), .B(start_instr), .C(data_txn_len[0]), 
         .Z(txn_len[0])) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_3_lut_adj_456.init = 16'hfefe;
    PFUMX i22543 (.BLUT(n25470), .ALUT(n25471), .C0(fsm_state[0]), .Z(n25472));
    qspi_controller q_ctrl (.n24335(n24335), .n1032(n1032), .clk_c(clk_c), 
            .n25154(n25154), .\addr_in[24] (addr_in[24]), .spi_ram_a_select_N_2040(spi_ram_a_select_N_2040), 
            .spi_ram_b_select_N_2044(spi_ram_b_select_N_2044), .spi_clk_pos(spi_clk_pos), 
            .is_writing(is_writing), .clk_c_enable_103(clk_c_enable_103), 
            .n23082(n23082), .\instr_data[8] (instr_data[8]), .n17515(n17515), 
            .fsm_state({fsm_state}), .n25174(n25174), .n25384(n25384), 
            .\read_cycles_count[1] (read_cycles_count[1]), .debug_stall_txn(debug_stall_txn), 
            .data_stall(data_stall), .n25355(n25355), .n21746(n21746), 
            .n23019(n23019), .n23020(n23020), .\write_qspi_data_byte_idx[1] (write_qspi_data_byte_idx[1]), 
            .n25151(n25151), .n25371(n25371), .n25470(n25470), .n23029(n23029), 
            .clk_c_enable_354(clk_c_enable_354), .qspi_data_ready(qspi_data_ready), 
            .n6595(n6595), .\write_qspi_data_byte_idx_1__N_1752[0] (write_qspi_data_byte_idx_1__N_1752[0]), 
            .n23022(n23022), .n23023(n23023), .\instr_data[13] (instr_data[13]), 
            .\instr_data[11] (instr_data[11]), .\instr_data[10] (instr_data[10]), 
            .n23013(n23013), .n23014(n23014), .n25150(n25150), .n57(n57), 
            .n18783(n18783), .n25159(n25159), .\instr_data[9] (instr_data[9]), 
            .\instr_data[12] (instr_data[12]), .\instr_data[14] (instr_data[14]), 
            .\instr_data[15] (instr_data[15]), .debug_stop_txn_N_1850(debug_stop_txn_N_1850), 
            .qspi_write_done(qspi_write_done), .rst_reg_n(rst_reg_n), .n6611(n6611), 
            .clk_c_enable_52(clk_c_enable_52), .n24195(n24195), .n25472(n25472), 
            .n23025(n23025), .n23028(n23028), .n23031(n23031), .n23034(n23034), 
            .n9278(n9278), .n25353(n25353), .n25342(n25342), .n25320(n25320), 
            .n8888(n8888), .start_instr(start_instr), .\addr_in[23] (\addr_in[23] ), 
            .\addr[24] (\addr[24] ), .instr_active(instr_active), .stop_txn_now_N_2094(stop_txn_now_N_2094), 
            .n5(n5), .n25170(n25170), .n334(n333[1]), .next_bit(next_bit), 
            .n25252(n25252), .uart_txd_N_2327(uart_txd_N_2327), .clk_c_enable_397(clk_c_enable_397), 
            .n22788(n22788), .n20638(n20638), .n25334(n25334), .clk_c_enable_208(clk_c_enable_208), 
            .n4(n4), .clk_c_enable_322(clk_c_enable_322), .\qv_data_read_n[1] (\qv_data_read_n[1] ), 
            .\qv_data_write_n[1] (\qv_data_write_n[1] ), .n25370(n25370), 
            .n20731(n20731), .n19413(n19413), .n25324(n25324), .n8460(n8460), 
            .instr_active_N_1837(instr_active_N_1837), .n23016(n23016), 
            .n25325(n25325), .n1002(n1002), .n26(n26), .n25172(n25172), 
            .n23032(n23032), .n23035(n23035), .n23026(n23026)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(112[21] 136[6])
    
endmodule
//
// Verilog Description of module qspi_controller
//

module qspi_controller (n24335, n1032, clk_c, n25154, \addr_in[24] , 
            spi_ram_a_select_N_2040, spi_ram_b_select_N_2044, spi_clk_pos, 
            is_writing, clk_c_enable_103, n23082, \instr_data[8] , n17515, 
            fsm_state, n25174, n25384, \read_cycles_count[1] , debug_stall_txn, 
            data_stall, n25355, n21746, n23019, n23020, \write_qspi_data_byte_idx[1] , 
            n25151, n25371, n25470, n23029, clk_c_enable_354, qspi_data_ready, 
            n6595, \write_qspi_data_byte_idx_1__N_1752[0] , n23022, n23023, 
            \instr_data[13] , \instr_data[11] , \instr_data[10] , n23013, 
            n23014, n25150, n57, n18783, n25159, \instr_data[9] , 
            \instr_data[12] , \instr_data[14] , \instr_data[15] , debug_stop_txn_N_1850, 
            qspi_write_done, rst_reg_n, n6611, clk_c_enable_52, n24195, 
            n25472, n23025, n23028, n23031, n23034, n9278, n25353, 
            n25342, n25320, n8888, start_instr, \addr_in[23] , \addr[24] , 
            instr_active, stop_txn_now_N_2094, n5, n25170, n334, next_bit, 
            n25252, uart_txd_N_2327, clk_c_enable_397, n22788, n20638, 
            n25334, clk_c_enable_208, n4, clk_c_enable_322, \qv_data_read_n[1] , 
            \qv_data_write_n[1] , n25370, n20731, n19413, n25324, 
            n8460, instr_active_N_1837, n23016, n25325, n1002, n26, 
            n25172, n23032, n23035, n23026) /* synthesis syn_module_defined=1 */ ;
    input n24335;
    output n1032;
    input clk_c;
    output n25154;
    input \addr_in[24] ;
    input spi_ram_a_select_N_2040;
    input spi_ram_b_select_N_2044;
    output spi_clk_pos;
    output is_writing;
    output clk_c_enable_103;
    input n23082;
    output \instr_data[8] ;
    output n17515;
    output [2:0]fsm_state;
    input n25174;
    output n25384;
    output \read_cycles_count[1] ;
    input debug_stall_txn;
    input data_stall;
    output n25355;
    output n21746;
    input n23019;
    input n23020;
    input \write_qspi_data_byte_idx[1] ;
    input n25151;
    output n25371;
    output n25470;
    input n23029;
    input clk_c_enable_354;
    output qspi_data_ready;
    output n6595;
    output \write_qspi_data_byte_idx_1__N_1752[0] ;
    input n23022;
    input n23023;
    output \instr_data[13] ;
    output \instr_data[11] ;
    output \instr_data[10] ;
    input n23013;
    input n23014;
    input n25150;
    input n57;
    output n18783;
    input n25159;
    output \instr_data[9] ;
    output \instr_data[12] ;
    output \instr_data[14] ;
    output \instr_data[15] ;
    input debug_stop_txn_N_1850;
    input qspi_write_done;
    input rst_reg_n;
    output n6611;
    output clk_c_enable_52;
    input n24195;
    input n25472;
    input n23025;
    input n23028;
    input n23031;
    input n23034;
    output n9278;
    output n25353;
    input n25342;
    input n25320;
    output n8888;
    input start_instr;
    input \addr_in[23] ;
    input \addr[24] ;
    input instr_active;
    input stop_txn_now_N_2094;
    output n5;
    input n25170;
    input n334;
    input next_bit;
    input n25252;
    input uart_txd_N_2327;
    output clk_c_enable_397;
    input n22788;
    input n20638;
    input n25334;
    output clk_c_enable_208;
    input n4;
    output clk_c_enable_322;
    input \qv_data_read_n[1] ;
    input \qv_data_write_n[1] ;
    input n25370;
    output n20731;
    input n19413;
    input n25324;
    output n8460;
    output instr_active_N_1837;
    input n23016;
    output n25325;
    output n1002;
    output n26;
    input n25172;
    input n23032;
    input n23035;
    input n23026;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n24339, n24340, spi_flash_select, clk_c_enable_83, spi_ram_a_select, 
        spi_ram_b_select, clk_c_enable_95, n21503, clk_c_enable_358;
    wire [7:0]data_out_7__N_1908;
    
    wire stop_txn_reg, stop_txn_reg_N_2091, clk_c_enable_282, n1024;
    wire [1:0]read_cycles_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(105[15:32])
    
    wire n1110;
    wire [1:0]n381;
    wire [1:0]n181;
    
    wire n20659, n25454, n25453, n13909, n26601, clk_c_enable_313;
    wire [1:0]n396;
    wire [3:0]spi_in_buffer;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(91[15:28])
    
    wire clk_c_enable_191, n23083, n21516, n25314;
    wire [55:0]instr_data_15__N_1690;
    wire [2:0]nibbles_remaining;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(86[15:32])
    
    wire n1033, data_ready_N_2069, last_ram_a_sel, last_ram_b_sel, n21583, 
        data_req_N_2049, n26600, n25400;
    wire [2:0]n4050;
    
    wire n14434, n25399, n25313, n25330, n25335, n25398, n9023, 
        n1026, n25455, n24196, n24193, n23363, n25356, n26602, 
        clk_c_enable_355, n25149;
    wire [1:0]n127;
    
    wire n8776, n25437, debug_stop_txn, n21820, n24194, n25374, 
        n25386, n22716;
    wire [7:0]data_out_7__N_2004;
    
    wire n23275, n22304, n25345, n25312, n25385, n24310, n4_c, 
        n21734, n21704, n5366, n21722, n5368;
    wire [2:0]n356;
    
    wire n21262, n9, n26599, n21840, n24192, n25303, n21501;
    
    PFUMX i22051 (.BLUT(n24339), .ALUT(n24335), .C0(n1032), .Z(n24340));
    FD1P3JX spi_flash_select_227 (.D(\addr_in[24] ), .SP(clk_c_enable_83), 
            .PD(n25154), .CK(clk_c), .Q(spi_flash_select)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_flash_select_227.GSR = "DISABLED";
    FD1P3JX spi_ram_a_select_228 (.D(spi_ram_a_select_N_2040), .SP(clk_c_enable_83), 
            .PD(n25154), .CK(clk_c), .Q(spi_ram_a_select)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_ram_a_select_228.GSR = "DISABLED";
    FD1P3JX spi_ram_b_select_229 (.D(spi_ram_b_select_N_2044), .SP(clk_c_enable_83), 
            .PD(n25154), .CK(clk_c), .Q(spi_ram_b_select)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_ram_b_select_229.GSR = "DISABLED";
    FD1P3AX spi_clk_pos_225 (.D(n21503), .SP(clk_c_enable_95), .CK(clk_c), 
            .Q(spi_clk_pos)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_clk_pos_225.GSR = "DISABLED";
    FD1P3IX is_writing_222 (.D(n23082), .SP(clk_c_enable_103), .CD(n25154), 
            .CK(clk_c), .Q(is_writing)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam is_writing_222.GSR = "DISABLED";
    FD1P3AX data_i1 (.D(data_out_7__N_1908[0]), .SP(clk_c_enable_358), .CK(clk_c), 
            .Q(\instr_data[8] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i1.GSR = "DISABLED";
    FD1S3IX stop_txn_reg_218 (.D(stop_txn_reg_N_2091), .CK(clk_c), .CD(n17515), 
            .Q(stop_txn_reg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(98[12] 103[8])
    defparam stop_txn_reg_218.GSR = "DISABLED";
    FD1P3IX fsm_state__i0 (.D(n1024), .SP(clk_c_enable_282), .CD(n25154), 
            .CK(clk_c), .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i0.GSR = "DISABLED";
    LUT4 mux_114_i1_4_lut_4_lut (.A(read_cycles_count[0]), .B(n25174), .C(n1110), 
         .D(n25384), .Z(n381[0])) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam mux_114_i1_4_lut_4_lut.init = 16'h5c50;
    LUT4 i11689_2_lut_3_lut_4_lut_4_lut (.A(read_cycles_count[0]), .B(\read_cycles_count[1] ), 
         .C(debug_stall_txn), .D(data_stall), .Z(n181[0])) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam i11689_2_lut_3_lut_4_lut_4_lut.init = 16'h5554;
    LUT4 i1_3_lut_4_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[0]), .C(fsm_state[2]), 
         .D(n25355), .Z(n21746)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+(C+(D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h0021;
    LUT4 n23019_bdd_4_lut (.A(n23019), .B(n23020), .C(\write_qspi_data_byte_idx[1] ), 
         .D(n20659), .Z(data_out_7__N_1908[2])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n23019_bdd_4_lut.init = 16'hca00;
    LUT4 mux_113_i3_4_lut_then_4_lut (.A(n25355), .B(fsm_state[2]), .C(fsm_state[1]), 
         .D(fsm_state[0]), .Z(n25454)) /* synthesis lut_function=(A (B (C (D)))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_113_i3_4_lut_then_4_lut.init = 16'hd454;
    LUT4 mux_113_i3_4_lut_else_4_lut (.A(n25355), .B(fsm_state[2]), .C(fsm_state[1]), 
         .D(fsm_state[0]), .Z(n25453)) /* synthesis lut_function=(A (B (C (D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_113_i3_4_lut_else_4_lut.init = 16'hd444;
    LUT4 i1_3_lut_4_lut (.A(n25151), .B(clk_c_enable_103), .C(n25371), 
         .D(n25154), .Z(clk_c_enable_95)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i1_3_lut_4_lut.init = 16'hfff8;
    LUT4 fsm_state_0__bdd_4_lut_22764 (.A(fsm_state[0]), .B(fsm_state[2]), 
         .C(fsm_state[1]), .D(is_writing), .Z(n13909)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam fsm_state_0__bdd_4_lut_22764.init = 16'h7f77;
    LUT4 i1_3_lut_3_lut_4_lut_then_4_lut (.A(fsm_state[0]), .B(fsm_state[1]), 
         .C(spi_clk_pos), .D(fsm_state[2]), .Z(n26601)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (D)))) */ ;
    defparam i1_3_lut_3_lut_4_lut_then_4_lut.init = 16'h6400;
    FD1P3IX read_cycles_count__i0 (.D(n396[0]), .SP(clk_c_enable_313), .CD(n25154), 
            .CK(clk_c), .Q(read_cycles_count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam read_cycles_count__i0.GSR = "DISABLED";
    LUT4 n24336_bdd_3_lut_rep_432_4_lut_else_4_lut_4_lut (.A(is_writing), 
         .B(spi_flash_select), .C(fsm_state[1]), .D(fsm_state[2]), .Z(n25470)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam n24336_bdd_3_lut_rep_432_4_lut_else_4_lut_4_lut.init = 16'hf010;
    FD1P3AX spi_in_buffer__i1 (.D(n23083), .SP(clk_c_enable_191), .CK(clk_c), 
            .Q(spi_in_buffer[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer__i1.GSR = "DISABLED";
    LUT4 i21455_3_lut (.A(n23029), .B(n21516), .C(n25314), .Z(instr_data_15__N_1690[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(238[18] 244[12])
    defparam i21455_3_lut.init = 16'hcaca;
    FD1P3IX nibbles_remaining__i0 (.D(n1033), .SP(clk_c_enable_354), .CD(n25154), 
            .CK(clk_c), .Q(nibbles_remaining[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i0.GSR = "DISABLED";
    FD1S3IX data_ready_224 (.D(data_ready_N_2069), .CK(clk_c), .CD(n6595), 
            .Q(qspi_data_ready)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam data_ready_224.GSR = "DISABLED";
    FD1S3JX last_ram_a_sel_235 (.D(spi_ram_a_select), .CK(clk_c), .PD(n17515), 
            .Q(last_ram_a_sel)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(272[12] 280[8])
    defparam last_ram_a_sel_235.GSR = "DISABLED";
    FD1S3JX last_ram_b_sel_236 (.D(spi_ram_b_select), .CK(clk_c), .PD(n17515), 
            .Q(last_ram_b_sel)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(272[12] 280[8])
    defparam last_ram_b_sel_236.GSR = "DISABLED";
    FD1S3IX data_req_230 (.D(data_req_N_2049), .CK(clk_c), .CD(n21583), 
            .Q(\write_qspi_data_byte_idx_1__N_1752[0] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam data_req_230.GSR = "DISABLED";
    LUT4 i1_3_lut_3_lut_4_lut_else_4_lut (.A(fsm_state[0]), .B(fsm_state[1]), 
         .C(spi_clk_pos), .D(fsm_state[2]), .Z(n26600)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;
    defparam i1_3_lut_3_lut_4_lut_else_4_lut.init = 16'hf4f0;
    LUT4 n23022_bdd_4_lut (.A(n23022), .B(n23023), .C(\write_qspi_data_byte_idx[1] ), 
         .D(n20659), .Z(data_out_7__N_1908[3])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n23022_bdd_4_lut.init = 16'hca00;
    LUT4 i21832_3_lut_4_lut (.A(n25400), .B(nibbles_remaining[0]), .C(n1032), 
         .D(n4050[1]), .Z(n14434)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam i21832_3_lut_4_lut.init = 16'h0d02;
    LUT4 mux_2546_i3_3_lut_4_lut (.A(fsm_state[2]), .B(n25399), .C(n25355), 
         .D(nibbles_remaining[2]), .Z(n4050[2])) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(180[37:57])
    defparam mux_2546_i3_3_lut_4_lut.init = 16'hf101;
    LUT4 i728_2_lut_rep_577_3_lut_4_lut (.A(fsm_state[2]), .B(n25399), .C(spi_clk_pos), 
         .D(n25355), .Z(n25313)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A ((D)+!C)) */ ;
    defparam i728_2_lut_rep_577_3_lut_4_lut.init = 16'hdf0f;
    LUT4 i1_3_lut_4_lut_adj_424 (.A(fsm_state[2]), .B(n25399), .C(is_writing), 
         .D(n25355), .Z(data_req_N_2049)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_424.init = 16'h0020;
    FD1P3AX data_i6 (.D(data_out_7__N_1908[5]), .SP(clk_c_enable_358), .CK(clk_c), 
            .Q(\instr_data[13] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i6.GSR = "DISABLED";
    FD1P3AX data_i4 (.D(data_out_7__N_1908[3]), .SP(clk_c_enable_358), .CK(clk_c), 
            .Q(\instr_data[11] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i4.GSR = "DISABLED";
    FD1P3AX data_i3 (.D(data_out_7__N_1908[2]), .SP(clk_c_enable_358), .CK(clk_c), 
            .Q(\instr_data[10] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i3.GSR = "DISABLED";
    LUT4 n23013_bdd_4_lut (.A(n23013), .B(n23014), .C(\write_qspi_data_byte_idx[1] ), 
         .D(n20659), .Z(data_out_7__N_1908[0])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n23013_bdd_4_lut.init = 16'hca00;
    LUT4 i1_2_lut_rep_594_3_lut_4_lut (.A(nibbles_remaining[0]), .B(n25400), 
         .C(n25399), .D(fsm_state[2]), .Z(n25330)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_2_lut_rep_594_3_lut_4_lut.init = 16'he0ee;
    LUT4 i1_2_lut_rep_599_3_lut_4_lut (.A(nibbles_remaining[0]), .B(n25400), 
         .C(n25399), .D(fsm_state[2]), .Z(n25335)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_2_lut_rep_599_3_lut_4_lut.init = 16'h0e00;
    LUT4 i1_3_lut_4_lut_adj_425 (.A(fsm_state[2]), .B(n25398), .C(is_writing), 
         .D(fsm_state[0]), .Z(n9023)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[102:126])
    defparam i1_3_lut_4_lut_adj_425.init = 16'hf2f0;
    FD1P3IX fsm_state__i1 (.D(n24340), .SP(clk_c_enable_282), .CD(n25154), 
            .CK(clk_c), .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i1.GSR = "DISABLED";
    FD1P3IX fsm_state__i2 (.D(n1026), .SP(clk_c_enable_282), .CD(n25154), 
            .CK(clk_c), .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i2.GSR = "DISABLED";
    LUT4 i11992_3_lut_4_lut (.A(n25150), .B(n25371), .C(n57), .D(n25455), 
         .Z(n1026)) /* synthesis lut_function=(A (B ((D)+!C))+!A ((D)+!C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i11992_3_lut_4_lut.init = 16'hdd0d;
    L6MUX21 i21970 (.D0(n24196), .D1(n24193), .SD(n23363), .Z(data_out_7__N_1908[1]));
    LUT4 i21_4_lut (.A(n25356), .B(n26602), .C(is_writing), .D(fsm_state[0]), 
         .Z(clk_c_enable_355)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i21_4_lut.init = 16'hc5c0;
    FD1P3IX read_cycles_count__i1 (.D(n396[1]), .SP(clk_c_enable_313), .CD(n25154), 
            .CK(clk_c), .Q(\read_cycles_count[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam read_cycles_count__i1.GSR = "DISABLED";
    LUT4 i4787_rep_413_3_lut_4_lut (.A(n18783), .B(n25159), .C(n25371), 
         .D(clk_c_enable_103), .Z(n25149)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i4787_rep_413_3_lut_4_lut.init = 16'h0800;
    LUT4 i12232_2_lut (.A(read_cycles_count[0]), .B(\read_cycles_count[1] ), 
         .Z(n127[1])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(151[22:69])
    defparam i12232_2_lut.init = 16'h8888;
    FD1P3IX nibbles_remaining__i1 (.D(n14434), .SP(clk_c_enable_354), .CD(n25154), 
            .CK(clk_c), .Q(nibbles_remaining[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i1.GSR = "DISABLED";
    FD1P3IX nibbles_remaining__i2 (.D(n8776), .SP(clk_c_enable_354), .CD(n25154), 
            .CK(clk_c), .Q(nibbles_remaining[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i2.GSR = "DISABLED";
    FD1P3AX data_i2 (.D(data_out_7__N_1908[1]), .SP(clk_c_enable_355), .CK(clk_c), 
            .Q(\instr_data[9] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i2.GSR = "DISABLED";
    FD1P3AX data_i5 (.D(data_out_7__N_1908[4]), .SP(clk_c_enable_358), .CK(clk_c), 
            .Q(\instr_data[12] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i5.GSR = "DISABLED";
    FD1P3AX data_i7 (.D(data_out_7__N_1908[6]), .SP(clk_c_enable_358), .CK(clk_c), 
            .Q(\instr_data[14] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i7.GSR = "DISABLED";
    FD1P3AX data_i8 (.D(data_out_7__N_1908[7]), .SP(clk_c_enable_358), .CK(clk_c), 
            .Q(\instr_data[15] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i8.GSR = "DISABLED";
    LUT4 i11498_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n25437), .C(debug_stop_txn_N_1850), 
         .D(qspi_write_done), .Z(debug_stop_txn)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(180[37:57])
    defparam i11498_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i21755_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(n25437), .C(rst_reg_n), 
         .D(qspi_write_done), .Z(n6611)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(180[37:57])
    defparam i21755_2_lut_3_lut_4_lut.init = 16'h0f1f;
    LUT4 i1_3_lut_4_lut_adj_426 (.A(fsm_state[2]), .B(n25437), .C(debug_stop_txn), 
         .D(rst_reg_n), .Z(clk_c_enable_52)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(180[37:57])
    defparam i1_3_lut_4_lut_adj_426.init = 16'hf1ff;
    LUT4 i1_3_lut_4_lut_adj_427 (.A(fsm_state[2]), .B(n25437), .C(stop_txn_reg), 
         .D(spi_clk_pos), .Z(n21820)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(180[37:57])
    defparam i1_3_lut_4_lut_adj_427.init = 16'hfff1;
    PFUMX i21968 (.BLUT(n24195), .ALUT(n24194), .C0(n25314), .Z(n24196));
    LUT4 i8005_1_lut_rep_638 (.A(is_writing), .Z(n25374)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i8005_1_lut_rep_638.init = 16'h5555;
    LUT4 i1_4_lut_4_lut (.A(is_writing), .B(spi_flash_select), .C(fsm_state[0]), 
         .D(n25386), .Z(n22716)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_4_lut_4_lut.init = 16'h00f4;
    LUT4 n10254_bdd_3_lut_22467_4_lut_4_lut (.A(is_writing), .B(n57), .C(n25355), 
         .D(n25472), .Z(n24339)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam n10254_bdd_3_lut_22467_4_lut_4_lut.init = 16'h1d11;
    LUT4 mux_180_i5_3_lut_3_lut (.A(is_writing), .B(\instr_data[8] ), .C(n23025), 
         .Z(data_out_7__N_2004[4])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i5_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i6_3_lut_3_lut (.A(is_writing), .B(\instr_data[9] ), .C(n23028), 
         .Z(data_out_7__N_2004[5])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i6_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i7_3_lut_3_lut (.A(is_writing), .B(\instr_data[10] ), .C(n23031), 
         .Z(data_out_7__N_2004[6])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i7_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i8_3_lut_3_lut (.A(is_writing), .B(\instr_data[11] ), .C(n23034), 
         .Z(data_out_7__N_2004[7])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i8_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_rep_648 (.A(fsm_state[2]), .B(fsm_state[0]), .Z(n25384)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_648.init = 16'h8888;
    LUT4 i21935_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(n25400), 
         .D(nibbles_remaining[0]), .Z(n23275)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i21935_2_lut_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_3_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(data_stall), 
         .Z(n22304)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h0808;
    LUT4 equal_118_i4_2_lut_rep_650 (.A(fsm_state[1]), .B(fsm_state[2]), 
         .Z(n25386)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(183[42:63])
    defparam equal_118_i4_2_lut_rep_650.init = 16'hdddd;
    LUT4 i7014_1_lut (.A(\write_qspi_data_byte_idx_1__N_1752[0] ), .Z(n9278)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i7014_1_lut.init = 16'h5555;
    LUT4 equal_118_i5_2_lut_rep_609_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(fsm_state[0]), .Z(n25345)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(183[42:63])
    defparam equal_118_i5_2_lut_rep_609_3_lut.init = 16'hfdfd;
    LUT4 i1_2_lut_rep_617_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[0]), 
         .Z(n25353)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_617_3_lut.init = 16'h8080;
    LUT4 i3_3_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(\read_cycles_count[1] ), 
         .D(read_cycles_count[0]), .Z(clk_c_enable_191)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0080;
    LUT4 i11480_2_lut_rep_662 (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .Z(n25398)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11480_2_lut_rep_662.init = 16'heeee;
    LUT4 i27_3_lut_4_lut (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .C(n13909), .D(spi_clk_pos), .Z(n25312)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam i27_3_lut_4_lut.init = 16'hf101;
    LUT4 equal_3124_i8_2_lut_rep_620_3_lut (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .C(fsm_state[2]), .Z(n25356)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam equal_3124_i8_2_lut_rep_620_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_663 (.A(fsm_state[1]), .B(fsm_state[0]), .Z(n25399)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[102:126])
    defparam i1_2_lut_rep_663.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_649_3_lut (.A(fsm_state[1]), .B(fsm_state[0]), .C(fsm_state[2]), 
         .Z(n25385)) /* synthesis lut_function=(!(A (B (C))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[102:126])
    defparam i1_2_lut_rep_649_3_lut.init = 16'h3b3b;
    LUT4 fsm_state_1__bdd_4_lut_4_lut_3_lut (.A(fsm_state[1]), .B(fsm_state[0]), 
         .C(fsm_state[2]), .Z(n24310)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[102:126])
    defparam fsm_state_1__bdd_4_lut_4_lut_3_lut.init = 16'h2121;
    LUT4 equal_113_i4_2_lut_rep_664 (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .Z(n25400)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam equal_113_i4_2_lut_rep_664.init = 16'heeee;
    LUT4 equal_113_i5_2_lut_rep_619_3_lut (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .C(nibbles_remaining[0]), .Z(n25355)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam equal_113_i5_2_lut_rep_619_3_lut.init = 16'hfefe;
    LUT4 i3653_2_lut_3_lut_4_lut (.A(nibbles_remaining[1]), .B(nibbles_remaining[2]), 
         .C(n4050[1]), .D(nibbles_remaining[0]), .Z(n4_c)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i3653_2_lut_3_lut_4_lut.init = 16'hfff1;
    LUT4 i1_4_lut (.A(qspi_data_ready), .B(data_stall), .C(n25342), .D(n25320), 
         .Z(n8888)) /* synthesis lut_function=(A+!(B (C)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_4_lut.init = 16'haeaf;
    LUT4 i1_4_lut_adj_428 (.A(n18783), .B(clk_c_enable_103), .C(n25159), 
         .D(n25371), .Z(n1032)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i1_4_lut_adj_428.init = 16'h0080;
    LUT4 i1_4_lut_adj_429 (.A(start_instr), .B(\addr_in[23] ), .C(\addr[24] ), 
         .D(n21734), .Z(n18783)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(109[49:72])
    defparam i1_4_lut_adj_429.init = 16'hffef;
    LUT4 i1_2_lut (.A(instr_active), .B(last_ram_a_sel), .Z(n21734)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(109[49:72])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_430 (.A(start_instr), .B(\addr_in[23] ), .C(\addr[24] ), 
         .D(n21704), .Z(clk_c_enable_103)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_430.init = 16'hffbf;
    LUT4 i1_2_lut_adj_431 (.A(instr_active), .B(last_ram_b_sel), .Z(n21704)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_431.init = 16'heeee;
    LUT4 i21895_4_lut (.A(rst_reg_n), .B(stop_txn_now_N_2094), .C(n21820), 
         .D(n5), .Z(n21503)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i21895_4_lut.init = 16'h0200;
    LUT4 i1_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[0]), 
         .Z(n5)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_3_lut.init = 16'hf7f7;
    LUT4 i2803_3_lut_4_lut (.A(n25151), .B(clk_c_enable_103), .C(n25371), 
         .D(n25170), .Z(n5366)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i2803_3_lut_4_lut.init = 16'h08f8;
    PFUMX mux_129_i1 (.BLUT(n181[0]), .ALUT(n381[0]), .C0(n5), .Z(n396[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 i1_3_lut_adj_432 (.A(debug_stop_txn), .B(stop_txn_now_N_2094), 
         .C(stop_txn_reg), .Z(stop_txn_reg_N_2091)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut_adj_432.init = 16'h0202;
    LUT4 i1_4_lut_adj_433 (.A(n25154), .B(n21722), .C(n5368), .D(n25149), 
         .Z(clk_c_enable_282)) /* synthesis lut_function=(A+(B (C (D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(123[13:34])
    defparam i1_4_lut_adj_433.init = 16'hfaba;
    LUT4 i1_4_lut_adj_434 (.A(n5), .B(n25353), .C(n25170), .D(n25355), 
         .Z(n21722)) /* synthesis lut_function=(!(A (B+!(D))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_434.init = 16'h3200;
    LUT4 i2802_4_lut (.A(n25312), .B(n5366), .C(n25371), .D(n5), .Z(n5368)) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i2802_4_lut.init = 16'haccc;
    LUT4 mux_622_i1_4_lut (.A(n356[0]), .B(\addr_in[24] ), .C(n1032), 
         .D(n57), .Z(n1024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam mux_622_i1_4_lut.init = 16'hcacf;
    PFUMX i12246 (.BLUT(n334), .ALUT(n127[1]), .C0(n21262), .Z(n396[1]));
    LUT4 i23_3_lut_4_lut_4_lut_4_lut (.A(fsm_state[0]), .B(n25345), .C(spi_flash_select), 
         .D(is_writing), .Z(n9)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(180[37:57])
    defparam i23_3_lut_4_lut_4_lut_4_lut.init = 16'h7745;
    LUT4 i1_2_lut_rep_707 (.A(is_writing), .B(spi_flash_select), .Z(n26599)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_rep_707.init = 16'heeee;
    LUT4 i1_3_lut_rep_418_3_lut (.A(rst_reg_n), .B(stop_txn_reg), .C(stop_txn_now_N_2094), 
         .Z(n25154)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_3_lut_rep_418_3_lut.init = 16'hfdfd;
    LUT4 n14378_bdd_2_lut_22106_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(n25355), 
         .C(n25399), .D(fsm_state[2]), .Z(n24194)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam n14378_bdd_2_lut_22106_3_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 i1_4_lut_rep_484_4_lut (.A(rst_reg_n), .B(next_bit), .C(n25252), 
         .D(uart_txd_N_2327), .Z(clk_c_enable_397)) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_rep_484_4_lut.init = 16'hfdf5;
    LUT4 i1_4_lut_4_lut_adj_435 (.A(rst_reg_n), .B(n22788), .C(n20638), 
         .D(n25334), .Z(clk_c_enable_208)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_435.init = 16'hd555;
    LUT4 i1_2_lut_1_lut_1_lut (.A(rst_reg_n), .Z(n17515)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_2_lut_1_lut_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_2_lut (.A(rst_reg_n), .B(n4), .Z(clk_c_enable_322)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut_adj_436 (.A(rst_reg_n), .B(stop_txn_reg), .C(n25371), 
         .D(stop_txn_now_N_2094), .Z(clk_c_enable_313)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_436.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_437 (.A(rst_reg_n), .B(\qv_data_read_n[1] ), 
         .C(\qv_data_write_n[1] ), .D(n25370), .Z(n20731)) /* synthesis lut_function=((B (C+(D))+!B (D))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_437.init = 16'hffd5;
    LUT4 i1_4_lut_4_lut_adj_438 (.A(rst_reg_n), .B(stop_txn_reg), .C(stop_txn_now_N_2094), 
         .D(n25371), .Z(n6595)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_438.init = 16'hfdff;
    LUT4 i1_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n1032), .C(stop_txn_reg), 
         .D(stop_txn_now_N_2094), .Z(clk_c_enable_83)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_2_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_439 (.A(rst_reg_n), .B(n21840), .C(stop_txn_now_N_2094), 
         .D(n25312), .Z(n21583)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_4_lut_4_lut_adj_439.init = 16'hfffd;
    PFUMX mux_113_i1 (.BLUT(n9), .ALUT(n19413), .C0(n23275), .Z(n356[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 n23016_bdd_4_lut_22105_4_lut (.A(rst_reg_n), .B(spi_in_buffer[1]), 
         .C(n25399), .D(n25356), .Z(n24192)) /* synthesis lut_function=(A (B (C+(D)))+!A (B+!(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam n23016_bdd_4_lut_22105_4_lut.init = 16'hccc5;
    LUT4 i20808_4_lut_4_lut (.A(rst_reg_n), .B(fsm_state[0]), .C(is_writing), 
         .D(spi_in_buffer[1]), .Z(n23083)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D)+!B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i20808_4_lut_4_lut.init = 16'hfd01;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(n25324), .C(qspi_write_done), 
         .D(n25371), .Z(n8460)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 rstn_N_1760_I_0_2_lut_2_lut (.A(rst_reg_n), .B(debug_stop_txn), 
         .Z(instr_active_N_1837)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(85[13:19])
    defparam rstn_N_1760_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i21829_2_lut_4_lut (.A(n25313), .B(n25314), .C(is_writing), .D(n9023), 
         .Z(clk_c_enable_358)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;
    defparam i21829_2_lut_4_lut.init = 16'h7f00;
    LUT4 i21911_3_lut (.A(is_writing), .B(n25314), .C(\write_qspi_data_byte_idx[1] ), 
         .Z(n23363)) /* synthesis lut_function=(!(A (B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(238[18] 244[12])
    defparam i21911_3_lut.init = 16'h5757;
    PFUMX i21966 (.BLUT(n23016), .ALUT(n24192), .C0(n25374), .Z(n24193));
    LUT4 i1_2_lut_rep_701 (.A(fsm_state[0]), .B(fsm_state[1]), .Z(n25437)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_rep_701.init = 16'heeee;
    LUT4 i1_2_lut_rep_635_3_lut (.A(fsm_state[0]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .Z(n25371)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_rep_635_3_lut.init = 16'hfefe;
    LUT4 qspi_busy_I_0_2_lut_rep_589_3_lut_4_lut (.A(fsm_state[0]), .B(fsm_state[1]), 
         .C(qspi_write_done), .D(fsm_state[2]), .Z(n25325)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam qspi_busy_I_0_2_lut_rep_589_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut_3_lut_4_lut_2_lut_3_lut (.A(fsm_state[0]), .B(fsm_state[1]), 
         .C(fsm_state[2]), .Z(n1002)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i2_2_lut_3_lut_4_lut_2_lut_3_lut.init = 16'h1010;
    LUT4 i2_2_lut_4_lut (.A(n1002), .B(n25174), .C(n25384), .D(n25303), 
         .Z(n1110)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;
    defparam i2_2_lut_4_lut.init = 16'hff35;
    LUT4 i29_4_lut (.A(n25150), .B(n25312), .C(n25371), .D(n5), .Z(n26)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i29_4_lut.init = 16'hca0a;
    LUT4 i11704_4_lut (.A(nibbles_remaining[0]), .B(n1032), .C(n25400), 
         .D(n24310), .Z(n1033)) /* synthesis lut_function=(A (B)+!A (B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i11704_4_lut.init = 16'hdcdd;
    LUT4 i1_4_lut_adj_440 (.A(is_writing), .B(n25170), .C(n21501), .D(n5), 
         .Z(data_ready_N_2069)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_440.init = 16'h5011;
    LUT4 i1_4_lut_adj_441 (.A(n25312), .B(debug_stall_txn), .C(n25355), 
         .D(n22304), .Z(n21501)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_441.init = 16'h0200;
    LUT4 i1_4_lut_adj_442 (.A(fsm_state[0]), .B(stop_txn_reg), .C(fsm_state[1]), 
         .D(fsm_state[2]), .Z(n21840)) /* synthesis lut_function=(A (B)+!A (B+(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam i1_4_lut_adj_442.init = 16'hdccd;
    LUT4 i1_2_lut_4_lut (.A(n25355), .B(n5), .C(n25313), .D(is_writing), 
         .Z(n20659)) /* synthesis lut_function=(!(A (B+!(D))+!A (B (C+!(D))+!B !(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h3700;
    LUT4 i1_3_lut_4_lut_adj_443 (.A(n25355), .B(n25312), .C(n5), .D(n25172), 
         .Z(n21262)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_443.init = 16'hbfff;
    LUT4 i1_2_lut_rep_567_4_lut (.A(spi_clk_pos), .B(n25398), .C(n13909), 
         .D(n25355), .Z(n25303)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[25:140])
    defparam i1_2_lut_rep_567_4_lut.init = 16'hff5c;
    LUT4 i1_3_lut_4_lut_adj_444 (.A(n25330), .B(spi_clk_pos), .C(\instr_data[9] ), 
         .D(n25335), .Z(n21516)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_3_lut_4_lut_adj_444.init = 16'h4000;
    PFUMX i23143 (.BLUT(n26600), .ALUT(n26601), .C0(n25355), .Z(n26602));
    PFUMX data_out_7__I_0_242_i8 (.BLUT(instr_data_15__N_1690[31]), .ALUT(data_out_7__N_2004[7]), 
          .C0(n23363), .Z(data_out_7__N_1908[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i7 (.BLUT(instr_data_15__N_1690[30]), .ALUT(data_out_7__N_2004[6]), 
          .C0(n23363), .Z(data_out_7__N_1908[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i6 (.BLUT(instr_data_15__N_1690[29]), .ALUT(data_out_7__N_2004[5]), 
          .C0(n23363), .Z(data_out_7__N_1908[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i5 (.BLUT(instr_data_15__N_1690[28]), .ALUT(data_out_7__N_2004[4]), 
          .C0(n23363), .Z(data_out_7__N_1908[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 i21457_3_lut_4_lut (.A(\instr_data[10] ), .B(n25335), .C(n25314), 
         .D(n23032), .Z(instr_data_15__N_1690[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam i21457_3_lut_4_lut.init = 16'h8f80;
    LUT4 i21459_3_lut_4_lut (.A(\instr_data[11] ), .B(n25335), .C(n25314), 
         .D(n23035), .Z(instr_data_15__N_1690[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam i21459_3_lut_4_lut.init = 16'h8f80;
    LUT4 i21453_3_lut_4_lut (.A(\instr_data[8] ), .B(n25335), .C(n25314), 
         .D(n23026), .Z(instr_data_15__N_1690[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam i21453_3_lut_4_lut.init = 16'h8f80;
    LUT4 i12154_3_lut_rep_578_3_lut (.A(n25355), .B(n5), .C(spi_clk_pos), 
         .Z(n25314)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam i12154_3_lut_rep_578_3_lut.init = 16'h8c8c;
    LUT4 mux_2546_i2_4_lut (.A(n22716), .B(nibbles_remaining[1]), .C(n25355), 
         .D(n25385), .Z(n4050[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_2546_i2_4_lut.init = 16'hcac0;
    LUT4 mux_629_i3_4_lut (.A(n4050[2]), .B(\addr_in[24] ), .C(n1032), 
         .D(n4_c), .Z(n8776)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam mux_629_i3_4_lut.init = 16'h3a35;
    PFUMX i22533 (.BLUT(n25453), .ALUT(n25454), .C0(n26599), .Z(n25455));
    
endmodule
//
// Verilog Description of module tinyqv_cpu
//

module tinyqv_cpu (clk_c, instr_data, \pc[10] , \pc[11] , qv_data_read_n, 
            \pc[12] , VCC_net, debug_instr_valid, n25370, n24935, 
            \mem_data_from_read[4] , counter_hi, \pc[13] , n24929, \mem_data_from_read[6] , 
            \instr_len[2] , instr_fetch_running, \pc[14] , \pc[1] , 
            addr, \pc[2] , \pc[3] , \pc[4] , \pc[5] , \pc[6] , \pc[7] , 
            \instr_write_offset[3] , \next_instr_write_offset[3] , rst_reg_n, 
            n25175, n2015, n2010, \data_from_read[2] , n8229, \gpio_out_sel[7] , 
            n1949, n1969, n26612, instr_complete_N_1378, n21541, n8146, 
            \qspi_data_buf[25] , \qspi_data_buf[29] , qspi_data_ready, 
            n25361, \mem_data_from_read[17] , \mem_data_from_read[21] , 
            debug_data_continue, n3597, data_to_write, \pc[15] , qv_data_write_n, 
            \pc[16] , \mem_data_from_read[27] , \mem_data_from_read[31] , 
            \pc[17] , instr_fetch_running_N_676, debug_stall_txn, n21800, 
            \next_pc_for_core[3] , \next_pc_for_core[7] , \pc[18] , \imm[19] , 
            \imm[23] , n17512, \imm[11] , \imm[15] , \imm[3] , \imm[7] , 
            \imm[18] , \imm[22] , n25363, \imm[10] , \imm[14] , \imm[2] , 
            \imm[6] , \imm[17] , \imm[21] , \imm[9] , \imm[13] , \imm[1] , 
            \imm[5] , mem_op_increment_reg, n23084, \imm[16] , \imm[20] , 
            \imm[8] , \imm[12] , \imm[4] , \next_pc_for_core[4] , \pc[9] , 
            \next_pc_for_core[9] , \next_pc_for_core[13] , \pc[19] , n10, 
            n22566, \pc[20] , \pc[8] , n25163, n25161, \instr_avail_len[3] , 
            \next_pc_for_core[8] , \next_pc_for_core[12] , n25194, n25336, 
            clk_c_enable_206, \next_pc_for_core[5] , \next_pc_for_core[6] , 
            \next_pc_for_core[10] , \next_pc_for_core[11] , n25417, \next_pc_for_core[14] , 
            \next_pc_for_core[15] , \next_pc_for_core[16] , \next_pc_for_core[17] , 
            \next_pc_for_core[18] , \next_pc_for_core[19] , \next_pc_for_core[20] , 
            \next_pc_for_core[21] , \next_pc_for_core[22] , data_txn_len, 
            \qspi_data_buf[14] , n25253, \pc[21] , \pc[22] , \pc[23] , 
            \next_pc_for_core[23] , \qspi_data_buf[10] , n25419, \mem_data_from_read[19] , 
            \mem_data_from_read[23] , n25431, n25432, n25324, n20582, 
            \mem_data_from_read[16] , \mem_data_from_read[20] , \mem_data_from_read[18] , 
            \mem_data_from_read[22] , \mem_data_from_read[3] , read_en, 
            \qspi_data_buf[12] , \instr_addr_23__N_49[22] , \early_branch_addr[23] , 
            \instr_addr[23] , instr_fetch_stopped, \early_branch_addr[5] , 
            \early_branch_addr[4] , \early_branch_addr[2] , \early_branch_addr[6] , 
            \early_branch_addr[3] , \early_branch_addr[7] , \early_branch_addr[8] , 
            \early_branch_addr[9] , \early_branch_addr[10] , \early_branch_addr[11] , 
            \early_branch_addr[12] , \early_branch_addr[13] , \early_branch_addr[14] , 
            \early_branch_addr[15] , \early_branch_addr[16] , \early_branch_addr[17] , 
            \early_branch_addr[18] , \early_branch_addr[19] , \early_branch_addr[20] , 
            \early_branch_addr[21] , \early_branch_addr[22] , \qspi_data_buf[8] , 
            n25304, instr_active, \txn_len[1] , n8527, n25403, \addr_in[23] , 
            spi_ram_b_select_N_2044, n23037, n23038, n1, n22873, \mem_data_from_read[1] , 
            \mem_data_from_read[5] , \mem_data_from_read[9] , \mem_data_from_read[13] , 
            n25272, n22334, n25337, \mem_data_from_read[24] , \mem_data_from_read[28] , 
            \mem_data_from_read[26] , \mem_data_from_read[30] , mem_data_ready, 
            \data_from_read[6] , \data_from_read[0] , start_instr, n24998, 
            mem_op_increment_reg_de, n25273, clk_c_enable_27, \next_fsm_state_3__N_2230[3] , 
            \cycle[0] , \ui_in_sync[1] , n1092, debug_rd, accum, d_3__N_1599, 
            \mul_out[1] , \mul_out[3] , n14111, n24186, \mul_out[2] , 
            \next_accum[6] , \next_accum[7] , \next_accum[8] , \next_accum[9] , 
            \next_accum[10] , \next_accum[11] , \next_accum[12] , \next_accum[13] , 
            \next_accum[14] , \next_accum[15] , GND_net, \next_accum[16] , 
            \next_accum[17] , \next_accum[18] , \next_accum[19] , \next_accum[5] , 
            \next_accum[4] ) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    input [15:0]instr_data;
    output \pc[10] ;
    output \pc[11] ;
    output [1:0]qv_data_read_n;
    output \pc[12] ;
    input VCC_net;
    output debug_instr_valid;
    input n25370;
    input n24935;
    input \mem_data_from_read[4] ;
    output [4:2]counter_hi;
    output \pc[13] ;
    input n24929;
    input \mem_data_from_read[6] ;
    output \instr_len[2] ;
    output instr_fetch_running;
    output \pc[14] ;
    output \pc[1] ;
    output [27:0]addr;
    output \pc[2] ;
    output \pc[3] ;
    output \pc[4] ;
    output \pc[5] ;
    output \pc[6] ;
    output \pc[7] ;
    output \instr_write_offset[3] ;
    output \next_instr_write_offset[3] ;
    input rst_reg_n;
    output n25175;
    output n2015;
    output n2010;
    input \data_from_read[2] ;
    input n8229;
    input \gpio_out_sel[7] ;
    input n1949;
    input n1969;
    input n26612;
    output instr_complete_N_1378;
    output n21541;
    output n8146;
    input \qspi_data_buf[25] ;
    input \qspi_data_buf[29] ;
    input qspi_data_ready;
    input n25361;
    input \mem_data_from_read[17] ;
    input \mem_data_from_read[21] ;
    output debug_data_continue;
    output n3597;
    output [31:0]data_to_write;
    output \pc[15] ;
    output [1:0]qv_data_write_n;
    output \pc[16] ;
    input \mem_data_from_read[27] ;
    input \mem_data_from_read[31] ;
    output \pc[17] ;
    input instr_fetch_running_N_676;
    input debug_stall_txn;
    output n21800;
    input \next_pc_for_core[3] ;
    input \next_pc_for_core[7] ;
    output \pc[18] ;
    output \imm[19] ;
    output \imm[23] ;
    output n17512;
    output \imm[11] ;
    output \imm[15] ;
    output \imm[3] ;
    output \imm[7] ;
    output \imm[18] ;
    output \imm[22] ;
    output n25363;
    output \imm[10] ;
    output \imm[14] ;
    output \imm[2] ;
    output \imm[6] ;
    output \imm[17] ;
    output \imm[21] ;
    output \imm[9] ;
    output \imm[13] ;
    output \imm[1] ;
    output \imm[5] ;
    output mem_op_increment_reg;
    input n23084;
    output \imm[16] ;
    output \imm[20] ;
    output \imm[8] ;
    output \imm[12] ;
    output \imm[4] ;
    input \next_pc_for_core[4] ;
    output \pc[9] ;
    input \next_pc_for_core[9] ;
    input \next_pc_for_core[13] ;
    output \pc[19] ;
    input n10;
    output n22566;
    output \pc[20] ;
    output \pc[8] ;
    output n25163;
    output n25161;
    input \instr_avail_len[3] ;
    input \next_pc_for_core[8] ;
    input \next_pc_for_core[12] ;
    input n25194;
    input n25336;
    output clk_c_enable_206;
    input \next_pc_for_core[5] ;
    input \next_pc_for_core[6] ;
    input \next_pc_for_core[10] ;
    input \next_pc_for_core[11] ;
    input n25417;
    input \next_pc_for_core[14] ;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[16] ;
    input \next_pc_for_core[17] ;
    input \next_pc_for_core[18] ;
    input \next_pc_for_core[19] ;
    input \next_pc_for_core[20] ;
    input \next_pc_for_core[21] ;
    input \next_pc_for_core[22] ;
    input [1:0]data_txn_len;
    input \qspi_data_buf[14] ;
    input n25253;
    output \pc[21] ;
    output \pc[22] ;
    output \pc[23] ;
    input \next_pc_for_core[23] ;
    input \qspi_data_buf[10] ;
    output n25419;
    input \mem_data_from_read[19] ;
    input \mem_data_from_read[23] ;
    input n25431;
    output n25432;
    output n25324;
    output n20582;
    input \mem_data_from_read[16] ;
    input \mem_data_from_read[20] ;
    input \mem_data_from_read[18] ;
    input \mem_data_from_read[22] ;
    input \mem_data_from_read[3] ;
    output read_en;
    input \qspi_data_buf[12] ;
    input \instr_addr_23__N_49[22] ;
    input \early_branch_addr[23] ;
    output \instr_addr[23] ;
    input instr_fetch_stopped;
    input \early_branch_addr[5] ;
    input \early_branch_addr[4] ;
    input \early_branch_addr[2] ;
    input \early_branch_addr[6] ;
    input \early_branch_addr[3] ;
    input \early_branch_addr[7] ;
    input \early_branch_addr[8] ;
    input \early_branch_addr[9] ;
    input \early_branch_addr[10] ;
    input \early_branch_addr[11] ;
    input \early_branch_addr[12] ;
    input \early_branch_addr[13] ;
    input \early_branch_addr[14] ;
    input \early_branch_addr[15] ;
    input \early_branch_addr[16] ;
    input \early_branch_addr[17] ;
    input \early_branch_addr[18] ;
    input \early_branch_addr[19] ;
    input \early_branch_addr[20] ;
    input \early_branch_addr[21] ;
    input \early_branch_addr[22] ;
    input \qspi_data_buf[8] ;
    input n25304;
    input instr_active;
    output \txn_len[1] ;
    input n8527;
    input n25403;
    input \addr_in[23] ;
    output spi_ram_b_select_N_2044;
    input n23037;
    input n23038;
    output n1;
    output n22873;
    input \mem_data_from_read[1] ;
    input \mem_data_from_read[5] ;
    input \mem_data_from_read[9] ;
    input \mem_data_from_read[13] ;
    output n25272;
    output n22334;
    input n25337;
    input \mem_data_from_read[24] ;
    input \mem_data_from_read[28] ;
    input \mem_data_from_read[26] ;
    input \mem_data_from_read[30] ;
    input mem_data_ready;
    input \data_from_read[6] ;
    input \data_from_read[0] ;
    output start_instr;
    input n24998;
    output mem_op_increment_reg_de;
    output n25273;
    input clk_c_enable_27;
    input \next_fsm_state_3__N_2230[3] ;
    output \cycle[0] ;
    input \ui_in_sync[1] ;
    output n1092;
    output [3:0]debug_rd;
    output [15:0]accum;
    output [19:0]d_3__N_1599;
    input \mul_out[1] ;
    input \mul_out[3] ;
    output n14111;
    input n24186;
    input \mul_out[2] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input GND_net;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[5] ;
    input \next_accum[4] ;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [15:0]n2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire clk_c_enable_219, is_store, clk_c_enable_203, n25424, is_store_de, 
        data_ready_latch, clk_c_enable_15, n21632, is_load, is_load_de;
    wire [3:0]alu_op;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    
    wire clk_c_enable_84;
    wire [3:0]alu_op_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(64[16:25])
    wire [15:0]n1629;
    wire [15:0]n1649;
    
    wire n25338;
    wire [31:0]instr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(47[17:22])
    wire [3:0]alu_op_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[16:25])
    
    wire n24943, n24942, n26597, n19, clk_c_enable_29;
    wire [63:0]instr_data_0__15__N_369;
    
    wire n24940, n24939, n25284, n24941, clk_c_enable_393;
    wire [20:0]pc_23__N_642;
    wire [3:0]rd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(119[15:17])
    
    wire clk_c_enable_312;
    wire [3:0]n3675;
    wire [15:0]n7;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire clk_c_enable_72;
    wire [2:1]instr_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(113[15:24])
    
    wire clk_c_enable_38, n25219;
    wire [2:0]mem_op;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(115[15:21])
    
    wire clk_c_enable_69;
    wire [2:0]mem_op_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(65[16:25])
    wire [3:0]rs1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(117[15:18])
    wire [3:0]n2089;
    
    wire clk_c_enable_56, n21389;
    wire [15:0]n9;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire clk_c_enable_93;
    wire [22:0]instr_addr_23__N_49;
    wire [2:0]instr_write_offset_3__N_665;
    wire [2:0]additional_mem_ops;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(120[15:33])
    wire [2:0]additional_mem_ops_2__N_480;
    
    wire load_started, clk_c_enable_54, n54, clk_c_enable_110, debug_instr_valid_N_167, 
        n21388, n24937, n24933, n24938, n24936, clk_c_enable_74, 
        n24931, n24927, n24932, clk_c_enable_91, n24930;
    wire [1:0]instr_len_2__N_307;
    
    wire was_early_branch, clk_c_enable_197, was_early_branch_N_759, is_branch, 
        is_branch_de, clk_c_enable_102, n5438, interrupt_core, n25179, 
        data_ready_sync, data_ready_core, is_alu_imm, is_alu_imm_de, 
        n24915, n24914, n24916;
    wire [1:0]pc_2__N_663;
    
    wire clk_c_enable_309;
    wire [27:0]addr_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(131[17:25])
    wire [3:0]rs2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(118[15:18])
    wire [3:0]n1729;
    wire [15:0]n14;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire clk_c_enable_216, is_auipc, is_auipc_de, n25407, n20739;
    wire [3:2]addr_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(121[15:26])
    wire [1:0]n17;
    
    wire n25207, n24876, n3615, n24877, n25434, is_alu_reg, is_alu_reg_de, 
        n5599, n25178, n27, n25171, n3989, n21916, n25190, n25167, 
        n24997, n26598, n25279, n25005, n25451, n25450, n25164, 
        n10_c, n21067, n3619, n21297, clk_c_enable_368, n21750, 
        n7955, n8, n25457, n25456, n26, n22286, n35, n22, n22298;
    wire [31:0]n2937;
    
    wire n24568;
    wire [31:0]n2978;
    
    wire n25166, n23265, n21978, n16, n1943, n25468, n25467, n22050, 
        n6, n22056;
    wire [3:1]next_pc_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[16:30])
    
    wire n6830, n5879, n25221, n25015, n5856, n21390;
    wire [31:0]n2890;
    
    wire n25028, n25177, n25182, n22126, n3613, n3605;
    wire [31:0]n2703;
    wire [31:0]n2414;
    wire [31:0]n2854;
    
    wire n25155, n23237, n25209;
    wire [30:0]n4516;
    
    wire n25311, n25027, n25415, n21962, n25406, n21884, n25409, 
        n21970, n25030, n25029, n25031, n25394, n21966;
    wire [15:0]n1950;
    
    wire is_timer_addr, data_out_3__N_1116, n23106, n23062, load_top_bit;
    wire [59:0]debug_branch_N_571;
    
    wire n21369, n22272, n3993, n23059;
    wire [15:0]n1970;
    
    wire n25169, n25438, n25439, n25440, is_jalr, is_jalr_de, n22996, 
        clk_c_enable_194, data_continue_N_694, is_jal, is_jal_de, n22990, 
        clk_c_enable_324;
    wire [3:0]data_out_slice;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(230[16:30])
    
    wire n25372, no_write_in_progress, no_write_in_progress_N_202, n20805, 
        clk_c_enable_314;
    wire [1:0]data_write_n_1__N_100;
    
    wire n25156, n21236, n3611, n25290;
    wire [31:0]n2813;
    
    wire is_system, is_system_de, is_lui, is_lui_de, n25181, n25176, 
        n20762, n21402, n22028, n21322, n25281, n20641, n24, n23065;
    wire [3:0]n5047;
    wire [59:0]debug_rd_3__N_136;
    
    wire n25381, n6657;
    wire [59:0]debug_branch_N_177;
    
    wire any_additional_mem_ops, n25180;
    wire [2:0]n4030;
    
    wire n24486, n24487, n24419, n24420, n25237, n25244, n21944, 
        n23060;
    wire [3:0]timer_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(143[16:26])
    
    wire n8755, n22_adj_2374, n4, n25196, n22324, n22992, n20952, 
        instr_fetch_restart_N_678, n25118, n25153, n21121, n25266, 
        n25119, n23063, n8759;
    wire [12:0]n4548;
    
    wire n24422, n22994, n22092, n3991, n23073;
    wire [31:0]imm;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(100[16:19])
    
    wire n23444, n23443, n22959, n22970, n24424, n24425, n24428, 
        n24427, n23442, n23441, n24429, n23437, n23436, n25420, 
        n23435, n23434, n23430, n23429, n26596, n25248, n25203, 
        n25278, n24431, n24432, n25210, n26286, n23428, n22282, 
        n1945, n23427, clk_c_enable_209, n25383, n25326, n26288, 
        n23423, n22978, n23422, n23421, clk_c_enable_392, n23420, 
        clk_c_enable_218, n25249, n22074, n23055, n24999, n23057, 
        n22966, n22972, n22038, n22964, n22974, n24450, n22062, 
        n22957, n22968, n22852, n149, n24449, n22955, n23155, 
        n22944, n22953, n25226, n25265;
    wire [2:0]additional_mem_ops_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(70[16:37])
    
    wire n24452, n24453, n23068, n25264, n22961, n24457, n23403, 
        n23405, n22963, n22977, n209, n25359, n23245, n209_adj_2376;
    wire [3:0]data_rs1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(83[16:24])
    
    wire n25402;
    wire [59:0]debug_branch_N_173;
    
    wire n22941, n25288, n22960, n25287, n22962, n149_adj_2377, 
        n24687, n24686, n24688, n21430, n25458, n25144, n25240, 
        n25263, n21152, n21150, n21148, n24661, n24660, n24662, 
        n157, n25158, n23220;
    wire [23:1]return_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(135[17:28])
    
    wire debug_ret;
    wire [20:0]n1742;
    
    wire n25206;
    wire [31:0]n2736;
    wire [1:0]n699;
    
    wire n21499, n25307;
    wire [2:0]n17_adj_2394;
    
    wire n22470, n22172;
    wire [31:0]n2772;
    
    wire n22010;
    wire [15:0]n4608;
    wire [3:0]n1708;
    
    wire n66, n12257, n25387, n25004;
    wire [3:0]n155;
    
    wire n25216, n25239;
    wire [3:0]alu_op_3__N_901;
    
    wire n25444, n25445, cmp;
    wire [3:0]alu_b_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[16:24])
    wire [3:0]alu_a_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[16:24])
    
    wire n21812, n25267, n23899;
    wire [31:0]n2627;
    
    wire n21260, n22878, n25195, n25260, n24919, n21575, n22646, 
        n22648, n22644, n22636, n22622, n23900, n22638, n22620, 
        n21269;
    wire [3:0]n2075;
    
    wire n2244, n3603;
    wire [31:0]n2666;
    
    wire n25211, n32, n25442, n25255;
    wire [3:0]alu_op_3__N_1068;
    
    wire n15_adj_2380, n21157, n21242, n27_adj_2381, n25441, n25429, 
        n25368, n25418, n23070, n5570, n21248, n24488;
    wire [1:0]n1768;
    
    wire n23395;
    wire [3:0]n234;
    wire [3:0]debug_rd_3__N_1298;
    
    wire n21960, n21113, n21954, n24617, n24616, n24618, n23064, 
        n24564, n24565, n21374, n21375, n21376, n25258, n24566, 
        n8768, n25257, n15_adj_2382, n25, n23066, n13814, n37, 
        n23058, n23061, n21212, n3589, n23039, n8735, n25277, 
        clk_c_enable_328, clk_c_enable_332, clk_c_enable_336, clk_c_enable_340, 
        clk_c_enable_344, clk_c_enable_348, clk_c_enable_352;
    wire [3:0]n2047;
    
    wire n2242, n21153, n25375, n25348, n26610, n26608, n11558, 
        n20807, n22112, n20, is_ret_de, n25350, n25202, n25208, 
        n22098, n25289, n22954, n23341, n15_adj_2383, n25227, is_jalr_N_1101, 
        n25121, clk_c_enable_370, n22016, n11, n23271;
    wire [3:0]n2066;
    wire [3:0]n3657;
    wire [3:0]n3665;
    
    wire n20605, n23319, n25412, n23322, n22160, n25349, n2240, 
        n2236, n25410, n23111, n25411;
    wire [1:0]n4455;
    wire [3:0]n2034;
    wire [3:0]n2042;
    
    wire n22354, n13;
    wire [3:0]n1718;
    wire [3:0]n3631;
    
    wire n25236, n25222, is_lui_N_1096, n20720, n25247, n8_adj_2384, 
        n22044;
    wire [3:0]data_rs2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(84[16:24])
    wire [3:0]n92;
    
    wire n24567, n22068, n21303, n22080, n21992, n26287, n24615, 
        n7734, n25475, n23011, n23012, n7775;
    wire [3:0]n4994;
    wire [3:0]n5029;
    
    wire n25408;
    wire [16:0]mie;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(323[16:19])
    
    wire n5, n22798, instr_fetch_running_N_674, n22030;
    wire [3:0]n2052;
    wire [3:0]n3636;
    wire [20:0]n1143;
    
    wire n25310, n21594, n25230, n24956, n25191, n25443, n25225, 
        n21868, n21864;
    wire [3:0]n3641;
    
    wire n22976, n23255, n23089, n7375, n6647, n25197, n25421, 
        n6638, n23067, n8154, n25422, n22022, load_done, instr_complete_N_1382, 
        n23898, n22839, n23897, n24659, n23896, n20820, n25241, 
        n23895, n24489, n24229, n24228, n24230, n23894, n25426, 
        n22939, n225, n226, n24264, n24685, n225_adj_2385, n25228, 
        n25261, n25262, n25243, n29, n25234, n20650, n25430, n25343, 
        n25341, n23424, n23425, n25319, n23431, n23432, n23438, 
        n23439, n23445, n23446, n25301, n25369, n25300, n25282, 
        n25269;
    wire [6:0]cycle_count_wide;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(279[16:32])
    
    wire cy;
    wire [4:0]increment_result_3__N_1642;
    wire [3:0]instrret_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(301[16:30])
    
    wire instr_retired, cy_adj_2386;
    wire [4:0]increment_result_3__N_1656;
    
    wire n23069, n25294, n25256, n24451, n25152, n25229, n24913, 
        n25352, cy_adj_2387, n25218, n25231, cy_adj_2388, time_pulse_r, 
        n25305, n3, n212, n8761, n25259, n24423, n22290, n21860, 
        n13701, n25238, n25245, n24430, n25189, n24894, n23379, 
        n22008, n25214, n22384, n23166, n21910;
    wire [31:0]mtimecmp;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(30[16:24])
    
    wire mtimecmp_1__N_1672, mtimecmp_0__N_1674, mtimecmp_2__N_1670, n25232;
    wire [3:0]debug_branch_N_181;
    
    wire n21998, n23399, n23400, n23, n26_adj_2389, n25162, n22398, 
        n26289, n10_adj_2390, debug_rd_3__N_1306, n21898, n22178, 
        n22238, n22132;
    wire [2:0]n1764;
    
    wire n25120, n25365, mstatus_mpie, mstatus_mie;
    wire [3:0]csr_read_3__N_1170;
    
    wire n25212, n22214, n22226, n21696, n24875, n25016, n28, 
        n22202, n24_adj_2391, n21230, n22146, n22004, n22933, n16_adj_2392, 
        n25014;
    wire [3:0]mtime_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(29[16:25])
    
    wire n25329, n25291, n22558, n22254, n22258, n25333, n25293, 
        n25316, clk_c_enable_111, n25344, n25271;
    wire [3:0]tmp_data_in_3__N_1245;
    wire [5:0]mcause;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(325[15:21])
    
    wire mstatus_mte, mtimecmp_3__N_1666, clk_c_enable_205, timer_interrupt, 
        n5_adj_2393;
    wire [3:0]\reg_access[3] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(30[16:26])
    wire [3:0]\reg_access[4] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(30[16:26])
    
    wire n25246, clk_c_enable_170, n22086, n12, n22208, n22152, 
        n22867, n22232, n22244, n22184, n22120, n22138, n22276, 
        n22220;
    
    FD1P3AX instr_data_3__i47 (.D(instr_data[14]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i47.GSR = "DISABLED";
    FD1P3AX instr_data_3__i46 (.D(instr_data[13]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i46.GSR = "DISABLED";
    FD1P3AX instr_data_3__i45 (.D(instr_data[12]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i45.GSR = "DISABLED";
    FD1P3AX instr_data_3__i44 (.D(instr_data[11]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i44.GSR = "DISABLED";
    FD1P3AX instr_data_3__i43 (.D(instr_data[10]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i43.GSR = "DISABLED";
    FD1P3AX instr_data_3__i42 (.D(instr_data[9]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i42.GSR = "DISABLED";
    FD1P3AX instr_data_3__i41 (.D(instr_data[8]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i41.GSR = "DISABLED";
    FD1P3AX instr_data_3__i40 (.D(instr_data[7]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i40.GSR = "DISABLED";
    FD1P3IX is_store_396 (.D(is_store_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_store)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_store_396.GSR = "DISABLED";
    FD1P3AX instr_data_3__i39 (.D(instr_data[6]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i39.GSR = "DISABLED";
    FD1P3AX data_ready_latch_416 (.D(n21632), .SP(clk_c_enable_15), .CK(clk_c), 
            .Q(data_ready_latch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(235[12] 256[8])
    defparam data_ready_latch_416.GSR = "DISABLED";
    FD1P3IX is_load_393 (.D(is_load_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_load)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_load_393.GSR = "DISABLED";
    FD1P3AX instr_data_3__i38 (.D(instr_data[5]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i38.GSR = "DISABLED";
    FD1P3AX instr_data_3__i37 (.D(instr_data[4]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i37.GSR = "DISABLED";
    FD1P3AX instr_data_3__i36 (.D(instr_data[3]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i36.GSR = "DISABLED";
    FD1P3AX instr_data_3__i35 (.D(instr_data[2]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i35.GSR = "DISABLED";
    FD1P3IX alu_op__i3 (.D(alu_op_de[3]), .SP(clk_c_enable_84), .CD(n25424), 
            .CK(clk_c), .Q(alu_op[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i3.GSR = "DISABLED";
    PFUMX mux_1013_i12 (.BLUT(n1629[11]), .ALUT(n1649[11]), .C0(n25338), 
          .Z(instr[27]));
    FD1P3IX alu_op__i2 (.D(alu_op_de[2]), .SP(clk_c_enable_84), .CD(n25424), 
            .CK(clk_c), .Q(alu_op_in[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i2.GSR = "DISABLED";
    FD1P3IX alu_op__i0 (.D(alu_op_de[0]), .SP(clk_c_enable_84), .CD(n25424), 
            .CK(clk_c), .Q(alu_op[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i0.GSR = "DISABLED";
    PFUMX i22403 (.BLUT(n24943), .ALUT(n24942), .C0(n26597), .Z(n19));
    FD1P3AX instr_data_3__i34 (.D(instr_data_0__15__N_369[49]), .SP(clk_c_enable_29), 
            .CK(clk_c), .Q(n2[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i34.GSR = "DISABLED";
    FD1P3AX instr_data_3__i33 (.D(instr_data_0__15__N_369[0]), .SP(clk_c_enable_29), 
            .CK(clk_c), .Q(n2[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i33.GSR = "DISABLED";
    PFUMX i22400 (.BLUT(n24940), .ALUT(n24939), .C0(n25284), .Z(n24941));
    PFUMX mux_1013_i10 (.BLUT(n1629[9]), .ALUT(n1649[9]), .C0(n25338), 
          .Z(instr[25]));
    FD1P3IX pc_offset__i10 (.D(pc_23__N_642[7]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[10] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i10.GSR = "DISABLED";
    FD1P3IX pc_offset__i11 (.D(pc_23__N_642[8]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[11] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i11.GSR = "DISABLED";
    FD1P3AX rd_i0_i0 (.D(n3675[0]), .SP(clk_c_enable_312), .CK(clk_c), 
            .Q(rd[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i0.GSR = "DISABLED";
    FD1P3AX instr_data_3__i32 (.D(instr_data[15]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i32.GSR = "DISABLED";
    FD1P3AX instr_data_3__i31 (.D(instr_data[14]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i31.GSR = "DISABLED";
    FD1P3AX instr_data_3__i30 (.D(instr_data[13]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i30.GSR = "DISABLED";
    FD1P3IX instr_len_i1 (.D(n25219), .SP(clk_c_enable_38), .CD(n25424), 
            .CK(clk_c), .Q(instr_len[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_len_i1.GSR = "DISABLED";
    FD1P3AX instr_data_3__i29 (.D(instr_data[12]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i29.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i0 (.D(mem_op_de[0]), .SP(clk_c_enable_69), .CK(clk_c), 
            .Q(mem_op[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i0.GSR = "DISABLED";
    FD1P3AX rs1_i0_i0 (.D(n2089[0]), .SP(clk_c_enable_69), .CK(clk_c), 
            .Q(rs1[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i0.GSR = "DISABLED";
    FD1P3AX data_read_n_i0_i0 (.D(n21389), .SP(clk_c_enable_56), .CK(clk_c), 
            .Q(qv_data_read_n[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_read_n_i0_i0.GSR = "DISABLED";
    FD1P3AX instr_data_3__i28 (.D(instr_data[11]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i28.GSR = "DISABLED";
    FD1P3IX alu_op__i1 (.D(alu_op_de[1]), .SP(clk_c_enable_84), .CD(n25424), 
            .CK(clk_c), .Q(alu_op[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i1.GSR = "DISABLED";
    FD1P3AX instr_data_3__i27 (.D(instr_data[10]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i27.GSR = "DISABLED";
    FD1P3IX pc_offset__i12 (.D(pc_23__N_642[9]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[12] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i12.GSR = "DISABLED";
    FD1P3AX instr_data_3__i26 (.D(instr_data[9]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i26.GSR = "DISABLED";
    FD1P3AX instr_data_3__i1 (.D(instr_data_0__15__N_369[0]), .SP(clk_c_enable_93), 
            .CK(clk_c), .Q(n9[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i1.GSR = "DISABLED";
    FD1P3AX instr_data_3__i25 (.D(instr_data[8]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i25.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i1 (.D(instr_write_offset_3__N_665[0]), .CK(clk_c), 
            .CD(n25424), .Q(instr_addr_23__N_49[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i1.GSR = "DISABLED";
    PFUMX mux_1013_i9 (.BLUT(n1629[8]), .ALUT(n1649[8]), .C0(n25338), 
          .Z(instr[24]));
    FD1S3IX additional_mem_ops__i0 (.D(additional_mem_ops_2__N_480[0]), .CK(clk_c), 
            .CD(n25424), .Q(additional_mem_ops[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i0.GSR = "DISABLED";
    FD1P3IX load_started_422 (.D(VCC_net), .SP(clk_c_enable_54), .CD(n54), 
            .CK(clk_c), .Q(load_started)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam load_started_422.GSR = "DISABLED";
    FD1P3IX instr_valid_392 (.D(debug_instr_valid_N_167), .SP(clk_c_enable_110), 
            .CD(n25424), .CK(clk_c), .Q(debug_instr_valid)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_valid_392.GSR = "DISABLED";
    FD1P3AX data_read_n_i0_i1 (.D(n21388), .SP(clk_c_enable_56), .CK(clk_c), 
            .Q(qv_data_read_n[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_read_n_i0_i1.GSR = "DISABLED";
    PFUMX i22397 (.BLUT(n24937), .ALUT(n24933), .C0(n25370), .Z(n24938));
    PFUMX i22395 (.BLUT(n24935), .ALUT(\mem_data_from_read[4] ), .C0(counter_hi[2]), 
          .Z(n24936));
    FD1P3IX pc_offset__i13 (.D(pc_23__N_642[10]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[13] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i13.GSR = "DISABLED";
    FD1P3AX rs1_i0_i3 (.D(n2089[3]), .SP(clk_c_enable_69), .CK(clk_c), 
            .Q(rs1[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i3.GSR = "DISABLED";
    FD1P3AX instr_data_3__i24 (.D(instr_data[7]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i24.GSR = "DISABLED";
    FD1P3AX instr_data_3__i23 (.D(instr_data[6]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i23.GSR = "DISABLED";
    FD1P3AX rs1_i0_i2 (.D(n2089[2]), .SP(clk_c_enable_69), .CK(clk_c), 
            .Q(rs1[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i2.GSR = "DISABLED";
    FD1P3AX instr_data_3__i22 (.D(instr_data[5]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i22.GSR = "DISABLED";
    FD1P3AX rs1_i0_i1 (.D(n2089[1]), .SP(clk_c_enable_69), .CK(clk_c), 
            .Q(rs1[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i1.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i2 (.D(mem_op_de[2]), .SP(clk_c_enable_69), .CK(clk_c), 
            .Q(mem_op[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i2.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i1 (.D(mem_op_de[1]), .SP(clk_c_enable_69), .CK(clk_c), 
            .Q(mem_op[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i1.GSR = "DISABLED";
    FD1P3AX instr_data_3__i21 (.D(instr_data[4]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i21.GSR = "DISABLED";
    FD1P3AX instr_data_3__i20 (.D(instr_data[3]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i20.GSR = "DISABLED";
    FD1P3AX instr_data_3__i19 (.D(instr_data[2]), .SP(clk_c_enable_72), 
            .CK(clk_c), .Q(n7[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i19.GSR = "DISABLED";
    FD1P3AX instr_data_3__i18 (.D(instr_data_0__15__N_369[49]), .SP(clk_c_enable_74), 
            .CK(clk_c), .Q(n7[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i18.GSR = "DISABLED";
    PFUMX i22392 (.BLUT(n24931), .ALUT(n24927), .C0(n25370), .Z(n24932));
    FD1P3AX instr_data_3__i17 (.D(instr_data_0__15__N_369[0]), .SP(clk_c_enable_74), 
            .CK(clk_c), .Q(n7[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i17.GSR = "DISABLED";
    FD1P3AX instr_data_3__i16 (.D(instr_data[15]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(n9[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i16.GSR = "DISABLED";
    FD1P3AX instr_data_3__i15 (.D(instr_data[14]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(n9[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i15.GSR = "DISABLED";
    FD1P3AX instr_data_3__i14 (.D(instr_data[13]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(n9[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i14.GSR = "DISABLED";
    PFUMX i22390 (.BLUT(n24929), .ALUT(\mem_data_from_read[6] ), .C0(counter_hi[2]), 
          .Z(n24930));
    FD1P3AX instr_data_3__i13 (.D(instr_data[12]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(n9[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i13.GSR = "DISABLED";
    FD1P3AX instr_data_3__i12 (.D(instr_data[11]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(n9[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i12.GSR = "DISABLED";
    PFUMX mux_1013_i4 (.BLUT(n1629[3]), .ALUT(n1649[3]), .C0(n25338), 
          .Z(instr[19]));
    FD1P3AX instr_data_3__i11 (.D(instr_data[10]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(n9[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i11.GSR = "DISABLED";
    FD1P3AX instr_data_3__i10 (.D(instr_data[9]), .SP(clk_c_enable_91), 
            .CK(clk_c), .Q(n9[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i10.GSR = "DISABLED";
    FD1P3AX instr_len_i2 (.D(instr_len_2__N_307[1]), .SP(clk_c_enable_84), 
            .CK(clk_c), .Q(\instr_len[2] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_len_i2.GSR = "DISABLED";
    FD1P3AX instr_data_3__i9 (.D(instr_data[8]), .SP(clk_c_enable_91), .CK(clk_c), 
            .Q(n9[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i9.GSR = "DISABLED";
    FD1P3AX instr_data_3__i8 (.D(instr_data[7]), .SP(clk_c_enable_91), .CK(clk_c), 
            .Q(n9[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i8.GSR = "DISABLED";
    FD1P3AX instr_data_3__i7 (.D(instr_data[6]), .SP(clk_c_enable_91), .CK(clk_c), 
            .Q(n9[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i7.GSR = "DISABLED";
    FD1P3AX instr_data_3__i6 (.D(instr_data[5]), .SP(clk_c_enable_91), .CK(clk_c), 
            .Q(n9[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i6.GSR = "DISABLED";
    FD1P3AX instr_data_3__i5 (.D(instr_data[4]), .SP(clk_c_enable_91), .CK(clk_c), 
            .Q(n9[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i5.GSR = "DISABLED";
    FD1P3AX instr_data_3__i4 (.D(instr_data[3]), .SP(clk_c_enable_91), .CK(clk_c), 
            .Q(n9[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i4.GSR = "DISABLED";
    FD1P3AX instr_data_3__i3 (.D(instr_data[2]), .SP(clk_c_enable_91), .CK(clk_c), 
            .Q(n9[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i3.GSR = "DISABLED";
    FD1P3IX was_early_branch_424 (.D(was_early_branch_N_759), .SP(clk_c_enable_197), 
            .CD(n25424), .CK(clk_c), .Q(was_early_branch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(315[12] 320[8])
    defparam was_early_branch_424.GSR = "DISABLED";
    FD1P3AX instr_data_3__i2 (.D(instr_data_0__15__N_369[49]), .SP(clk_c_enable_93), 
            .CK(clk_c), .Q(n9[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i2.GSR = "DISABLED";
    FD1P3IX is_branch_399 (.D(is_branch_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_branch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_branch_399.GSR = "DISABLED";
    FD1P3AX rd_i0_i3 (.D(n3675[3]), .SP(clk_c_enable_312), .CK(clk_c), 
            .Q(rd[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i3.GSR = "DISABLED";
    FD1P3AX rd_i0_i2 (.D(n3675[2]), .SP(clk_c_enable_312), .CK(clk_c), 
            .Q(rd[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i2.GSR = "DISABLED";
    FD1P3AX rd_i0_i1 (.D(n3675[1]), .SP(clk_c_enable_312), .CK(clk_c), 
            .Q(rd[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i1.GSR = "DISABLED";
    FD1P3AX instr_fetch_running_429 (.D(n5438), .SP(clk_c_enable_102), .CK(clk_c), 
            .Q(instr_fetch_running)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_fetch_running_429.GSR = "DISABLED";
    FD1P3IX pc_offset__i14 (.D(pc_23__N_642[11]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[14] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i14.GSR = "DISABLED";
    FD1P3IX interrupt_core_408 (.D(n25179), .SP(clk_c_enable_110), .CD(n25424), 
            .CK(clk_c), .Q(interrupt_core)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam interrupt_core_408.GSR = "DISABLED";
    FD1S3IX data_ready_sync_415 (.D(data_ready_core), .CK(clk_c), .CD(n25424), 
            .Q(data_ready_sync)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(235[12] 256[8])
    defparam data_ready_sync_415.GSR = "DISABLED";
    FD1P3IX is_alu_imm_394 (.D(is_alu_imm_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_alu_imm)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_alu_imm_394.GSR = "DISABLED";
    PFUMX i22379 (.BLUT(n24915), .ALUT(n24914), .C0(n25284), .Z(n24916));
    FD1P3IX pc_offset__i1 (.D(pc_2__N_663[0]), .SP(clk_c_enable_393), .CD(n25424), 
            .CK(clk_c), .Q(\pc[1] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i1.GSR = "DISABLED";
    FD1P3IX data_addr__i0 (.D(addr_out[0]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i0.GSR = "DISABLED";
    FD1P3AX rs2_i0_i0 (.D(n1729[0]), .SP(clk_c_enable_312), .CK(clk_c), 
            .Q(rs2[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i0.GSR = "DISABLED";
    FD1P3AX instr_data_3__i64 (.D(instr_data[15]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i64.GSR = "DISABLED";
    FD1P3IX pc_offset__i2 (.D(pc_2__N_663[1]), .SP(clk_c_enable_393), .CD(n25424), 
            .CK(clk_c), .Q(\pc[2] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i2.GSR = "DISABLED";
    FD1P3IX pc_offset__i3 (.D(pc_23__N_642[0]), .SP(clk_c_enable_393), .CD(n25424), 
            .CK(clk_c), .Q(\pc[3] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i3.GSR = "DISABLED";
    FD1P3IX pc_offset__i4 (.D(pc_23__N_642[1]), .SP(clk_c_enable_393), .CD(n25424), 
            .CK(clk_c), .Q(\pc[4] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i4.GSR = "DISABLED";
    FD1P3AX instr_data_3__i63 (.D(instr_data[14]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i63.GSR = "DISABLED";
    FD1P3AX instr_data_3__i62 (.D(instr_data[13]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i62.GSR = "DISABLED";
    FD1P3AX instr_data_3__i61 (.D(instr_data[12]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i61.GSR = "DISABLED";
    FD1P3AX instr_data_3__i60 (.D(instr_data[11]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i60.GSR = "DISABLED";
    FD1P3AX instr_data_3__i59 (.D(instr_data[10]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i59.GSR = "DISABLED";
    FD1P3AX instr_data_3__i58 (.D(instr_data[9]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i58.GSR = "DISABLED";
    FD1P3AX instr_data_3__i57 (.D(instr_data[8]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i57.GSR = "DISABLED";
    FD1P3IX is_auipc_395 (.D(is_auipc_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_auipc)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_auipc_395.GSR = "DISABLED";
    FD1S3IX counter_hi_3136__i2 (.D(n25407), .CK(clk_c), .CD(n25424), 
            .Q(counter_hi[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3136__i2.GSR = "DISABLED";
    FD1P3IX pc_offset__i5 (.D(pc_23__N_642[2]), .SP(clk_c_enable_393), .CD(n25424), 
            .CK(clk_c), .Q(\pc[5] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i5.GSR = "DISABLED";
    FD1P3IX pc_offset__i6 (.D(pc_23__N_642[3]), .SP(clk_c_enable_393), .CD(n25424), 
            .CK(clk_c), .Q(\pc[6] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i6.GSR = "DISABLED";
    FD1P3IX pc_offset__i7 (.D(pc_23__N_642[4]), .SP(clk_c_enable_393), .CD(n25424), 
            .CK(clk_c), .Q(\pc[7] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i7.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i2 (.D(additional_mem_ops_2__N_480[2]), .CK(clk_c), 
            .CD(n25424), .Q(additional_mem_ops[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i2.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i1 (.D(additional_mem_ops_2__N_480[1]), .CK(clk_c), 
            .CD(n25424), .Q(additional_mem_ops[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i1.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i3 (.D(\next_instr_write_offset[3] ), .CK(clk_c), 
            .CD(n20739), .Q(\instr_write_offset[3] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i3.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i2 (.D(instr_write_offset_3__N_665[1]), .CK(clk_c), 
            .CD(n25424), .Q(instr_addr_23__N_49[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i2.GSR = "DISABLED";
    FD1S3IX addr_offset_3137__i2 (.D(n17[0]), .CK(clk_c), .CD(n25424), 
            .Q(addr_offset[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam addr_offset_3137__i2.GSR = "DISABLED";
    PFUMX i22359 (.BLUT(n25207), .ALUT(n24876), .C0(n3615), .Z(n24877));
    LUT4 i3564_2_lut_rep_698 (.A(rd[1]), .B(rd[0]), .Z(n25434)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(180[19:31])
    defparam i3564_2_lut_rep_698.init = 16'h8888;
    FD1P3IX is_alu_reg_397 (.D(is_alu_reg_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_alu_reg)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_alu_reg_397.GSR = "DISABLED";
    LUT4 i3571_2_lut_3_lut (.A(rd[1]), .B(rd[0]), .C(rd[2]), .Z(n5599)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(180[19:31])
    defparam i3571_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_4_lut (.A(n25178), .B(rst_reg_n), .C(n27), .D(n25171), 
         .Z(n3989)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h4000;
    LUT4 i3_4_lut_rep_431_4_lut (.A(n25178), .B(n25175), .C(n21916), .D(n25190), 
         .Z(n25167)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_4_lut_rep_431_4_lut.init = 16'h4000;
    LUT4 i1274_2_lut_3_lut_4_lut_4_lut (.A(\instr_len[2] ), .B(\pc[2] ), 
         .C(\pc[1] ), .D(instr_len[1]), .Z(n2015)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (B+(C (D)+!C !(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1274_2_lut_3_lut_4_lut_4_lut.init = 16'h0990;
    LUT4 i1269_2_lut_3_lut_4_lut_4_lut (.A(\instr_len[2] ), .B(\pc[2] ), 
         .C(\pc[1] ), .D(instr_len[1]), .Z(n2010)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A ((C (D)+!C !(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1269_2_lut_3_lut_4_lut_4_lut.init = 16'h0660;
    LUT4 n4956_bdd_3_lut_22427 (.A(\data_from_read[2] ), .B(n8229), .C(\gpio_out_sel[7] ), 
         .Z(n24997)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam n4956_bdd_3_lut_22427.init = 16'heaea;
    LUT4 mux_1003_i13_3_lut (.A(n2[12]), .B(n7[12]), .C(n1949), .Z(n1629[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1007_i14_3_lut (.A(n9[13]), .B(n14[13]), .C(n1969), .Z(n1649[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i14_3_lut.init = 16'hcaca;
    LUT4 instr_1__bdd_4_lut (.A(n26598), .B(n25284), .C(n25279), .D(n26597), 
         .Z(n25005)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !((C)+!B)) */ ;
    defparam instr_1__bdd_4_lut.init = 16'h8c8e;
    LUT4 mux_1003_i14_3_lut (.A(n2[13]), .B(n7[13]), .C(n1949), .Z(n1629[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1266_i5_3_lut_then_3_lut (.A(n9[4]), .B(n7[4]), .C(n1969), 
         .Z(n25451)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i5_3_lut_then_3_lut.init = 16'hacac;
    LUT4 mux_1266_i5_3_lut_else_3_lut (.A(n14[4]), .B(n2[4]), .C(n1949), 
         .Z(n25450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i5_3_lut_else_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_319 (.A(n25178), .B(n26612), .C(n25164), .D(n10_c), 
         .Z(n21067)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_319.init = 16'h4000;
    LUT4 i16_4_lut (.A(n3619), .B(clk_c_enable_38), .C(rst_reg_n), .D(n21297), 
         .Z(clk_c_enable_368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i16_4_lut.init = 16'hcfca;
    LUT4 i1_4_lut (.A(n21750), .B(n25178), .C(n7955), .D(instr_complete_N_1378), 
         .Z(n8)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut.init = 16'hfefc;
    LUT4 i1_4_lut_then_4_lut (.A(instr_len[1]), .B(\pc[1] ), .C(instr_addr_23__N_49[1]), 
         .D(instr_addr_23__N_49[0]), .Z(n25457)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_4_lut_then_4_lut.init = 16'h781e;
    LUT4 i1_4_lut_else_4_lut (.A(instr_len[1]), .B(\pc[1] ), .C(instr_addr_23__N_49[1]), 
         .D(instr_addr_23__N_49[0]), .Z(n25456)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_4_lut_else_4_lut.init = 16'h87e1;
    LUT4 i1_4_lut_adj_320 (.A(n26), .B(n22286), .C(n35), .D(n22), .Z(n22298)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_320.init = 16'hccc8;
    LUT4 mux_1568_i2_3_lut (.A(n2937[1]), .B(n24568), .C(n3619), .Z(n2978[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1568_i2_3_lut.init = 16'hcaca;
    LUT4 i21940_3_lut (.A(n3615), .B(n25166), .C(n25338), .Z(n23265)) /* synthesis lut_function=(A+!((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21940_3_lut.init = 16'haeae;
    LUT4 i1_4_lut_4_lut_adj_321 (.A(n25178), .B(n21978), .C(n16), .D(n25171), 
         .Z(n1943)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_321.init = 16'h4000;
    LUT4 mux_1266_i13_3_lut_then_3_lut (.A(n9[12]), .B(n7[12]), .C(n1969), 
         .Z(n25468)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i13_3_lut_then_3_lut.init = 16'hacac;
    LUT4 mux_1266_i13_3_lut_else_3_lut (.A(n14[12]), .B(n2[12]), .C(n1949), 
         .Z(n25467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i13_3_lut_else_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_322 (.A(n25178), .B(n22050), .C(n6), .D(n25171), 
         .Z(n22056)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_322.init = 16'h4000;
    LUT4 i1_4_lut_adj_323 (.A(next_pc_offset[3]), .B(n6830), .C(\instr_write_offset[3] ), 
         .D(n5879), .Z(n21541)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C)+!B (C (D)+!C !(D)))) */ ;
    defparam i1_4_lut_adj_323.init = 16'ha596;
    LUT4 n15_bdd_4_lut (.A(n26598), .B(n25284), .C(n25221), .D(n26597), 
         .Z(n25015)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;
    defparam n15_bdd_4_lut.init = 16'hc800;
    LUT4 i1_4_lut_adj_324 (.A(\instr_write_offset[3] ), .B(instr_addr_23__N_49[1]), 
         .C(n5856), .D(n21390), .Z(n8146)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_324.init = 16'h565a;
    LUT4 mux_1568_i4_3_lut (.A(n2937[3]), .B(n2890[3]), .C(n3619), .Z(n2978[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1568_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1568_i6_3_lut (.A(n2937[5]), .B(n2890[5]), .C(n3619), .Z(n2978[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1568_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1568_i7_3_lut (.A(n2937[6]), .B(n2890[6]), .C(n3619), .Z(n2978[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1568_i7_3_lut.init = 16'hcaca;
    LUT4 mem_data_ready_bdd_3_lut_22487 (.A(\qspi_data_buf[25] ), .B(\qspi_data_buf[29] ), 
         .C(counter_hi[2]), .Z(n25028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mem_data_ready_bdd_3_lut_22487.init = 16'hcaca;
    LUT4 i11740_2_lut_rep_428_3_lut_4_lut (.A(n25177), .B(n25182), .C(n25178), 
         .D(n22126), .Z(n25164)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i11740_2_lut_rep_428_3_lut_4_lut.init = 16'hf0fe;
    LUT4 mux_1540_i10_3_lut_4_lut (.A(n3613), .B(n3605), .C(n2703[9]), 
         .D(n2414[9]), .Z(n2854[9])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1540_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i21947_2_lut_3_lut_4_lut (.A(n3613), .B(n3605), .C(n3619), .D(n25155), 
         .Z(n23237)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21947_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 mux_2749_i25_3_lut (.A(instr[31]), .B(instr[24]), .C(n25209), 
         .Z(n4516[24])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2749_i25_3_lut.init = 16'hacac;
    LUT4 i3976_2_lut_rep_575_4_lut (.A(qspi_data_ready), .B(n25361), .C(instr_fetch_running), 
         .D(instr_addr_23__N_49[0]), .Z(n25311)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[64:98])
    defparam i3976_2_lut_rep_575_4_lut.init = 16'h8000;
    LUT4 mux_2749_i26_3_lut (.A(instr[31]), .B(instr[25]), .C(n25209), 
         .Z(n4516[25])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2749_i26_3_lut.init = 16'hacac;
    LUT4 mem_data_ready_bdd_3_lut_22452 (.A(counter_hi[2]), .B(instr_data[9]), 
         .C(instr_data[13]), .Z(n25027)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mem_data_ready_bdd_3_lut_22452.init = 16'he4e4;
    LUT4 i1_2_lut_4_lut (.A(qspi_data_ready), .B(n25361), .C(instr_fetch_running), 
         .D(n25415), .Z(n21962)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[64:98])
    defparam i1_2_lut_4_lut.init = 16'hff7f;
    LUT4 i1_2_lut_4_lut_adj_325 (.A(qspi_data_ready), .B(n25361), .C(instr_fetch_running), 
         .D(n25406), .Z(n21884)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[64:98])
    defparam i1_2_lut_4_lut_adj_325.init = 16'h8000;
    LUT4 i409_2_lut_rep_429_3_lut_4_lut (.A(n25177), .B(n25182), .C(n25178), 
         .D(n22126), .Z(clk_c_enable_38)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i409_2_lut_rep_429_3_lut_4_lut.init = 16'h000e;
    LUT4 mux_2749_i28_3_lut (.A(instr[31]), .B(instr[27]), .C(n25209), 
         .Z(n4516[27])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2749_i28_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_4_lut_adj_326 (.A(qspi_data_ready), .B(n25361), .C(instr_fetch_running), 
         .D(n25409), .Z(n21970)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[64:98])
    defparam i1_2_lut_4_lut_adj_326.init = 16'hff7f;
    LUT4 mem_data_from_read_17__bdd_3_lut_22491 (.A(\mem_data_from_read[17] ), 
         .B(counter_hi[2]), .C(\mem_data_from_read[21] ), .Z(n25030)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam mem_data_from_read_17__bdd_3_lut_22491.init = 16'he2e2;
    LUT4 n25030_bdd_3_lut (.A(n25030), .B(n25029), .C(counter_hi[3]), 
         .Z(n25031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25030_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_327 (.A(qspi_data_ready), .B(n25361), .C(instr_fetch_running), 
         .D(n25394), .Z(n21966)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[64:98])
    defparam i1_2_lut_4_lut_adj_327.init = 16'hff7f;
    LUT4 mux_1256_i9_3_lut (.A(n14[8]), .B(n2[8]), .C(n1949), .Z(n1950[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i9_3_lut.init = 16'hcaca;
    LUT4 i21923_3_lut_4_lut (.A(n25370), .B(counter_hi[3]), .C(is_timer_addr), 
         .D(data_out_3__N_1116), .Z(n23106)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam i21923_3_lut_4_lut.init = 16'hff04;
    LUT4 mux_2749_i29_3_lut (.A(instr[31]), .B(instr[28]), .C(n25209), 
         .Z(n4516[28])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2749_i29_3_lut.init = 16'hacac;
    LUT4 shift_right_317_i271_3_lut (.A(n23062), .B(load_top_bit), .C(data_out_3__N_1116), 
         .Z(debug_branch_N_571[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam shift_right_317_i271_3_lut.init = 16'hcaca;
    LUT4 mux_2749_i30_3_lut (.A(instr[31]), .B(instr[29]), .C(n25209), 
         .Z(n4516[29])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2749_i30_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n25177), .B(n25182), .C(n21369), .D(n22126), 
         .Z(clk_c_enable_203)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 i1_4_lut_adj_328 (.A(clk_c_enable_312), .B(n25178), .C(n22272), 
         .D(n25175), .Z(n3993)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_328.init = 16'ha888;
    LUT4 shift_right_317_i269_3_lut (.A(n23059), .B(load_top_bit), .C(data_out_3__N_1116), 
         .Z(debug_branch_N_571[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam shift_right_317_i269_3_lut.init = 16'hcaca;
    LUT4 mux_1260_i9_3_lut (.A(n7[8]), .B(n9[8]), .C(n1969), .Z(n1970[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i9_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_433_4_lut (.A(n25177), .B(n25182), .C(n22126), .D(n25178), 
         .Z(n25169)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i1_3_lut_rep_433_4_lut.init = 16'hfff1;
    PFUMX i22523 (.BLUT(n25438), .ALUT(n25439), .C0(counter_hi[2]), .Z(n25440));
    FD1P3IX is_jalr_400 (.D(is_jalr_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_jalr)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_jalr_400.GSR = "DISABLED";
    LUT4 mux_1003_i1_rep_117_3_lut (.A(n2[0]), .B(n7[0]), .C(n1949), .Z(n22996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i1_rep_117_3_lut.init = 16'hcaca;
    FD1P3AX data_continue_420 (.D(data_continue_N_694), .SP(clk_c_enable_194), 
            .CK(clk_c), .Q(debug_data_continue)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_continue_420.GSR = "DISABLED";
    FD1P3IX is_jal_401 (.D(is_jal_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_jal)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_jal_401.GSR = "DISABLED";
    LUT4 mux_1256_i8_3_lut (.A(n14[7]), .B(n2[7]), .C(n1949), .Z(n1950[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1013_i1_rep_111_3_lut (.A(n1649[0]), .B(instr[31]), .C(n3597), 
         .Z(n22990)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i1_rep_111_3_lut.init = 16'hcaca;
    FD1P3IX data_out__i0 (.D(data_out_slice[0]), .SP(clk_c_enable_324), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i0.GSR = "DISABLED";
    LUT4 mux_1260_i8_3_lut (.A(n7[7]), .B(n9[7]), .C(n1969), .Z(n1970[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i8_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(n25372), .B(rst_reg_n), .C(data_ready_latch), 
         .D(clk_c_enable_54), .Z(clk_c_enable_15)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_3_lut_4_lut.init = 16'hff7f;
    FD1P3JX no_write_in_progress_419 (.D(no_write_in_progress_N_202), .SP(clk_c_enable_197), 
            .PD(n25424), .CK(clk_c), .Q(no_write_in_progress)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam no_write_in_progress_419.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_329 (.A(n25372), .B(rst_reg_n), .C(data_ready_latch), 
         .D(n20805), .Z(n21632)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_329.init = 16'h0008;
    LUT4 mux_1007_i1_3_lut (.A(n9[0]), .B(n14[0]), .C(n1969), .Z(n1649[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i1_3_lut.init = 16'hcaca;
    FD1P3IX pc_offset__i15 (.D(pc_23__N_642[12]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[15] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i15.GSR = "DISABLED";
    FD1P3AX data_write_n_i0 (.D(data_write_n_1__N_100[0]), .SP(clk_c_enable_314), 
            .CK(clk_c), .Q(qv_data_write_n[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_write_n_i0.GSR = "DISABLED";
    LUT4 mux_1013_i1_3_lut (.A(n22996), .B(n1649[0]), .C(n25338), .Z(instr[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i1_3_lut.init = 16'hcaca;
    LUT4 i21658_3_lut_4_lut_4_lut (.A(n25156), .B(n21236), .C(n3611), 
         .D(n25290), .Z(n2813[7])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i21658_3_lut_4_lut_4_lut.init = 16'hc5c0;
    FD1P3IX pc_offset__i16 (.D(pc_23__N_642[13]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[16] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i16.GSR = "DISABLED";
    FD1P3IX is_system_402 (.D(is_system_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_system)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_system_402.GSR = "DISABLED";
    FD1P3IX is_lui_398 (.D(is_lui_de), .SP(clk_c_enable_203), .CD(n25424), 
            .CK(clk_c), .Q(is_lui)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_lui_398.GSR = "DISABLED";
    LUT4 mux_1003_i15_3_lut (.A(n2[14]), .B(n7[14]), .C(n1949), .Z(n1629[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i15_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_440 (.A(clk_c_enable_54), .B(n25181), .C(is_load), 
         .Z(n25176)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_440.init = 16'h2020;
    LUT4 i1_2_lut_4_lut_adj_330 (.A(clk_c_enable_54), .B(n25181), .C(is_load), 
         .D(n20762), .Z(clk_c_enable_194)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;
    defparam i1_2_lut_4_lut_adj_330.init = 16'hff20;
    LUT4 i1_3_lut_4_lut_adj_331 (.A(n21402), .B(n25181), .C(n22028), .D(n8), 
         .Z(n21322)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[22:78])
    defparam i1_3_lut_4_lut_adj_331.init = 16'h00d0;
    LUT4 i43_3_lut (.A(n25281), .B(n25279), .C(n20641), .Z(n24)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;
    defparam i43_3_lut.init = 16'h6464;
    LUT4 i1_2_lut_rep_435_3_lut_4_lut (.A(n21402), .B(n25181), .C(n22126), 
         .D(n25182), .Z(n25171)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[22:78])
    defparam i1_2_lut_rep_435_3_lut_4_lut.init = 16'h0f0d;
    LUT4 i21469_3_lut (.A(\mem_data_from_read[27] ), .B(\mem_data_from_read[31] ), 
         .C(counter_hi[2]), .Z(n23065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam i21469_3_lut.init = 16'hcaca;
    LUT4 next_pc_for_core_23__I_0_i271_4_lut (.A(n5047[2]), .B(debug_rd_3__N_136[30]), 
         .C(n25381), .D(n6657), .Z(debug_branch_N_177[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i271_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut_3_lut (.A(any_additional_mem_ops), .B(n25180), .C(n4030[0]), 
         .Z(additional_mem_ops_2__N_480[0])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i1_2_lut_3_lut.init = 16'h7878;
    LUT4 i1_3_lut_4_lut_adj_332 (.A(any_additional_mem_ops), .B(n25180), 
         .C(n4030[0]), .D(n4030[1]), .Z(additional_mem_ops_2__N_480[1])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i1_3_lut_4_lut_adj_332.init = 16'hf708;
    LUT4 gnd_bdd_2_lut_22140_2_lut_3_lut (.A(any_additional_mem_ops), .B(n25180), 
         .C(n24486), .Z(n24487)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam gnd_bdd_2_lut_22140_2_lut_3_lut.init = 16'h7070;
    LUT4 n24419_bdd_3_lut (.A(n24419), .B(instr[31]), .C(n25209), .Z(n24420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24419_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_1256_i10_3_lut (.A(n14[9]), .B(n2[9]), .C(n1949), .Z(n1950[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i10_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_333 (.A(n25237), .B(n25279), .C(n25244), .D(n26612), 
         .Z(n21944)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_333.init = 16'h4000;
    LUT4 mux_1260_i10_3_lut (.A(n7[9]), .B(n9[9]), .C(n1969), .Z(n1970[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i10_3_lut.init = 16'hcaca;
    LUT4 i21477_3_lut (.A(n23060), .B(timer_data[0]), .C(is_timer_addr), 
         .Z(n8755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam i21477_3_lut.init = 16'hcaca;
    FD1P3IX pc_offset__i17 (.D(pc_23__N_642[14]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[17] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i17.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_334 (.A(n22_adj_2374), .B(n7955), .C(n4), .D(n25196), 
         .Z(n22324)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_334.init = 16'h0200;
    LUT4 mux_1013_i3_3_lut (.A(n22992), .B(n1649[2]), .C(n25338), .Z(instr[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i3_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_335 (.A(n20952), .B(instr_fetch_running_N_676), .C(instr_fetch_restart_N_678), 
         .D(debug_stall_txn), .Z(n21800)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(435[34:115])
    defparam i1_4_lut_adj_335.init = 16'h5010;
    LUT4 mux_1256_i11_3_lut (.A(n14[10]), .B(n2[10]), .C(n1949), .Z(n1950[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i11_3_lut.init = 16'hcaca;
    LUT4 n2733_bdd_4_lut_22506 (.A(n2703[2]), .B(n3613), .C(n26598), .D(instr[4]), 
         .Z(n25118)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B (C (D)))) */ ;
    defparam n2733_bdd_4_lut_22506.init = 16'he222;
    LUT4 mux_1260_i11_3_lut (.A(n7[10]), .B(n9[10]), .C(n1969), .Z(n1970[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i11_3_lut.init = 16'hcaca;
    LUT4 n2733_bdd_4_lut (.A(n25153), .B(n3611), .C(n21121), .D(n25266), 
         .Z(n25119)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (C))) */ ;
    defparam n2733_bdd_4_lut.init = 16'he2c0;
    LUT4 i21481_3_lut (.A(n23063), .B(timer_data[2]), .C(is_timer_addr), 
         .Z(n8759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam i21481_3_lut.init = 16'hcaca;
    LUT4 mux_2750_i9_3_lut (.A(n25284), .B(instr[31]), .C(n3597), .Z(n4548[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2750_i9_3_lut.init = 16'hcaca;
    LUT4 mux_2750_i8_3_lut (.A(n26598), .B(instr[31]), .C(n3597), .Z(n4548[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2750_i8_3_lut.init = 16'hcaca;
    LUT4 mux_2750_i7_3_lut (.A(n25279), .B(instr[31]), .C(n3597), .Z(n4548[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2750_i7_3_lut.init = 16'hcaca;
    LUT4 mux_2750_i6_3_lut (.A(instr[12]), .B(instr[31]), .C(n3597), .Z(n4548[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2750_i6_3_lut.init = 16'hcaca;
    LUT4 n24421_bdd_3_lut (.A(n24419), .B(instr[31]), .C(n3597), .Z(n24422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24421_bdd_3_lut.init = 16'hcaca;
    LUT4 n1664_bdd_3_lut (.A(n1649[1]), .B(n25338), .C(n22994), .Z(n24419)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n1664_bdd_3_lut.init = 16'hb8b8;
    LUT4 i1_4_lut_adj_336 (.A(clk_c_enable_312), .B(n25178), .C(n22092), 
         .D(n25175), .Z(n3991)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_336.init = 16'ha888;
    LUT4 next_pc_for_core_23__I_0_i270_4_lut (.A(n5047[1]), .B(debug_rd_3__N_136[29]), 
         .C(n25381), .D(n6657), .Z(debug_branch_N_177[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i270_4_lut.init = 16'hcac0;
    LUT4 next_pc_for_core_23__I_0_i272_4_lut (.A(n5047[3]), .B(debug_rd_3__N_136[31]), 
         .C(n25381), .D(n6657), .Z(debug_branch_N_177[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i272_4_lut.init = 16'hcac0;
    LUT4 i20798_3_lut (.A(\next_pc_for_core[3] ), .B(\next_pc_for_core[7] ), 
         .C(counter_hi[2]), .Z(n23073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20798_3_lut.init = 16'hcaca;
    FD1P3IX pc_offset__i18 (.D(pc_23__N_642[15]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[18] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i18.GSR = "DISABLED";
    LUT4 i21169_3_lut (.A(imm[27]), .B(imm[31]), .C(counter_hi[2]), .Z(n23444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21169_3_lut.init = 16'hcaca;
    LUT4 i21168_3_lut (.A(\imm[19] ), .B(\imm[23] ), .C(counter_hi[2]), 
         .Z(n23443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21168_3_lut.init = 16'hcaca;
    LUT4 mux_1013_i5_3_lut (.A(n22959), .B(n22970), .C(n25338), .Z(instr[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i5_3_lut.init = 16'hcaca;
    LUT4 n2952_bdd_3_lut_22104 (.A(n2937[17]), .B(n24424), .C(n3619), 
         .Z(n24425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n2952_bdd_3_lut_22104.init = 16'hcaca;
    LUT4 i1_2_lut (.A(qv_data_read_n[0]), .B(qv_data_read_n[1]), .Z(n17512)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 n24426_bdd_3_lut (.A(n24428), .B(instr[31]), .C(n25209), .Z(n24427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24426_bdd_3_lut.init = 16'hcaca;
    LUT4 i21167_3_lut (.A(\imm[11] ), .B(\imm[15] ), .C(counter_hi[2]), 
         .Z(n23442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21167_3_lut.init = 16'hcaca;
    LUT4 i21166_3_lut (.A(\imm[3] ), .B(\imm[7] ), .C(counter_hi[2]), 
         .Z(n23441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21166_3_lut.init = 16'hcaca;
    LUT4 n3597_bdd_3_lut_22175 (.A(n1649[2]), .B(n25338), .C(n22992), 
         .Z(n24428)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n3597_bdd_3_lut_22175.init = 16'hb8b8;
    LUT4 mux_1568_i25_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n4516[24]), .Z(n2978[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1568_i25_3_lut_4_lut.init = 16'hf870;
    LUT4 n24428_bdd_3_lut (.A(n24428), .B(instr[31]), .C(n3597), .Z(n24429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24428_bdd_3_lut.init = 16'hcaca;
    LUT4 i21162_3_lut (.A(imm[26]), .B(imm[30]), .C(counter_hi[2]), .Z(n23437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21162_3_lut.init = 16'hcaca;
    LUT4 i21161_3_lut (.A(\imm[18] ), .B(\imm[22] ), .C(counter_hi[2]), 
         .Z(n23436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21161_3_lut.init = 16'hcaca;
    LUT4 i4615_3_lut_4_lut (.A(instr_addr_23__N_49[0]), .B(n25420), .C(n25363), 
         .D(instr_addr_23__N_49[1]), .Z(n6830)) /* synthesis lut_function=(A (D)+!A !(B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i4615_3_lut_4_lut.init = 16'hbf00;
    LUT4 i21160_3_lut (.A(\imm[10] ), .B(\imm[14] ), .C(counter_hi[2]), 
         .Z(n23435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21160_3_lut.init = 16'hcaca;
    LUT4 i21159_3_lut (.A(\imm[2] ), .B(\imm[6] ), .C(counter_hi[2]), 
         .Z(n23434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21159_3_lut.init = 16'hcaca;
    LUT4 i21155_3_lut (.A(imm[25]), .B(imm[29]), .C(counter_hi[2]), .Z(n23430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21155_3_lut.init = 16'hcaca;
    LUT4 i21154_3_lut (.A(\imm[17] ), .B(\imm[21] ), .C(counter_hi[2]), 
         .Z(n23429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21154_3_lut.init = 16'hcaca;
    LUT4 i11754_3_lut (.A(any_additional_mem_ops), .B(rst_reg_n), .C(n25176), 
         .Z(data_continue_N_694)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i11754_3_lut.init = 16'ha8a8;
    LUT4 mux_1568_i26_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n4516[25]), .Z(n2978[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1568_i26_3_lut_4_lut.init = 16'hf870;
    LUT4 i29_4_lut (.A(n26596), .B(n25248), .C(n25203), .D(n25278), 
         .Z(n16)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)+!B !(C+(D))))) */ ;
    defparam i29_4_lut.init = 16'h3534;
    LUT4 mux_1568_i30_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n4516[29]), .Z(n2978[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1568_i30_3_lut_4_lut.init = 16'hf870;
    LUT4 n2952_bdd_3_lut_22120 (.A(n2937[17]), .B(n24431), .C(n3619), 
         .Z(n24432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n2952_bdd_3_lut_22120.init = 16'hcaca;
    LUT4 mux_1568_i28_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n4516[27]), .Z(n2978[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1568_i28_3_lut_4_lut.init = 16'hf870;
    LUT4 n25283_bdd_4_lut_22958 (.A(n25210), .B(n25284), .C(n25279), .D(n26598), 
         .Z(n26286)) /* synthesis lut_function=(!(A (B (D)+!B !((D)+!C))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam n25283_bdd_4_lut_22958.init = 16'h33cb;
    LUT4 i21153_3_lut (.A(\imm[9] ), .B(\imm[13] ), .C(counter_hi[2]), 
         .Z(n23428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21153_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_337 (.A(clk_c_enable_312), .B(n25178), .C(n22282), 
         .D(n25175), .Z(n1945)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_337.init = 16'ha888;
    LUT4 i21152_3_lut (.A(\imm[1] ), .B(\imm[5] ), .C(counter_hi[2]), 
         .Z(n23427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21152_3_lut.init = 16'hcaca;
    FD1P3AX mem_op_increment_reg_413 (.D(n23084), .SP(clk_c_enable_209), 
            .CK(clk_c), .Q(mem_op_increment_reg)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_increment_reg_413.GSR = "DISABLED";
    LUT4 stall_core_I_0_438_2_lut_rep_590_4_lut (.A(debug_instr_valid), .B(n25383), 
         .C(no_write_in_progress), .D(interrupt_core), .Z(n25326)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(148[23:87])
    defparam stall_core_I_0_438_2_lut_rep_590_4_lut.init = 16'h005d;
    LUT4 n25283_bdd_4_lut_23028 (.A(n25284), .B(n1950[0]), .C(n1970[0]), 
         .D(n25338), .Z(n26288)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam n25283_bdd_4_lut_23028.init = 16'h5044;
    LUT4 i21148_3_lut (.A(imm[24]), .B(imm[28]), .C(counter_hi[2]), .Z(n23423)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21148_3_lut.init = 16'hcaca;
    LUT4 mux_1568_i29_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n4516[28]), .Z(n2978[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1568_i29_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_1013_i11_3_lut (.A(n22978), .B(n1649[10]), .C(n25338), .Z(instr[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i11_3_lut.init = 16'hcaca;
    LUT4 i21147_3_lut (.A(\imm[16] ), .B(\imm[20] ), .C(counter_hi[2]), 
         .Z(n23422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21147_3_lut.init = 16'hcaca;
    FD1P3AX instr_data_3__i56 (.D(instr_data[7]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i56.GSR = "DISABLED";
    FD1P3AX instr_data_3__i55 (.D(instr_data[6]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i55.GSR = "DISABLED";
    LUT4 i21146_3_lut (.A(\imm[8] ), .B(\imm[12] ), .C(counter_hi[2]), 
         .Z(n23421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21146_3_lut.init = 16'hcaca;
    FD1P3AX imm_i0_i0 (.D(n2978[0]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(imm[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i0.GSR = "DISABLED";
    LUT4 i21145_3_lut (.A(imm[0]), .B(\imm[4] ), .C(counter_hi[2]), .Z(n23420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21145_3_lut.init = 16'hcaca;
    FD1P3AX instr_data_3__i54 (.D(instr_data[5]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i54.GSR = "DISABLED";
    LUT4 mux_1544_i27_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n22978), .Z(n2890[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1544_i27_3_lut_4_lut.init = 16'hf870;
    FD1P3AX instr_data_3__i53 (.D(instr_data[4]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i53.GSR = "DISABLED";
    FD1P3AX instr_data_3__i52 (.D(instr_data[3]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i52.GSR = "DISABLED";
    FD1P3AX instr_data_3__i51 (.D(instr_data[2]), .SP(clk_c_enable_216), 
            .CK(clk_c), .Q(n14[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i51.GSR = "DISABLED";
    FD1P3AX instr_data_3__i50 (.D(instr_data_0__15__N_369[49]), .SP(clk_c_enable_218), 
            .CK(clk_c), .Q(n14[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i50.GSR = "DISABLED";
    FD1P3AX instr_data_3__i49 (.D(instr_data_0__15__N_369[0]), .SP(clk_c_enable_218), 
            .CK(clk_c), .Q(n14[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i49.GSR = "DISABLED";
    FD1P3AX instr_data_3__i48 (.D(instr_data[15]), .SP(clk_c_enable_219), 
            .CK(clk_c), .Q(n2[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i48.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_338 (.A(n25248), .B(n25249), .C(instr[23]), .D(n26612), 
         .Z(n22074)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_338.init = 16'h1000;
    LUT4 i21515_3_lut (.A(n23055), .B(n24999), .C(counter_hi[2]), .Z(n23057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam i21515_3_lut.init = 16'hcaca;
    LUT4 mux_1013_i8_3_lut (.A(n22966), .B(n22972), .C(n25338), .Z(instr[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i8_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_339 (.A(n25248), .B(n25249), .C(instr[22]), .D(n26612), 
         .Z(n22038)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_339.init = 16'h1000;
    LUT4 mux_1013_i7_3_lut (.A(n22964), .B(n22974), .C(n25338), .Z(instr[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i7_3_lut.init = 16'hcaca;
    LUT4 n3609_bdd_3_lut_22367 (.A(n3597), .B(instr[31]), .C(instr[19]), 
         .Z(n24450)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n3609_bdd_3_lut_22367.init = 16'hd8d8;
    L6MUX21 mux_1568_i1 (.D0(n2937[0]), .D1(n2890[0]), .SD(n3619), .Z(n2978[0]));
    LUT4 i1_4_lut_adj_340 (.A(n25248), .B(n25249), .C(instr[21]), .D(n26612), 
         .Z(n22062)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_340.init = 16'h1000;
    LUT4 mux_1013_i6_3_lut (.A(n22957), .B(n22968), .C(n25338), .Z(instr[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i6_3_lut.init = 16'hcaca;
    L6MUX21 mux_1568_i5 (.D0(n2937[4]), .D1(n2890[4]), .SD(n3619), .Z(n2978[4]));
    PFUMX mux_1559_i1 (.BLUT(n2813[0]), .ALUT(n22852), .C0(n25155), .Z(n2937[0]));
    LUT4 i11649_2_lut (.A(\next_pc_for_core[4] ), .B(counter_hi[2]), .Z(n149)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i11649_2_lut.init = 16'h8888;
    LUT4 n3609_bdd_3_lut_22116 (.A(n25209), .B(instr[31]), .C(instr[19]), 
         .Z(n24449)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n3609_bdd_3_lut_22116.init = 16'hd8d8;
    FD1P3IX pc_offset__i9 (.D(pc_23__N_642[6]), .SP(clk_c_enable_393), .CD(n25424), 
            .CK(clk_c), .Q(\pc[9] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i9.GSR = "DISABLED";
    PFUMX mux_1568_i21 (.BLUT(n22955), .ALUT(n2890[20]), .C0(n23155), 
          .Z(n2978[20]));
    LUT4 i1_4_lut_adj_341 (.A(n25248), .B(n25249), .C(instr[20]), .D(n26612), 
         .Z(n22050)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_341.init = 16'h1000;
    LUT4 debug_branch_I_23_i4_rep_65_3_lut (.A(timer_data[3]), .B(load_top_bit), 
         .C(data_out_3__N_1116), .Z(n22944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_23_i4_rep_65_3_lut.init = 16'hcaca;
    PFUMX mux_1568_i22 (.BLUT(n22953), .ALUT(n2890[21]), .C0(n23155), 
          .Z(n2978[21]));
    LUT4 i4449_4_lut_4_lut (.A(clk_c_enable_38), .B(n25226), .C(additional_mem_ops[0]), 
         .D(n25265), .Z(additional_mem_ops_de[0])) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i4449_4_lut_4_lut.init = 16'hd850;
    LUT4 n2952_bdd_3_lut_22122 (.A(n2937[17]), .B(n24452), .C(n3619), 
         .Z(n24453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n2952_bdd_3_lut_22122.init = 16'hcaca;
    LUT4 i20793_3_lut (.A(\next_pc_for_core[9] ), .B(\next_pc_for_core[13] ), 
         .C(counter_hi[2]), .Z(n23068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20793_3_lut.init = 16'hcaca;
    LUT4 mux_1544_i24_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n22966), .Z(n2890[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1544_i24_3_lut_4_lut.init = 16'hf870;
    LUT4 i5146_4_lut_4_lut (.A(clk_c_enable_38), .B(n25226), .C(additional_mem_ops[1]), 
         .D(n25264), .Z(additional_mem_ops_de[1])) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i5146_4_lut_4_lut.init = 16'hd850;
    LUT4 mux_1544_i23_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n22964), .Z(n2890[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1544_i23_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_1544_i22_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n22957), .Z(n2890[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1544_i22_3_lut_4_lut.init = 16'hf870;
    PFUMX mux_1568_i23 (.BLUT(n22961), .ALUT(n2890[22]), .C0(n23155), 
          .Z(n2978[22]));
    LUT4 n2952_bdd_3_lut (.A(n2937[17]), .B(n24877), .C(n3619), .Z(n24457)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n2952_bdd_3_lut.init = 16'hcaca;
    LUT4 i21130_3_lut (.A(n23403), .B(n25031), .C(counter_hi[4]), .Z(n23405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21130_3_lut.init = 16'hcaca;
    PFUMX mux_1568_i24 (.BLUT(n22963), .ALUT(n2890[23]), .C0(n23155), 
          .Z(n2978[23]));
    FD1P3IX pc_offset__i19 (.D(pc_23__N_642[16]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[19] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i19.GSR = "DISABLED";
    LUT4 instr_len_2__bdd_4_lut (.A(\instr_len[2] ), .B(\pc[1] ), .C(instr_len[1]), 
         .D(\pc[2] ), .Z(next_pc_offset[3])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B (C (D)))) */ ;
    defparam instr_len_2__bdd_4_lut.init = 16'hea80;
    LUT4 i18654_3_lut (.A(n10), .B(addr[27]), .C(addr[26]), .Z(n20805)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i18654_3_lut.init = 16'heaea;
    PFUMX mux_1568_i27 (.BLUT(n22977), .ALUT(n2890[26]), .C0(n23155), 
          .Z(n2978[26]));
    LUT4 next_pc_for_core_23__I_0_i269_4_lut (.A(n209), .B(n5047[0]), .C(n25359), 
         .D(n6657), .Z(debug_branch_N_177[28])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i269_4_lut.init = 16'haca0;
    L6MUX21 mux_1559_i6 (.D0(n2813[5]), .D1(n2854[5]), .SD(n25155), .Z(n2937[5]));
    LUT4 i1_2_lut_adj_342 (.A(addr[4]), .B(addr[5]), .Z(n22566)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_342.init = 16'h8888;
    PFUMX mux_1559_i5 (.BLUT(n2813[4]), .ALUT(n2854[4]), .C0(n25155), 
          .Z(n2937[4]));
    FD1P3IX pc_offset__i20 (.D(pc_23__N_642[17]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[20] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i20.GSR = "DISABLED";
    L6MUX21 mux_1568_i8 (.D0(n2937[7]), .D1(n2890[7]), .SD(n3619), .Z(n2978[7]));
    PFUMX mux_1568_i9 (.BLUT(n2854[8]), .ALUT(n2937[8]), .C0(n23245), 
          .Z(n2978[8]));
    LUT4 pc_23__I_0_450_i269_3_lut (.A(n209_adj_2376), .B(data_rs1[0]), 
         .C(n25402), .Z(debug_branch_N_173[28])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam pc_23__I_0_450_i269_3_lut.init = 16'hacac;
    PFUMX mux_1568_i10 (.BLUT(n2854[9]), .ALUT(n2937[9]), .C0(n23245), 
          .Z(n2978[9]));
    LUT4 pc_23__I_0_450_i157_rep_62_3_lut (.A(\pc[8] ), .B(\pc[12] ), .C(counter_hi[2]), 
         .Z(n22941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam pc_23__I_0_450_i157_rep_62_3_lut.init = 16'hcaca;
    LUT4 mux_1013_i7_rep_81_3_lut_3_lut (.A(n25166), .B(n25288), .C(n22974), 
         .Z(n22960)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1013_i7_rep_81_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_1013_i8_rep_83_3_lut_3_lut (.A(n25166), .B(n25287), .C(n22972), 
         .Z(n22962)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1013_i8_rep_83_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_1544_i21_3_lut_4_lut (.A(n3619), .B(n3615), .C(n4516[21]), 
         .D(n22959), .Z(n2890[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1544_i21_3_lut_4_lut.init = 16'hf870;
    LUT4 i11618_2_lut (.A(\pc[4] ), .B(counter_hi[2]), .Z(n149_adj_2377)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam i11618_2_lut.init = 16'h8888;
    LUT4 i21797_2_lut_rep_427 (.A(instr_fetch_running), .B(was_early_branch_N_759), 
         .Z(n25163)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21797_2_lut_rep_427.init = 16'h1111;
    PFUMX mux_1568_i11 (.BLUT(n2854[10]), .ALUT(n2937[10]), .C0(n23237), 
          .Z(n2978[10]));
    PFUMX i22243 (.BLUT(n24687), .ALUT(n24686), .C0(counter_hi[2]), .Z(n24688));
    PFUMX mux_1568_i12 (.BLUT(n2937[11]), .ALUT(n2890[11]), .C0(n3619), 
          .Z(n2978[11]));
    LUT4 i1_3_lut_rep_425_4_lut (.A(instr_fetch_running), .B(was_early_branch_N_759), 
         .C(instr_fetch_restart_N_678), .D(n20952), .Z(n25161)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_rep_425_4_lut.init = 16'h0010;
    LUT4 n21430_bdd_4_lut (.A(n21430), .B(n25458), .C(debug_instr_valid), 
         .D(\instr_avail_len[3] ), .Z(n25144)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n21430_bdd_4_lut.init = 16'hca00;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n25240), .B(n21067), .C(instr[4]), .D(n25263), 
         .Z(n21152)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut.init = 16'h0040;
    PFUMX mux_1568_i13 (.BLUT(n2937[12]), .ALUT(n2890[12]), .C0(n3619), 
          .Z(n2978[12]));
    PFUMX mux_1568_i14 (.BLUT(n2937[13]), .ALUT(n2890[13]), .C0(n3619), 
          .Z(n2978[13]));
    LUT4 i1_4_lut_4_lut_4_lut_adj_343 (.A(n25240), .B(n21067), .C(n25265), 
         .D(n25263), .Z(n21150)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_343.init = 16'h0040;
    PFUMX mux_1568_i15 (.BLUT(n2937[14]), .ALUT(n2890[14]), .C0(n3619), 
          .Z(n2978[14]));
    LUT4 i1_4_lut_4_lut_4_lut_adj_344 (.A(n25240), .B(n21067), .C(n25264), 
         .D(n25263), .Z(n21148)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_4_lut_adj_344.init = 16'h0040;
    PFUMX i22229 (.BLUT(n24661), .ALUT(n24660), .C0(counter_hi[2]), .Z(n24662));
    LUT4 next_pc_for_core_23__I_0_i157_3_lut (.A(\next_pc_for_core[8] ), .B(\next_pc_for_core[12] ), 
         .C(counter_hi[2]), .Z(n157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i157_3_lut.init = 16'hcaca;
    LUT4 i21952_3_lut_4_lut (.A(n26), .B(n25158), .C(n3605), .D(n3613), 
         .Z(n23220)) /* synthesis lut_function=(!(A (B (C+(D))))) */ ;
    defparam i21952_3_lut_4_lut.init = 16'h777f;
    LUT4 mux_345_i1_3_lut (.A(\next_pc_for_core[3] ), .B(return_addr[3]), 
         .C(debug_ret), .Z(n1742[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i1_3_lut.init = 16'hcaca;
    PFUMX mux_1568_i16 (.BLUT(n2937[15]), .ALUT(n2890[15]), .C0(n3619), 
          .Z(n2978[15]));
    LUT4 mux_1256_i16_3_lut (.A(n14[15]), .B(n2[15]), .C(n1949), .Z(n1950[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i16_3_lut.init = 16'hcaca;
    LUT4 i12007_2_lut_rep_470_3_lut (.A(n25281), .B(n26598), .C(instr[12]), 
         .Z(n25206)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12007_2_lut_rep_470_3_lut.init = 16'h4040;
    LUT4 mux_1260_i16_3_lut (.A(n7[15]), .B(n9[15]), .C(n1969), .Z(n1970[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i16_3_lut.init = 16'hcaca;
    LUT4 i12006_2_lut_3_lut (.A(n25281), .B(n26598), .C(n25264), .Z(n2736[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i12006_2_lut_3_lut.init = 16'h4040;
    L6MUX21 mux_1568_i17 (.D0(n2937[16]), .D1(n2890[16]), .SD(n3619), 
            .Z(n2978[16]));
    LUT4 mux_1540_i19_3_lut_3_lut_4_lut (.A(n26), .B(n25158), .C(n25206), 
         .D(n2813[10]), .Z(n2854[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1540_i19_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1517_i12_4_lut_4_lut_4_lut (.A(n25281), .B(n26598), .C(n3613), 
         .D(instr[12]), .Z(n2703[11])) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (C (D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1517_i12_4_lut_4_lut_4_lut.init = 16'h4300;
    LUT4 mux_1256_i1_3_lut (.A(n14[0]), .B(n2[0]), .C(n1949), .Z(n1950[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i1_3_lut.init = 16'hcaca;
    FD1P3IX data_addr__i1 (.D(addr_out[1]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i1.GSR = "DISABLED";
    LUT4 mux_1260_i1_3_lut (.A(n7[0]), .B(n9[0]), .C(n1969), .Z(n1970[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i1_3_lut.init = 16'hcaca;
    FD1P3IX data_addr__i2 (.D(n699[0]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i2.GSR = "DISABLED";
    FD1P3IX data_addr__i3 (.D(n21499), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i3.GSR = "DISABLED";
    FD1P3IX data_addr__i4 (.D(addr_out[4]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i4.GSR = "DISABLED";
    FD1P3IX data_addr__i5 (.D(addr_out[5]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i5.GSR = "DISABLED";
    FD1P3IX data_addr__i6 (.D(addr_out[6]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i6.GSR = "DISABLED";
    FD1P3IX data_addr__i7 (.D(addr_out[7]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i7.GSR = "DISABLED";
    FD1P3IX data_addr__i8 (.D(addr_out[8]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i8.GSR = "DISABLED";
    FD1P3IX data_addr__i9 (.D(addr_out[9]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i9.GSR = "DISABLED";
    FD1P3IX data_addr__i10 (.D(addr_out[10]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i10.GSR = "DISABLED";
    FD1P3IX data_addr__i11 (.D(addr_out[11]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i11.GSR = "DISABLED";
    FD1P3IX data_addr__i12 (.D(addr_out[12]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i12.GSR = "DISABLED";
    FD1P3IX data_addr__i13 (.D(addr_out[13]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i13.GSR = "DISABLED";
    FD1P3IX data_addr__i14 (.D(addr_out[14]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i14.GSR = "DISABLED";
    FD1P3IX data_addr__i15 (.D(addr_out[15]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i15.GSR = "DISABLED";
    FD1P3IX data_addr__i16 (.D(addr_out[16]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[16])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i16.GSR = "DISABLED";
    FD1P3IX data_addr__i17 (.D(addr_out[17]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[17])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i17.GSR = "DISABLED";
    FD1P3IX data_addr__i18 (.D(addr_out[18]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[18])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i18.GSR = "DISABLED";
    FD1P3IX data_addr__i19 (.D(addr_out[19]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[19])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i19.GSR = "DISABLED";
    FD1P3IX data_addr__i20 (.D(addr_out[20]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[20])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i20.GSR = "DISABLED";
    FD1P3IX data_addr__i21 (.D(addr_out[21]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[21])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i21.GSR = "DISABLED";
    FD1P3IX data_addr__i22 (.D(addr_out[22]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[22])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i22.GSR = "DISABLED";
    FD1P3IX data_addr__i23 (.D(addr_out[23]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[23])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i23.GSR = "DISABLED";
    FD1P3IX data_addr__i24 (.D(addr_out[24]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i24.GSR = "DISABLED";
    FD1P3IX data_addr__i25 (.D(addr_out[25]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i25.GSR = "DISABLED";
    FD1P3IX data_addr__i26 (.D(addr_out[26]), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i26.GSR = "DISABLED";
    FD1P3IX data_addr__i27 (.D(n25307), .SP(clk_c_enable_309), .CD(n25424), 
            .CK(clk_c), .Q(addr[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i27.GSR = "DISABLED";
    FD1P3AX rs2_i0_i1 (.D(n1729[1]), .SP(clk_c_enable_312), .CK(clk_c), 
            .Q(rs2[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i1.GSR = "DISABLED";
    FD1P3AX rs2_i0_i2 (.D(n1729[2]), .SP(clk_c_enable_312), .CK(clk_c), 
            .Q(rs2[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i2.GSR = "DISABLED";
    FD1P3AX rs2_i0_i3 (.D(n1729[3]), .SP(clk_c_enable_312), .CK(clk_c), 
            .Q(rs2[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i3.GSR = "DISABLED";
    FD1S3IX counter_hi_3136__i3 (.D(n17_adj_2394[1]), .CK(clk_c), .CD(n25424), 
            .Q(counter_hi[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3136__i3.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_adj_345 (.A(n26598), .B(n24), .C(n22286), .D(n22470), 
         .Z(n22172)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_4_lut_adj_345.init = 16'hf040;
    LUT4 mux_1522_i17_3_lut_4_lut (.A(n25167), .B(n25194), .C(n4548[9]), 
         .D(n22996), .Z(n2772[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1522_i17_3_lut_4_lut.init = 16'hf870;
    LUT4 i21809_4_lut (.A(n25182), .B(n20952), .C(n25336), .D(n22010), 
         .Z(clk_c_enable_219)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i21809_4_lut.init = 16'h0010;
    LUT4 mux_1540_i13_3_lut_3_lut_4_lut (.A(n26), .B(n25158), .C(n4608[11]), 
         .D(n2813[10]), .Z(n2854[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1540_i13_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1026_i1_4_lut (.A(n25265), .B(rs2[0]), .C(n25178), .D(mem_op_increment_reg), 
         .Z(n1708[0])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1026_i1_4_lut.init = 16'h3aca;
    LUT4 n928_bdd_4_lut_22417_4_lut (.A(n26598), .B(n25279), .C(n25281), 
         .D(n25284), .Z(n24943)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam n928_bdd_4_lut_22417_4_lut.init = 16'h0040;
    LUT4 mux_1540_i14_3_lut_3_lut_4_lut (.A(n26), .B(n25158), .C(n4608[12]), 
         .D(n2813[10]), .Z(n2854[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1540_i14_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1540_i17_3_lut_3_lut_4_lut (.A(n26), .B(n25158), .C(n4608[15]), 
         .D(n2813[10]), .Z(n2854[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1540_i17_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i2_3_lut (.A(\next_pc_for_core[4] ), .B(return_addr[4]), 
         .C(debug_ret), .Z(n1742[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i2_3_lut.init = 16'hcaca;
    LUT4 i15_4_lut (.A(n66), .B(n12257), .C(clk_c_enable_206), .D(n25387), 
         .Z(no_write_in_progress_N_202)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i15_4_lut.init = 16'hcaaa;
    LUT4 mux_345_i3_3_lut (.A(\next_pc_for_core[5] ), .B(return_addr[5]), 
         .C(debug_ret), .Z(n1742[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i3_3_lut.init = 16'hcaca;
    LUT4 instr_1__bdd_4_lut_22434_4_lut (.A(n26598), .B(n26597), .C(n25279), 
         .D(n25284), .Z(n25004)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam instr_1__bdd_4_lut_22434_4_lut.init = 16'h0010;
    LUT4 mux_1007_i15_3_lut (.A(n9[14]), .B(n14[14]), .C(n1969), .Z(n1649[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i15_3_lut.init = 16'hcaca;
    LUT4 mux_29_i3_3_lut_4_lut_4_lut (.A(n26598), .B(n155[2]), .C(n25216), 
         .D(n25239), .Z(alu_op_3__N_901[2])) /* synthesis lut_function=(A (B (C+(D)))+!A (B+!(C+(D)))) */ ;
    defparam mux_29_i3_3_lut_4_lut_4_lut.init = 16'hccc5;
    LUT4 mux_345_i4_3_lut (.A(\next_pc_for_core[6] ), .B(return_addr[6]), 
         .C(debug_ret), .Z(n1742[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i3_4_lut_4_lut (.A(n26598), .B(n3605), .C(n25284), .D(instr[4]), 
         .Z(n2703[2])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_1517_i3_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_1517_i6_4_lut_4_lut (.A(n26598), .B(n3605), .C(n25284), .D(n25265), 
         .Z(n2703[5])) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C+(D))+!B (D))) */ ;
    defparam mux_1517_i6_4_lut_4_lut.init = 16'hddc0;
    LUT4 mux_345_i5_3_lut (.A(\next_pc_for_core[7] ), .B(return_addr[7]), 
         .C(debug_ret), .Z(n1742[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i5_3_lut.init = 16'hcaca;
    PFUMX i22527 (.BLUT(n25444), .ALUT(n25445), .C0(n25338), .Z(instr[31]));
    LUT4 mux_1007_i2_3_lut (.A(n9[1]), .B(n14[1]), .C(n1969), .Z(n1649[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i2_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n25372), .B(cmp), .C(alu_b_in[1]), .D(alu_a_in[1]), 
         .Z(n21812)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd00d;
    LUT4 mux_1517_i4_4_lut_4_lut (.A(n26598), .B(n3605), .C(n25284), .D(n25267), 
         .Z(n2703[3])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_1517_i4_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_345_i6_3_lut (.A(\next_pc_for_core[8] ), .B(return_addr[8]), 
         .C(debug_ret), .Z(n1742[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i6_3_lut.init = 16'hcaca;
    LUT4 mux_345_i7_3_lut (.A(\next_pc_for_core[9] ), .B(return_addr[9]), 
         .C(debug_ret), .Z(n1742[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i7_3_lut.init = 16'hcaca;
    LUT4 mux_345_i8_3_lut (.A(\next_pc_for_core[10] ), .B(return_addr[10]), 
         .C(debug_ret), .Z(n1742[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i8_3_lut.init = 16'hcaca;
    LUT4 mux_1266_i2_rep_127_3_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .Z(n23899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i2_rep_127_3_lut.init = 16'hcaca;
    LUT4 mux_1517_i2_4_lut_4_lut (.A(n26598), .B(n3605), .C(n25284), .D(n25264), 
         .Z(n2703[1])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_1517_i2_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_345_i9_3_lut (.A(\next_pc_for_core[11] ), .B(return_addr[11]), 
         .C(debug_ret), .Z(n1742[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i9_3_lut.init = 16'hcaca;
    PFUMX mux_1531_i6 (.BLUT(n2627[5]), .ALUT(n21260), .C0(n3611), .Z(n2813[5]));
    FD1S3IX counter_hi_3136__i4 (.D(n17_adj_2394[2]), .CK(clk_c), .CD(n25424), 
            .Q(counter_hi[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3136__i4.GSR = "DISABLED";
    FD1S3IX addr_offset_3137__i3 (.D(n22878), .CK(clk_c), .CD(n25424), 
            .Q(addr_offset[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam addr_offset_3137__i3.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_459_4_lut (.A(n25284), .B(n25279), .C(n26598), .D(n25210), 
         .Z(n25195)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_3_lut_rep_459_4_lut.init = 16'h0002;
    LUT4 mux_345_i10_3_lut (.A(\next_pc_for_core[12] ), .B(return_addr[12]), 
         .C(debug_ret), .Z(n1742[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i10_3_lut.init = 16'hcaca;
    LUT4 mux_345_i11_3_lut (.A(\next_pc_for_core[13] ), .B(return_addr[13]), 
         .C(debug_ret), .Z(n1742[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i11_3_lut.init = 16'hcaca;
    LUT4 is_alu_imm_N_1098_bdd_3_lut_4_lut_4_lut (.A(n25279), .B(n26598), 
         .C(n25260), .D(n25290), .Z(n24919)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;
    defparam is_alu_imm_N_1098_bdd_3_lut_4_lut_4_lut.init = 16'h5d55;
    LUT4 i1_4_lut_adj_346 (.A(n21575), .B(n25417), .C(addr[3]), .D(addr[6]), 
         .Z(is_timer_addr)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_346.init = 16'h0002;
    LUT4 i1_4_lut_adj_347 (.A(n22646), .B(addr[7]), .C(n22648), .D(n22644), 
         .Z(n21575)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_347.init = 16'h2000;
    LUT4 i1_4_lut_adj_348 (.A(addr[13]), .B(n22636), .C(n22622), .D(addr[14]), 
         .Z(n22646)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_348.init = 16'h8000;
    LUT4 mux_1266_i2_rep_128_3_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .Z(n23900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i2_rep_128_3_lut.init = 16'hcaca;
    PFUMX mux_1559_i17 (.BLUT(n2703[16]), .ALUT(n2854[16]), .C0(n23220), 
          .Z(n2937[16]));
    LUT4 mux_345_i12_3_lut (.A(\next_pc_for_core[14] ), .B(return_addr[14]), 
         .C(debug_ret), .Z(n1742[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1540_i15_3_lut_3_lut_4_lut (.A(n26), .B(n25158), .C(n4608[13]), 
         .D(n2813[10]), .Z(n2854[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1540_i15_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i13_3_lut (.A(\next_pc_for_core[15] ), .B(return_addr[15]), 
         .C(debug_ret), .Z(n1742[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i13_3_lut.init = 16'hcaca;
    LUT4 mux_345_i14_3_lut (.A(\next_pc_for_core[16] ), .B(return_addr[16]), 
         .C(debug_ret), .Z(n1742[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1540_i11_3_lut_3_lut_4_lut (.A(n26), .B(n25158), .C(n2703[10]), 
         .D(n2813[10]), .Z(n2854[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1540_i11_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i15_3_lut (.A(\next_pc_for_core[17] ), .B(return_addr[17]), 
         .C(debug_ret), .Z(n1742[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i15_3_lut.init = 16'hcaca;
    PFUMX mux_1559_i8 (.BLUT(n2813[7]), .ALUT(n2854[7]), .C0(n25155), 
          .Z(n2937[7]));
    LUT4 mux_345_i16_3_lut (.A(\next_pc_for_core[18] ), .B(return_addr[18]), 
         .C(debug_ret), .Z(n1742[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1256_i2_3_lut (.A(n14[1]), .B(n2[1]), .C(n1949), .Z(n1950[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_349 (.A(n22638), .B(n22620), .C(addr[8]), .D(addr[25]), 
         .Z(n22648)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_349.init = 16'h8000;
    LUT4 mux_1540_i12_3_lut_3_lut_4_lut (.A(n26), .B(n25158), .C(n2703[11]), 
         .D(n2813[10]), .Z(n2854[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1540_i12_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1260_i2_3_lut (.A(n7[1]), .B(n9[1]), .C(n1969), .Z(n1970[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i2_3_lut.init = 16'hcaca;
    LUT4 mux_345_i17_3_lut (.A(\next_pc_for_core[19] ), .B(return_addr[19]), 
         .C(debug_ret), .Z(n1742[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i17_3_lut.init = 16'hcaca;
    L6MUX21 mux_1559_i7 (.D0(n2813[6]), .D1(n2854[6]), .SD(n25155), .Z(n2937[6]));
    L6MUX21 mux_1559_i4 (.D0(n2813[3]), .D1(n2854[3]), .SD(n25155), .Z(n2937[3]));
    LUT4 i1_4_lut_adj_350 (.A(addr[24]), .B(addr[26]), .C(addr[27]), .D(addr[23]), 
         .Z(n22644)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_350.init = 16'h8000;
    L6MUX21 mux_1559_i2 (.D0(n2813[1]), .D1(n2854[1]), .SD(n25155), .Z(n2937[1]));
    PFUMX mux_1323_i3 (.BLUT(n21269), .ALUT(n2075[2]), .C0(n2244), .Z(n2089[2]));
    LUT4 mux_1256_i15_3_lut (.A(n14[14]), .B(n2[14]), .C(n1949), .Z(n1950[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i15_3_lut.init = 16'hcaca;
    LUT4 mux_345_i18_3_lut (.A(\next_pc_for_core[20] ), .B(return_addr[20]), 
         .C(debug_ret), .Z(n1742[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i18_3_lut.init = 16'hcaca;
    LUT4 mux_1512_i2_4_lut_4_lut (.A(n25279), .B(n3603), .C(n25264), .D(n25267), 
         .Z(n2666[1])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;
    defparam mux_1512_i2_4_lut_4_lut.init = 16'h7340;
    LUT4 i1_4_lut_adj_351 (.A(addr[17]), .B(addr[15]), .C(addr[18]), .D(addr[21]), 
         .Z(n22636)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_351.init = 16'h8000;
    LUT4 mux_1260_i15_3_lut (.A(n7[14]), .B(n9[14]), .C(n1969), .Z(n1970[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i15_3_lut.init = 16'hcaca;
    LUT4 mux_345_i19_3_lut (.A(\next_pc_for_core[21] ), .B(return_addr[21]), 
         .C(debug_ret), .Z(n1742[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i19_3_lut.init = 16'hcaca;
    FD1P3AX data_write_n_i1 (.D(data_write_n_1__N_100[1]), .SP(clk_c_enable_314), 
            .CK(clk_c), .Q(qv_data_write_n[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_write_n_i1.GSR = "DISABLED";
    LUT4 i53_4_lut_4_lut (.A(n25279), .B(n25281), .C(n25211), .D(n26597), 
         .Z(n32)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam i53_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_345_i20_3_lut (.A(\next_pc_for_core[22] ), .B(return_addr[22]), 
         .C(debug_ret), .Z(n1742[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i20_3_lut.init = 16'hcaca;
    LUT4 mem_data_from_read_6__bdd_3_lut_22389_then_4_lut (.A(data_txn_len[0]), 
         .B(\qspi_data_buf[14] ), .C(instr_data[14]), .D(n25253), .Z(n25442)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B)) */ ;
    defparam mem_data_from_read_6__bdd_3_lut_22389_then_4_lut.init = 16'he4cc;
    FD1P3IX pc_offset__i21 (.D(pc_23__N_642[18]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[21] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i21.GSR = "DISABLED";
    FD1P3IX pc_offset__i22 (.D(pc_23__N_642[19]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[22] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i22.GSR = "DISABLED";
    FD1P3IX pc_offset__i23 (.D(pc_23__N_642[20]), .SP(clk_c_enable_393), 
            .CD(n25424), .CK(clk_c), .Q(\pc[23] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i23.GSR = "DISABLED";
    LUT4 i12041_4_lut_4_lut (.A(n25279), .B(n26598), .C(n25255), .D(alu_op_3__N_1068[2]), 
         .Z(n15_adj_2380)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i12041_4_lut_4_lut.init = 16'hd0c0;
    LUT4 mux_345_i21_3_lut (.A(\next_pc_for_core[23] ), .B(return_addr[23]), 
         .C(debug_ret), .Z(n1742[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i21_3_lut.init = 16'hcaca;
    PFUMX mux_1531_i9 (.BLUT(n21157), .ALUT(n21242), .C0(n3611), .Z(n2813[8]));
    LUT4 mux_1540_i16_3_lut_3_lut_4_lut (.A(n26), .B(n25158), .C(n4608[14]), 
         .D(n2813[10]), .Z(n2854[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1540_i16_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1256_i14_3_lut (.A(n14[13]), .B(n2[13]), .C(n1949), .Z(n1950[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1260_i14_3_lut (.A(n7[13]), .B(n9[13]), .C(n1969), .Z(n1970[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i14_3_lut.init = 16'hcaca;
    LUT4 i42_4_lut_4_lut (.A(n25279), .B(n26598), .C(n26597), .D(n25281), 
         .Z(n27_adj_2381)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C)))) */ ;
    defparam i42_4_lut_4_lut.init = 16'h404a;
    LUT4 mem_data_from_read_6__bdd_3_lut_22389_else_4_lut (.A(data_txn_len[0]), 
         .B(n25253), .C(instr_data[10]), .D(\qspi_data_buf[10] ), .Z(n25441)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mem_data_from_read_6__bdd_3_lut_22389_else_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_352 (.A(addr[9]), .B(addr[20]), .Z(n22622)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_352.init = 16'h8888;
    LUT4 i1_4_lut_adj_353 (.A(addr[19]), .B(addr[10]), .C(addr[12]), .D(addr[11]), 
         .Z(n22638)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_353.init = 16'h8000;
    LUT4 mux_1026_i2_4_lut (.A(n25264), .B(rs2[1]), .C(n25178), .D(n25429), 
         .Z(n1708[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1026_i2_4_lut.init = 16'h3aca;
    LUT4 mux_1026_i3_4_lut (.A(instr[4]), .B(rs2[2]), .C(n25178), .D(n25368), 
         .Z(n1708[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1026_i3_4_lut.init = 16'h3aca;
    LUT4 mux_1007_i13_3_lut (.A(n9[12]), .B(n14[12]), .C(n1969), .Z(n1649[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i13_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_354 (.A(addr[22]), .B(addr[16]), .Z(n22620)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_354.init = 16'h8888;
    LUT4 i20795_3_lut_4_lut (.A(n25419), .B(n25418), .C(counter_hi[2]), 
         .D(\next_pc_for_core[6] ), .Z(n23070)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i20795_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_1026_i4_4_lut (.A(n25267), .B(rs2[3]), .C(n25178), .D(n5570), 
         .Z(n1708[3])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1026_i4_4_lut.init = 16'h3aca;
    LUT4 mux_1256_i12_3_lut (.A(n14[11]), .B(n2[11]), .C(n1949), .Z(n1950[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i12_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_3_lut_4_lut (.A(n22), .B(n25158), .C(n25288), .D(rst_reg_n), 
         .Z(n21157)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam i1_3_lut_3_lut_4_lut.init = 16'h7000;
    PFUMX mux_1531_i7 (.BLUT(n2627[6]), .ALUT(n21248), .C0(n3611), .Z(n2813[6]));
    LUT4 mux_1260_i12_3_lut (.A(n7[11]), .B(n9[11]), .C(n1969), .Z(n1970[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i12_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(any_additional_mem_ops), .B(n25180), .C(n26612), 
         .Z(n21369)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i3851_2_lut_3_lut_4_lut (.A(n25419), .B(n25418), .C(n25420), 
         .D(instr_addr_23__N_49[0]), .Z(n5879)) /* synthesis lut_function=(A (B ((D)+!C))+!A !(B+!((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i3851_2_lut_3_lut_4_lut.init = 16'h9909;
    LUT4 n3601_bdd_3_lut_22143_4_lut (.A(n22), .B(n25158), .C(rst_reg_n), 
         .D(n25287), .Z(n24488)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam n3601_bdd_3_lut_22143_4_lut.init = 16'h7000;
    LUT4 i5262_4_lut (.A(n22978), .B(instr[26]), .C(n3615), .D(n25209), 
         .Z(n2772[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i5262_4_lut.init = 16'hca0a;
    LUT4 mux_347_i2_3_lut_4_lut (.A(n25419), .B(n25418), .C(debug_ret), 
         .D(return_addr[2]), .Z(n1768[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam mux_347_i2_3_lut_4_lut.init = 16'hf606;
    LUT4 i1_2_lut_adj_355 (.A(n25179), .B(n7955), .Z(n22126)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_355.init = 16'heeee;
    LUT4 i21542_4_lut_4_lut (.A(n25381), .B(n23395), .C(n234[0]), .D(debug_branch_N_177[28]), 
         .Z(debug_rd_3__N_1298[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i21542_4_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_356 (.A(n25279), .B(n25281), .C(n25267), .D(n26597), 
         .Z(n21960)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_356.init = 16'h0010;
    PFUMX mux_1531_i4 (.BLUT(n2627[3]), .ALUT(n21113), .C0(n3611), .Z(n2813[3]));
    LUT4 i1_3_lut_4_lut_adj_357 (.A(n25279), .B(n25281), .C(n25287), .D(n26597), 
         .Z(n21954)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_357.init = 16'h0010;
    PFUMX mux_1531_i2 (.BLUT(n2627[1]), .ALUT(n2666[1]), .C0(n3611), .Z(n2813[1]));
    PFUMX i22206 (.BLUT(n24617), .ALUT(n24616), .C0(counter_hi[2]), .Z(n24618));
    LUT4 i20789_3_lut (.A(\mem_data_from_read[19] ), .B(\mem_data_from_read[23] ), 
         .C(counter_hi[2]), .Z(n23064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20789_3_lut.init = 16'hcaca;
    LUT4 n24564_bdd_3_lut (.A(n24564), .B(n25290), .C(n3597), .Z(n24565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24564_bdd_3_lut.init = 16'hcaca;
    PFUMX mux_1540_i7 (.BLUT(n2703[6]), .ALUT(n2736[6]), .C0(n3613), .Z(n2854[6]));
    LUT4 i1_4_lut_adj_358 (.A(any_additional_mem_ops), .B(n25180), .C(rd[1]), 
         .D(rd[0]), .Z(n21374)) /* synthesis lut_function=(!(((C (D)+!C !(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i1_4_lut_adj_358.init = 16'h0880;
    PFUMX mux_1540_i6 (.BLUT(n2703[5]), .ALUT(n2736[5]), .C0(n3613), .Z(n2854[5]));
    LUT4 mux_1522_i12_3_lut_4_lut (.A(n3615), .B(n25167), .C(n4548[4]), 
         .D(n22959), .Z(n2772[11])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1522_i12_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_4_lut_adj_359 (.A(rd[2]), .B(n25180), .C(any_additional_mem_ops), 
         .D(n25434), .Z(n21375)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i1_4_lut_adj_359.init = 16'h4080;
    LUT4 i1_4_lut_adj_360 (.A(rd[3]), .B(n25180), .C(any_additional_mem_ops), 
         .D(n5599), .Z(n21376)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i1_4_lut_adj_360.init = 16'h4080;
    LUT4 n3597_bdd_4_lut_22186 (.A(n25258), .B(n22968), .C(n22957), .D(n25338), 
         .Z(n24566)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n3597_bdd_4_lut_22186.init = 16'h88a0;
    LUT4 i21814_4_lut (.A(n25182), .B(rst_reg_n), .C(n20952), .D(n21962), 
         .Z(clk_c_enable_29)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i21814_4_lut.init = 16'h3337;
    LUT4 i6512_3_lut (.A(n26598), .B(n25290), .C(n25260), .Z(n8768)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam i6512_3_lut.init = 16'h4c4c;
    LUT4 i12035_2_lut_3_lut_4_lut (.A(n26598), .B(n25279), .C(instr[4]), 
         .D(n25257), .Z(n15_adj_2382)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i12035_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i31_4_lut_4_lut (.A(n25284), .B(n26598), .C(n20641), .D(n25279), 
         .Z(n25)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(C+(D))))) */ ;
    defparam i31_4_lut_4_lut.init = 16'h11fc;
    LUT4 i2_3_lut_4_lut_3_lut_4_lut (.A(n25284), .B(n26598), .C(n25279), 
         .D(n25258), .Z(n6)) /* synthesis lut_function=(A (D)+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i2_3_lut_4_lut_3_lut_4_lut.init = 16'hff01;
    LUT4 i6507_3_lut_4_lut (.A(addr[27]), .B(n25431), .C(\data_from_read[2] ), 
         .D(n23405), .Z(debug_branch_N_571[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i6507_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21823_3_lut_rep_588_4_lut (.A(addr[27]), .B(n25431), .C(n25432), 
         .D(n17512), .Z(n25324)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i21823_3_lut_rep_588_4_lut.init = 16'h0111;
    LUT4 i20791_3_lut_4_lut (.A(addr[27]), .B(n25431), .C(\data_from_read[2] ), 
         .D(n23064), .Z(n23066)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i20791_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21675_3_lut (.A(n2772[12]), .B(n4516[12]), .C(n3615), .Z(n2890[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21675_3_lut.init = 16'hcaca;
    LUT4 i21673_3_lut (.A(n2772[13]), .B(n4516[13]), .C(n3615), .Z(n2890[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21673_3_lut.init = 16'hcaca;
    LUT4 i21671_3_lut (.A(n2772[14]), .B(n4516[14]), .C(n3615), .Z(n2890[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21671_3_lut.init = 16'hcaca;
    LUT4 i52_4_lut_4_lut (.A(n26597), .B(n25279), .C(n13814), .D(n26598), 
         .Z(n37)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (D)+!B !(C+(D))))) */ ;
    defparam i52_4_lut_4_lut.init = 16'h4403;
    LUT4 i1_2_lut_3_lut_4_lut_adj_361 (.A(addr[27]), .B(n25431), .C(addr[3]), 
         .D(n25432), .Z(n20582)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_4_lut_adj_361.init = 16'h00e0;
    LUT4 i21669_3_lut (.A(n2772[15]), .B(n4516[15]), .C(n3615), .Z(n2890[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21669_3_lut.init = 16'hcaca;
    LUT4 i20783_3_lut (.A(\mem_data_from_read[16] ), .B(\mem_data_from_read[20] ), 
         .C(counter_hi[2]), .Z(n23058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20783_3_lut.init = 16'hcaca;
    LUT4 i20786_3_lut (.A(\mem_data_from_read[18] ), .B(\mem_data_from_read[22] ), 
         .C(counter_hi[2]), .Z(n23061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20786_3_lut.init = 16'hcaca;
    LUT4 i20785_3_lut_4_lut (.A(addr[27]), .B(n25431), .C(\data_from_read[2] ), 
         .D(n23058), .Z(n23060)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i20785_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i20695_3_lut_rep_504 (.A(n25281), .B(n25279), .C(n26597), .Z(n25240)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i20695_3_lut_rep_504.init = 16'hfefe;
    LUT4 i20788_3_lut_4_lut (.A(addr[27]), .B(n25431), .C(\data_from_read[2] ), 
         .D(n23061), .Z(n23063)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i20788_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2_2_lut_4_lut (.A(n25281), .B(n25279), .C(n26597), .D(n21212), 
         .Z(n3589)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_2_lut_4_lut.init = 16'h0100;
    LUT4 i20780_3_lut_4_lut (.A(addr[27]), .B(n25431), .C(\data_from_read[2] ), 
         .D(\mem_data_from_read[3] ), .Z(n23055)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i20780_3_lut_4_lut.init = 16'hf1e0;
    PFUMX mux_1540_i4 (.BLUT(n2703[3]), .ALUT(n2736[3]), .C0(n3613), .Z(n2854[3]));
    LUT4 i6479_3_lut_4_lut (.A(addr[27]), .B(n25431), .C(\data_from_read[2] ), 
         .D(n23039), .Z(n8735)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i6479_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX data_out__i1 (.D(data_out_slice[1]), .SP(clk_c_enable_324), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i1.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_362 (.A(addr[27]), .B(n25431), .C(qv_data_read_n[1]), 
         .D(qv_data_read_n[0]), .Z(read_en)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_3_lut_4_lut_adj_362.init = 16'h00e0;
    FD1P3IX data_out__i2 (.D(data_out_slice[2]), .SP(clk_c_enable_324), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i2.GSR = "DISABLED";
    FD1P3IX data_out__i3 (.D(n25277), .SP(clk_c_enable_324), .CD(n25424), 
            .CK(clk_c), .Q(data_to_write[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i3.GSR = "DISABLED";
    FD1P3IX data_out__i4 (.D(data_out_slice[0]), .SP(clk_c_enable_328), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i4.GSR = "DISABLED";
    FD1P3IX data_out__i5 (.D(data_out_slice[1]), .SP(clk_c_enable_328), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i5.GSR = "DISABLED";
    FD1P3IX data_out__i6 (.D(data_out_slice[2]), .SP(clk_c_enable_328), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i6.GSR = "DISABLED";
    FD1P3IX data_out__i7 (.D(n25277), .SP(clk_c_enable_328), .CD(n25424), 
            .CK(clk_c), .Q(data_to_write[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i7.GSR = "DISABLED";
    FD1P3IX data_out__i8 (.D(data_out_slice[0]), .SP(clk_c_enable_332), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i8.GSR = "DISABLED";
    FD1P3IX data_out__i9 (.D(data_out_slice[1]), .SP(clk_c_enable_332), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i9.GSR = "DISABLED";
    FD1P3IX data_out__i10 (.D(data_out_slice[2]), .SP(clk_c_enable_332), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i10.GSR = "DISABLED";
    FD1P3IX data_out__i11 (.D(n25277), .SP(clk_c_enable_332), .CD(n25424), 
            .CK(clk_c), .Q(data_to_write[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i11.GSR = "DISABLED";
    FD1P3IX data_out__i12 (.D(data_out_slice[0]), .SP(clk_c_enable_336), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i12.GSR = "DISABLED";
    FD1P3IX data_out__i13 (.D(data_out_slice[1]), .SP(clk_c_enable_336), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i13.GSR = "DISABLED";
    FD1P3IX data_out__i14 (.D(data_out_slice[2]), .SP(clk_c_enable_336), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i14.GSR = "DISABLED";
    FD1P3IX data_out__i15 (.D(n25277), .SP(clk_c_enable_336), .CD(n25424), 
            .CK(clk_c), .Q(data_to_write[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i15.GSR = "DISABLED";
    FD1P3IX data_out__i16 (.D(data_out_slice[0]), .SP(clk_c_enable_340), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[16])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i16.GSR = "DISABLED";
    FD1P3IX data_out__i17 (.D(data_out_slice[1]), .SP(clk_c_enable_340), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[17])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i17.GSR = "DISABLED";
    FD1P3IX data_out__i18 (.D(data_out_slice[2]), .SP(clk_c_enable_340), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[18])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i18.GSR = "DISABLED";
    FD1P3IX data_out__i19 (.D(n25277), .SP(clk_c_enable_340), .CD(n25424), 
            .CK(clk_c), .Q(data_to_write[19])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i19.GSR = "DISABLED";
    FD1P3IX data_out__i20 (.D(data_out_slice[0]), .SP(clk_c_enable_344), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[20])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i20.GSR = "DISABLED";
    FD1P3IX data_out__i21 (.D(data_out_slice[1]), .SP(clk_c_enable_344), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[21])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i21.GSR = "DISABLED";
    FD1P3IX data_out__i22 (.D(data_out_slice[2]), .SP(clk_c_enable_344), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[22])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i22.GSR = "DISABLED";
    FD1P3IX data_out__i23 (.D(n25277), .SP(clk_c_enable_344), .CD(n25424), 
            .CK(clk_c), .Q(data_to_write[23])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i23.GSR = "DISABLED";
    FD1P3IX data_out__i24 (.D(data_out_slice[0]), .SP(clk_c_enable_348), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i24.GSR = "DISABLED";
    FD1P3IX data_out__i25 (.D(data_out_slice[1]), .SP(clk_c_enable_348), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i25.GSR = "DISABLED";
    FD1P3IX data_out__i26 (.D(data_out_slice[2]), .SP(clk_c_enable_348), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i26.GSR = "DISABLED";
    FD1P3IX data_out__i27 (.D(n25277), .SP(clk_c_enable_348), .CD(n25424), 
            .CK(clk_c), .Q(data_to_write[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i27.GSR = "DISABLED";
    FD1P3IX data_out__i28 (.D(data_out_slice[0]), .SP(clk_c_enable_352), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i28.GSR = "DISABLED";
    FD1P3IX data_out__i29 (.D(data_out_slice[1]), .SP(clk_c_enable_352), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i29.GSR = "DISABLED";
    FD1P3IX data_out__i30 (.D(data_out_slice[2]), .SP(clk_c_enable_352), 
            .CD(n25424), .CK(clk_c), .Q(data_to_write[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i30.GSR = "DISABLED";
    FD1P3IX data_out__i31 (.D(n25277), .SP(clk_c_enable_352), .CD(n25424), 
            .CK(clk_c), .Q(data_to_write[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i31.GSR = "DISABLED";
    LUT4 mux_1313_i4_4_lut (.A(n2047[3]), .B(instr[18]), .C(n2242), .D(n25258), 
         .Z(n2075[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam mux_1313_i4_4_lut.init = 16'hca0a;
    PFUMX mux_1540_i2 (.BLUT(n2703[1]), .ALUT(n2736[1]), .C0(n3613), .Z(n2854[1]));
    LUT4 n3597_bdd_3_lut_22183 (.A(n22968), .B(n22957), .C(n25338), .Z(n24564)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n3597_bdd_3_lut_22183.init = 16'hacac;
    LUT4 mux_1013_i16_3_lut_then_3_lut (.A(n14[15]), .B(n9[15]), .C(n1969), 
         .Z(n25445)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i16_3_lut_then_3_lut.init = 16'hacac;
    LUT4 mux_1013_i16_3_lut_else_3_lut (.A(n2[15]), .B(n7[15]), .C(n1949), 
         .Z(n25444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i16_3_lut_else_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_363 (.A(n25263), .B(n21067), .C(n25240), .Z(n21153)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_3_lut_adj_363.init = 16'h0404;
    FD1P3AX imm_i0_i1 (.D(n2978[1]), .SP(clk_c_enable_368), .CK(clk_c), 
            .Q(\imm[1] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i1.GSR = "DISABLED";
    LUT4 i16407_3_lut_4_lut (.A(n25178), .B(n25175), .C(n22126), .D(addr_offset[2]), 
         .Z(n17[0])) /* synthesis lut_function=(!(A (D)+!A !(B (C (D))+!B (D)))) */ ;
    defparam i16407_3_lut_4_lut.init = 16'h51aa;
    LUT4 equal_148_i4_2_lut_rep_639 (.A(counter_hi[3]), .B(counter_hi[4]), 
         .Z(n25375)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam equal_148_i4_2_lut_rep_639.init = 16'hbbbb;
    PFUMX mux_1544_i4 (.BLUT(n22962), .ALUT(n2772[3]), .C0(n23265), .Z(n2890[3]));
    LUT4 equal_149_i5_2_lut_rep_612_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(n25348)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam equal_149_i5_2_lut_rep_612_3_lut.init = 16'hfbfb;
    PFUMX mux_1544_i3 (.BLUT(n22960), .ALUT(n2772[2]), .C0(n23265), .Z(n2890[2]));
    LUT4 mux_1522_i5_3_lut (.A(n25278), .B(instr[24]), .C(n25166), .Z(n2772[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1522_i5_3_lut.init = 16'hcaca;
    LUT4 i21820_2_lut_3_lut (.A(n26610), .B(n26608), .C(counter_hi[2]), 
         .Z(n11558)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i21820_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_4_lut_adj_364 (.A(n25177), .B(n20807), .C(n8), .D(n22112), 
         .Z(n20739)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam i1_4_lut_adj_364.init = 16'h3b33;
    LUT4 i1_3_lut_4_lut_3_lut (.A(n25281), .B(n26597), .C(n25284), .Z(n20)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'hd9d9;
    LUT4 i1_2_lut_adj_365 (.A(is_ret_de), .B(n26612), .Z(n22112)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_365.init = 16'h8888;
    LUT4 i21870_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n25350), .D(counter_hi[2]), .Z(clk_c_enable_340)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i21870_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i3828_2_lut_3_lut (.A(instr_addr_23__N_49[0]), .B(\pc[1] ), .C(\pc[2] ), 
         .Z(n5856)) /* synthesis lut_function=(!(A (C)+!A (B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i3828_2_lut_3_lut.init = 16'h0b0b;
    LUT4 i1_2_lut_3_lut_adj_366 (.A(instr_addr_23__N_49[0]), .B(\pc[1] ), 
         .C(\pc[2] ), .Z(n21390)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i1_2_lut_3_lut_adj_366.init = 16'hbfbf;
    LUT4 i1_3_lut_4_lut_adj_367 (.A(n25209), .B(n25202), .C(n25208), .D(n7955), 
         .Z(n22098)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_adj_367.init = 16'h0070;
    LUT4 mux_1013_i5_rep_75_3_lut (.A(n22970), .B(n25289), .C(n3597), 
         .Z(n22954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i5_rep_75_3_lut.init = 16'hcaca;
    PFUMX mux_1559_i20 (.BLUT(n2703[17]), .ALUT(n2854[19]), .C0(n23341), 
          .Z(n2937[17]));
    LUT4 i11632_2_lut_3_lut (.A(n25281), .B(n26597), .C(n15_adj_2383), 
         .Z(mem_op_de[0])) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam i11632_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i1_3_lut_4_lut_adj_368 (.A(instr_addr_23__N_49[0]), .B(\pc[1] ), 
         .C(\pc[2] ), .D(instr_addr_23__N_49[1]), .Z(n21430)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i1_3_lut_4_lut_adj_368.init = 16'hb44b;
    LUT4 i11814_2_lut_3_lut_4_lut (.A(n25281), .B(n26597), .C(n25227), 
         .D(n25195), .Z(is_jalr_N_1101)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i11814_2_lut_3_lut_4_lut.init = 16'h2000;
    FD1P3AX imm_i0_i2 (.D(n25121), .SP(clk_c_enable_368), .CK(clk_c), 
            .Q(\imm[2] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i2.GSR = "DISABLED";
    FD1P3AX imm_i0_i3 (.D(n2978[3]), .SP(clk_c_enable_368), .CK(clk_c), 
            .Q(\imm[3] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i3.GSR = "DISABLED";
    FD1P3AX imm_i0_i4 (.D(n2978[4]), .SP(clk_c_enable_368), .CK(clk_c), 
            .Q(\imm[4] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i4.GSR = "DISABLED";
    FD1P3AX imm_i0_i5 (.D(n2978[5]), .SP(clk_c_enable_368), .CK(clk_c), 
            .Q(\imm[5] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i5.GSR = "DISABLED";
    FD1P3AX imm_i0_i6 (.D(n2978[6]), .SP(clk_c_enable_368), .CK(clk_c), 
            .Q(\imm[6] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i6.GSR = "DISABLED";
    FD1P3AX imm_i0_i7 (.D(n2978[7]), .SP(clk_c_enable_368), .CK(clk_c), 
            .Q(\imm[7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i7.GSR = "DISABLED";
    FD1P3AX imm_i0_i8 (.D(n2978[8]), .SP(clk_c_enable_370), .CK(clk_c), 
            .Q(\imm[8] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i8.GSR = "DISABLED";
    FD1P3AX imm_i0_i9 (.D(n2978[9]), .SP(clk_c_enable_370), .CK(clk_c), 
            .Q(\imm[9] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i9.GSR = "DISABLED";
    FD1P3AX imm_i0_i10 (.D(n2978[10]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[10] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i10.GSR = "DISABLED";
    FD1P3AX imm_i0_i11 (.D(n2978[11]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[11] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i11.GSR = "DISABLED";
    FD1P3AX imm_i0_i12 (.D(n2978[12]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[12] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i12.GSR = "DISABLED";
    FD1P3AX imm_i0_i13 (.D(n2978[13]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[13] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i13.GSR = "DISABLED";
    FD1P3AX imm_i0_i14 (.D(n2978[14]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[14] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i14.GSR = "DISABLED";
    FD1P3AX imm_i0_i15 (.D(n2978[15]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[15] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i15.GSR = "DISABLED";
    FD1P3AX imm_i0_i16 (.D(n2978[16]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[16] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i16.GSR = "DISABLED";
    FD1P3AX imm_i0_i17 (.D(n24425), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[17] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i17.GSR = "DISABLED";
    FD1P3AX imm_i0_i18 (.D(n24432), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i18.GSR = "DISABLED";
    FD1P3AX imm_i0_i19 (.D(n24453), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i19.GSR = "DISABLED";
    FD1P3AX imm_i0_i20 (.D(n2978[20]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i20.GSR = "DISABLED";
    FD1P3AX imm_i0_i21 (.D(n2978[21]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i21.GSR = "DISABLED";
    FD1P3AX imm_i0_i22 (.D(n2978[22]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i22.GSR = "DISABLED";
    FD1P3AX imm_i0_i23 (.D(n2978[23]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(\imm[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i23.GSR = "DISABLED";
    FD1P3AX imm_i0_i24 (.D(n2978[24]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(imm[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i24.GSR = "DISABLED";
    FD1P3AX imm_i0_i25 (.D(n2978[25]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(imm[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i25.GSR = "DISABLED";
    FD1P3AX imm_i0_i26 (.D(n2978[26]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(imm[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i26.GSR = "DISABLED";
    FD1P3AX imm_i0_i27 (.D(n2978[27]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(imm[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i27.GSR = "DISABLED";
    FD1P3AX imm_i0_i28 (.D(n2978[28]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(imm[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i28.GSR = "DISABLED";
    FD1P3AX imm_i0_i29 (.D(n2978[29]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(imm[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i29.GSR = "DISABLED";
    FD1P3AX imm_i0_i30 (.D(n24457), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(imm[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i30.GSR = "DISABLED";
    FD1P3AX imm_i0_i31 (.D(n4516[21]), .SP(clk_c_enable_392), .CK(clk_c), 
            .Q(imm[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i31.GSR = "DISABLED";
    LUT4 i21806_4_lut (.A(n25182), .B(n20952), .C(n25336), .D(n22016), 
         .Z(clk_c_enable_72)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i21806_4_lut.init = 16'h0010;
    LUT4 i2_2_lut_3_lut (.A(n25281), .B(n26597), .C(n25284), .Z(n11)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_2_lut_3_lut.init = 16'h2020;
    LUT4 i21677_3_lut (.A(n22954), .B(n2772[11]), .C(n23271), .Z(n2890[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21677_3_lut.init = 16'hcaca;
    LUT4 is_jalr_N_1103_bdd_2_lut_3_lut (.A(n25281), .B(n26597), .C(n25279), 
         .Z(n24915)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam is_jalr_N_1103_bdd_2_lut_3_lut.init = 16'h2020;
    L6MUX21 mux_1323_i2 (.D0(n2066[1]), .D1(n2075[1]), .SD(n2244), .Z(n2089[1]));
    L6MUX21 mux_2209_i2 (.D0(n3657[1]), .D1(n3665[1]), .SD(n3993), .Z(n3675[1]));
    L6MUX21 mux_2209_i3 (.D0(n3657[2]), .D1(n3665[2]), .SD(n3993), .Z(n3675[2]));
    L6MUX21 mux_2209_i4 (.D0(n3657[3]), .D1(n3665[3]), .SD(n3993), .Z(n3675[3]));
    PFUMX mux_1323_i1 (.BLUT(n2066[0]), .ALUT(n2075[0]), .C0(n2244), .Z(n2089[0]));
    LUT4 is_lui_I_0_473_2_lut_rep_645 (.A(is_lui), .B(debug_instr_valid), 
         .Z(n25381)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam is_lui_I_0_473_2_lut_rep_645.init = 16'h8888;
    LUT4 mux_91_i1_3_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(debug_rd_3__N_136[28]), 
         .D(n157), .Z(n234[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam mux_91_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_adj_369 (.A(n20605), .B(n25181), .C(clk_c_enable_54), 
         .Z(clk_c_enable_56)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_adj_369.init = 16'hfefe;
    LUT4 i1_3_lut_adj_370 (.A(n20605), .B(n25181), .C(mem_op[0]), .Z(n21389)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_adj_370.init = 16'hfefe;
    LUT4 i21047_3_lut_4_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(n23319), 
         .D(n25412), .Z(n23322)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i21047_3_lut_4_lut_4_lut.init = 16'h4000;
    L6MUX21 mux_2209_i1 (.D0(n3657[0]), .D1(n3665[0]), .SD(n3993), .Z(n3675[0]));
    LUT4 i1_3_lut_4_lut_adj_371 (.A(n25249), .B(n25195), .C(n26612), .D(n25227), 
         .Z(n22160)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_371.init = 16'h0080;
    PFUMX mux_1544_i17 (.BLUT(n2772[16]), .ALUT(n4516[16]), .C0(n3615), 
          .Z(n2890[16]));
    FD1P3IX pc_offset__i8 (.D(pc_23__N_642[5]), .SP(clk_c_enable_393), .CD(n25424), 
            .CK(clk_c), .Q(\pc[8] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i8.GSR = "DISABLED";
    LUT4 i1_3_lut_adj_372 (.A(is_load), .B(n20805), .C(load_started), 
         .Z(n20605)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_adj_372.init = 16'h7575;
    LUT4 i1_2_lut_rep_647 (.A(is_store), .B(is_load), .Z(n25383)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_rep_647.init = 16'heeee;
    LUT4 debug_instr_valid_N_164_I_0_3_lut_rep_613_4_lut (.A(is_store), .B(is_load), 
         .C(no_write_in_progress), .D(debug_instr_valid), .Z(n25349)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam debug_instr_valid_N_164_I_0_3_lut_rep_613_4_lut.init = 16'h0eff;
    LUT4 mux_1313_i1_4_lut (.A(n2047[0]), .B(n25284), .C(n2242), .D(n25258), 
         .Z(n2075[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam mux_1313_i1_4_lut.init = 16'hca0a;
    LUT4 i11668_3_lut (.A(n25289), .B(n2240), .C(n2236), .Z(n2066[0])) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam i11668_3_lut.init = 16'hc8c8;
    LUT4 i1_3_lut_rep_651 (.A(no_write_in_progress), .B(debug_instr_valid), 
         .C(is_store), .Z(n25387)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_3_lut_rep_651.init = 16'h8080;
    LUT4 i21922_2_lut_4_lut (.A(no_write_in_progress), .B(debug_instr_valid), 
         .C(is_store), .D(n25410), .Z(n23111)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i21922_2_lut_4_lut.init = 16'hff80;
    LUT4 i21726_4_lut (.A(n25182), .B(rst_reg_n), .C(n20952), .D(n21884), 
         .Z(clk_c_enable_93)) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;
    defparam i21726_4_lut.init = 16'h3733;
    LUT4 mux_1522_i3_4_lut (.A(n22964), .B(n25288), .C(n3615), .D(n25209), 
         .Z(n2772[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1522_i3_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_373 (.A(n25177), .B(n8), .C(n25182), .D(n22112), 
         .Z(debug_ret)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_373.init = 16'h0200;
    LUT4 mux_2704_i1_4_lut (.A(addr_out[1]), .B(\imm[1] ), .C(n25411), 
         .D(\pc[1] ), .Z(n4455[0])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(403[26] 407[20])
    defparam mux_2704_i1_4_lut.init = 16'h3aca;
    LUT4 mux_1522_i4_4_lut (.A(n22966), .B(n25287), .C(n3615), .D(n25209), 
         .Z(n2772[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1522_i4_4_lut.init = 16'hca0a;
    PFUMX mux_1544_i5 (.BLUT(n2772[4]), .ALUT(n4516[4]), .C0(n3615), .Z(n2890[4]));
    LUT4 pc_3__bdd_3_lut_22205 (.A(\pc[7] ), .B(\pc[15] ), .C(counter_hi[3]), 
         .Z(n24616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_3__bdd_3_lut_22205.init = 16'hcaca;
    LUT4 i1_2_lut_rep_658 (.A(instr_addr_23__N_49[1]), .B(instr_addr_23__N_49[0]), 
         .Z(n25394)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_rep_658.init = 16'heeee;
    PFUMX mux_1308_i2 (.BLUT(n2034[1]), .ALUT(n2042[1]), .C0(n2240), .Z(n2066[1]));
    PFUMX mux_1517_i8 (.BLUT(n4608[6]), .ALUT(n2414[7]), .C0(n3605), .Z(n2703[7]));
    LUT4 mem_data_from_read_4__bdd_3_lut_22394_then_4_lut (.A(data_txn_len[0]), 
         .B(\qspi_data_buf[12] ), .C(instr_data[12]), .D(n25253), .Z(n25439)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B)) */ ;
    defparam mem_data_from_read_4__bdd_3_lut_22394_then_4_lut.init = 16'he4cc;
    LUT4 i1_4_lut_adj_374 (.A(n25181), .B(n21369), .C(n25179), .D(n22354), 
         .Z(clk_c_enable_110)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;
    defparam i1_4_lut_adj_374.init = 16'h3332;
    LUT4 i21712_4_lut (.A(n25182), .B(n25179), .C(is_ret_de), .D(n7955), 
         .Z(debug_instr_valid_N_167)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21712_4_lut.init = 16'h0001;
    LUT4 i1_3_lut_adj_375 (.A(n20605), .B(n25181), .C(mem_op[1]), .Z(n21388)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_adj_375.init = 16'hfefe;
    LUT4 i30_3_lut_4_lut_3_lut (.A(n26597), .B(n25284), .C(n25281), .Z(n13)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam i30_3_lut_4_lut_3_lut.init = 16'h1818;
    PFUMX mux_1517_i5 (.BLUT(n4608[3]), .ALUT(n2414[4]), .C0(n3605), .Z(n2703[4]));
    LUT4 i21600_3_lut_4_lut (.A(n25265), .B(n26596), .C(n1943), .D(n22056), 
         .Z(n1718[0])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21600_3_lut_4_lut.init = 16'hefe0;
    PFUMX mux_2199_i4 (.BLUT(n21153), .ALUT(n3631[3]), .C0(n3989), .Z(n3657[3]));
    LUT4 i1_4_lut_4_lut_adj_376 (.A(n25284), .B(n25236), .C(n25244), .D(n25222), 
         .Z(is_lui_N_1096)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_376.init = 16'h4000;
    LUT4 i22_4_lut_4_lut (.A(n25284), .B(n26597), .C(n20720), .D(n25247), 
         .Z(n8_adj_2384)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam i22_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i11896_2_lut_3_lut_4_lut (.A(n22), .B(n25158), .C(instr[12]), 
         .D(n3589), .Z(n2627[5])) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i11896_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i11904_4_lut (.A(n25287), .B(n26598), .C(n25267), .D(n25281), 
         .Z(n2736[3])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i11904_4_lut.init = 16'hc088;
    PFUMX mux_2199_i3 (.BLUT(n21152), .ALUT(n3631[2]), .C0(n3989), .Z(n3657[2]));
    LUT4 i21605_3_lut_4_lut_4_lut (.A(n26596), .B(n22044), .C(n1943), 
         .D(instr[4]), .Z(n1718[2])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam i21605_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_40_i4_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_136[31]), 
         .D(data_rs2[3]), .Z(n92[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i4_3_lut_4_lut.init = 16'hf780;
    PFUMX i22176 (.BLUT(n24566), .ALUT(n24565), .C0(n25167), .Z(n24567));
    LUT4 mux_1266_i1_3_lut_rep_705 (.A(n1950[0]), .B(n1970[0]), .C(n25338), 
         .Z(n26597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i1_3_lut_rep_705.init = 16'hcaca;
    LUT4 i21607_3_lut_4_lut_4_lut (.A(n26596), .B(n22068), .C(n1943), 
         .D(n25264), .Z(n1718[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam i21607_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_40_i1_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_136[28]), 
         .D(data_rs2[0]), .Z(n92[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_40_i2_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_136[29]), 
         .D(data_rs2[1]), .Z(n92[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_40_i3_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_136[30]), 
         .D(data_rs2[2]), .Z(n92[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i11905_4_lut (.A(n25278), .B(n26598), .C(n25266), .D(n25281), 
         .Z(n2736[4])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i11905_4_lut.init = 16'hc088;
    LUT4 pc_3__bdd_3_lut_22771 (.A(\pc[3] ), .B(\pc[11] ), .C(counter_hi[3]), 
         .Z(n24617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_3__bdd_3_lut_22771.init = 16'hcaca;
    PFUMX mux_2199_i2 (.BLUT(n21148), .ALUT(n3631[1]), .C0(n3989), .Z(n3657[1]));
    LUT4 mux_2789_i1_3_lut (.A(\instr_addr_23__N_49[22] ), .B(\early_branch_addr[23] ), 
         .C(was_early_branch), .Z(\instr_addr[23] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[25:119])
    defparam mux_2789_i1_3_lut.init = 16'hcaca;
    PFUMX mux_1323_i4 (.BLUT(n21303), .ALUT(n2075[3]), .C0(n2244), .Z(n2089[3]));
    LUT4 i21772_4_lut (.A(n25182), .B(rst_reg_n), .C(n20952), .D(n21970), 
         .Z(clk_c_enable_74)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i21772_4_lut.init = 16'h3337;
    LUT4 i21603_3_lut_4_lut_4_lut (.A(n26596), .B(n22080), .C(n1943), 
         .D(n25267), .Z(n1718[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam i21603_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 i1_4_lut_adj_377 (.A(n25182), .B(n20952), .C(n25336), .D(n21992), 
         .Z(clk_c_enable_91)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(410[18] 430[16])
    defparam i1_4_lut_adj_377.init = 16'h1000;
    LUT4 i11906_4_lut (.A(n25265), .B(n26598), .C(instr[12]), .D(n25281), 
         .Z(n2736[5])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i11906_4_lut.init = 16'hc088;
    LUT4 n26286_bdd_2_lut_4_lut (.A(n1950[0]), .B(n1970[0]), .C(n25338), 
         .D(n26286), .Z(n26287)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam n26286_bdd_2_lut_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_rep_670 (.A(instr_addr_23__N_49[1]), .B(instr_addr_23__N_49[0]), 
         .Z(n25406)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_670.init = 16'h8888;
    LUT4 i11907_4_lut (.A(n25267), .B(n26598), .C(n25265), .D(n25281), 
         .Z(n2736[6])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i11907_4_lut.init = 16'hc088;
    LUT4 i1_2_lut_3_lut_adj_378 (.A(instr_addr_23__N_49[1]), .B(instr_addr_23__N_49[0]), 
         .C(n26612), .Z(n21992)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_378.init = 16'h8080;
    LUT4 mux_1517_i7_4_lut (.A(n2047[0]), .B(n25267), .C(n3605), .D(n25284), 
         .Z(n2703[6])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1517_i7_4_lut.init = 16'hfaca;
    LUT4 i11908_4_lut (.A(n25266), .B(n26598), .C(n25264), .D(n25281), 
         .Z(n2736[7])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i11908_4_lut.init = 16'hc088;
    PFUMX mux_2199_i1 (.BLUT(n21150), .ALUT(n3631[0]), .C0(n3989), .Z(n3657[0]));
    LUT4 n24618_bdd_3_lut (.A(n24618), .B(n24615), .C(n26608), .Z(debug_branch_N_173[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24618_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i9_4_lut (.A(n2813[8]), .B(instr[28]), .C(n3619), .D(n7734), 
         .Z(n2937[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1559_i9_4_lut.init = 16'hca0a;
    LUT4 i21432_3_lut_3_lut (.A(\imm[10] ), .B(n25475), .C(n23011), .Z(n23012)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i21432_3_lut_3_lut.init = 16'he4e4;
    LUT4 i21408_3_lut_3_lut (.A(\imm[10] ), .B(n7775), .C(n4994[2]), .Z(n5029[2])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i21408_3_lut_3_lut.init = 16'he4e4;
    LUT4 counter_2__I_0_i1_1_lut_rep_671 (.A(counter_hi[2]), .Z(n25407)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam counter_2__I_0_i1_1_lut_rep_671.init = 16'h5555;
    LUT4 mux_1505_i4_4_lut (.A(n25267), .B(n21954), .C(n25156), .D(n21212), 
         .Z(n2627[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1505_i4_4_lut.init = 16'hca0a;
    LUT4 i9_4_lut_4_lut (.A(counter_hi[2]), .B(n25408), .C(mie[0]), .D(mie[8]), 
         .Z(n5)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i9_4_lut_4_lut.init = 16'h7340;
    LUT4 i1_2_lut_3_lut_3_lut (.A(counter_hi[2]), .B(counter_hi[4]), .C(counter_hi[3]), 
         .Z(n22798)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 mux_1266_i15_3_lut_rep_706 (.A(n1950[14]), .B(n1970[14]), .C(n25338), 
         .Z(n26598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i15_3_lut_rep_706.init = 16'hcaca;
    LUT4 mux_1505_i7_4_lut (.A(n25289), .B(n21960), .C(n25156), .D(n21212), 
         .Z(n2627[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1505_i7_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_rep_673 (.A(instr_addr_23__N_49[0]), .B(instr_addr_23__N_49[1]), 
         .Z(n25409)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_rep_673.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_379 (.A(n20807), .B(n21322), .C(instr_fetch_running_N_676), 
         .D(instr_fetch_stopped), .Z(clk_c_enable_102)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_379.init = 16'hfffd;
    LUT4 i11492_4_lut (.A(instr_fetch_running_N_674), .B(rst_reg_n), .C(was_early_branch), 
         .D(n25182), .Z(n5438)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam i11492_4_lut.init = 16'hc088;
    LUT4 i11751_4_lut (.A(instr_fetch_running_N_676), .B(n25177), .C(n8), 
         .D(n22030), .Z(instr_fetch_running_N_674)) /* synthesis lut_function=(A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam i11751_4_lut.init = 16'ha2aa;
    LUT4 i1_3_lut_adj_380 (.A(is_jal_de), .B(rst_reg_n), .C(is_ret_de), 
         .Z(n22028)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut_adj_380.init = 16'hc8c8;
    LUT4 mux_1540_i8_3_lut (.A(n2703[7]), .B(n2736[7]), .C(n3613), .Z(n2854[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1540_i8_3_lut.init = 16'hcaca;
    PFUMX mux_1313_i2 (.BLUT(n8768), .ALUT(n2052[1]), .C0(n2242), .Z(n2075[1]));
    PFUMX mux_2203_i4 (.BLUT(n3636[3]), .ALUT(n21376), .C0(n3991), .Z(n3665[3]));
    LUT4 i21878_2_lut_4_lut (.A(n25178), .B(n25175), .C(n22126), .D(rst_reg_n), 
         .Z(clk_c_enable_370)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B (D)))) */ ;
    defparam i21878_2_lut_4_lut.init = 16'h04ff;
    LUT4 i21939_3_lut_4_lut (.A(n3597), .B(n25338), .C(n25167), .D(n3615), 
         .Z(n23271)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21939_3_lut_4_lut.init = 16'hff1f;
    PFUMX mux_2203_i3 (.BLUT(n3636[2]), .ALUT(n21375), .C0(n3991), .Z(n3665[2]));
    LUT4 is_branch_I_0_475_2_lut_rep_675 (.A(is_branch), .B(debug_instr_valid), 
         .Z(n25411)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam is_branch_I_0_475_2_lut_rep_675.init = 16'h8888;
    LUT4 mux_733_i3_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[5] ), 
         .D(addr_out[5]), .Z(n1143[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i2_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[4] ), 
         .D(addr_out[4]), .Z(n1143[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_2704_i2_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[2] ), .D(n25310), .Z(n4455[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_2704_i2_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_2203_i2 (.BLUT(n3636[1]), .ALUT(n21374), .C0(n3991), .Z(n3665[1]));
    LUT4 mux_733_i4_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[6] ), 
         .D(addr_out[6]), .Z(n1143[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i1_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[3] ), 
         .D(addr_out[3]), .Z(n1143[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i5_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[7] ), 
         .D(addr_out[7]), .Z(n1143[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_381 (.A(n2240), .B(n25158), .C(n25288), .D(n4), 
         .Z(n21269)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;
    defparam i1_4_lut_adj_381.init = 16'h20a0;
    LUT4 mux_733_i6_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[8] ), 
         .D(addr_out[8]), .Z(n1143[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i7_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[9] ), 
         .D(addr_out[9]), .Z(n1143[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 i21909_3_lut_4_lut (.A(n25209), .B(n25338), .C(n3615), .D(n3619), 
         .Z(n23155)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21909_3_lut_4_lut.init = 16'h1fff;
    LUT4 mux_733_i8_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[10] ), 
         .D(addr_out[10]), .Z(n1143[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i9_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[11] ), 
         .D(addr_out[11]), .Z(n1143[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i10_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[12] ), .D(addr_out[12]), .Z(n1143[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i10_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_1544_i1 (.BLUT(n21594), .ALUT(n4516[0]), .C0(n3615), .Z(n2890[0]));
    LUT4 mux_733_i11_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[13] ), .D(addr_out[13]), .Z(n1143[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i12_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[14] ), .D(addr_out[14]), .Z(n1143[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i13_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[15] ), .D(addr_out[15]), .Z(n1143[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i13_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_1039_i2 (.BLUT(n1718[1]), .ALUT(n1708[1]), .C0(n1945), .Z(n1729[1]));
    LUT4 mux_733_i14_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[16] ), .D(addr_out[16]), .Z(n1143[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 n20725_bdd_2_lut_22411_4_lut (.A(n25230), .B(n25210), .C(n26598), 
         .D(n25227), .Z(n24956)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam n20725_bdd_2_lut_22411_4_lut.init = 16'h0002;
    LUT4 mux_733_i15_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[17] ), .D(addr_out[17]), .Z(n1143[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_455_4_lut (.A(n25230), .B(n25210), .C(n26598), .D(n25249), 
         .Z(n25191)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_rep_455_4_lut.init = 16'h0200;
    LUT4 mux_733_i16_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[18] ), .D(addr_out[18]), .Z(n1143[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i17_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[19] ), .D(addr_out[19]), .Z(n1143[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i18_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[20] ), .D(addr_out[20]), .Z(n1143[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i19_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[21] ), .D(addr_out[21]), .Z(n1143[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1540_i5_3_lut (.A(n2703[4]), .B(n2736[4]), .C(n3613), .Z(n2854[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1540_i5_3_lut.init = 16'hcaca;
    PFUMX i22525 (.BLUT(n25441), .ALUT(n25442), .C0(counter_hi[2]), .Z(n25443));
    LUT4 mux_733_i20_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[22] ), .D(addr_out[22]), .Z(n1143[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_733_i21_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[23] ), .D(addr_out[23]), .Z(n1143[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_733_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_489_3_lut_4_lut (.A(n25279), .B(n25284), .C(n26597), 
         .D(n26598), .Z(n25225)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_rep_489_3_lut_4_lut.init = 16'h0002;
    PFUMX mux_1039_i3 (.BLUT(n1718[2]), .ALUT(n1708[2]), .C0(n1945), .Z(n1729[2]));
    LUT4 i1_4_lut_adj_382 (.A(n21868), .B(n21864), .C(instr_complete_N_1378), 
         .D(n25349), .Z(\next_instr_write_offset[3] )) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i1_4_lut_adj_382.init = 16'haa6a;
    PFUMX mux_1039_i4 (.BLUT(n1718[3]), .ALUT(n1708[3]), .C0(n1945), .Z(n1729[3]));
    PFUMX mux_2203_i1 (.BLUT(n3636[0]), .ALUT(n3641[0]), .C0(n3991), .Z(n3665[0]));
    PFUMX mux_1039_i1 (.BLUT(n1718[0]), .ALUT(n1708[0]), .C0(n1945), .Z(n1729[0]));
    PFUMX mux_1544_i7 (.BLUT(n22976), .ALUT(n2772[6]), .C0(n23255), .Z(n2890[6]));
    LUT4 i1_2_lut_rep_679 (.A(instr_addr_23__N_49[1]), .B(instr_addr_23__N_49[0]), 
         .Z(n25415)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_rep_679.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_383 (.A(instr_addr_23__N_49[1]), .B(instr_addr_23__N_49[0]), 
         .C(n26612), .Z(n22010)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_3_lut_adj_383.init = 16'hbfbf;
    LUT4 i21931_2_lut_3_lut_4_lut (.A(n22126), .B(n25175), .C(n25281), 
         .D(n25178), .Z(n23089)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i21931_2_lut_3_lut_4_lut.init = 16'hffbf;
    PFUMX mux_55_i2 (.BLUT(n7375), .ALUT(additional_mem_ops_de[1]), .C0(n23089), 
          .Z(n4030[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    PFUMX mux_55_i1 (.BLUT(n6647), .ALUT(additional_mem_ops_de[0]), .C0(n23089), 
          .Z(n4030[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i1_3_lut_rep_461 (.A(is_timer_addr), .B(n20805), .C(data_ready_latch), 
         .Z(n25197)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(258[53:106])
    defparam i1_3_lut_rep_461.init = 16'hfbfb;
    LUT4 i1_2_lut_rep_682 (.A(\instr_len[2] ), .B(\pc[2] ), .Z(n25418)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_2_lut_rep_682.init = 16'h6666;
    LUT4 i1276_3_lut_rep_602_4_lut_4_lut (.A(\instr_len[2] ), .B(\pc[2] ), 
         .C(debug_instr_valid), .D(n25419), .Z(n25338)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C (D))+!B !(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1276_3_lut_rep_602_4_lut_4_lut.init = 16'h9c6c;
    LUT4 i3598_2_lut_rep_683 (.A(\pc[1] ), .B(instr_len[1]), .Z(n25419)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i3598_2_lut_rep_683.init = 16'h8888;
    LUT4 i4439_2_lut_4_lut (.A(is_timer_addr), .B(n20805), .C(data_ready_latch), 
         .D(n25421), .Z(n6638)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(258[53:106])
    defparam i4439_2_lut_4_lut.init = 16'hfb00;
    LUT4 i2_2_lut_rep_627_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), .C(\pc[2] ), 
         .D(\instr_len[2] ), .Z(n25363)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i2_2_lut_rep_627_3_lut_4_lut.init = 16'h8778;
    LUT4 i3596_2_lut_rep_684 (.A(\pc[1] ), .B(instr_len[1]), .Z(n25420)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i3596_2_lut_rep_684.init = 16'h6666;
    LUT4 i20792_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), .C(counter_hi[2]), 
         .D(\next_pc_for_core[5] ), .Z(n23067)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i20792_3_lut_4_lut.init = 16'hf606;
    LUT4 i1_4_lut_4_lut_adj_384 (.A(\pc[1] ), .B(instr_len[1]), .C(debug_instr_valid), 
         .D(instr_addr_23__N_49[0]), .Z(n8154)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_4_lut_4_lut_adj_384.init = 16'h956a;
    LUT4 mux_347_i1_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), .C(debug_ret), 
         .D(return_addr[1]), .Z(n1768[0])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam mux_347_i1_3_lut_4_lut.init = 16'hf606;
    PFUMX mux_1544_i8 (.BLUT(n2772[7]), .ALUT(n4516[7]), .C0(n3615), .Z(n2890[7]));
    LUT4 i1_2_lut_rep_686 (.A(debug_instr_valid), .B(no_write_in_progress), 
         .Z(n25422)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_2_lut_rep_686.init = 16'h8888;
    LUT4 i21762_4_lut (.A(n25182), .B(n20952), .C(n25336), .D(n22022), 
         .Z(clk_c_enable_216)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i21762_4_lut.init = 16'h0010;
    LUT4 i411_2_lut_rep_424_3_lut_4_lut (.A(n22126), .B(n25175), .C(n26612), 
         .D(n25178), .Z(clk_c_enable_69)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i411_2_lut_rep_424_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_3_lut_4_lut_adj_385 (.A(debug_instr_valid), .B(no_write_in_progress), 
         .C(load_done), .D(is_load), .Z(instr_complete_N_1382)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_3_lut_4_lut_adj_385.init = 16'h8000;
    LUT4 mux_1559_i16_3_lut (.A(n2703[12]), .B(n2854[15]), .C(n23220), 
         .Z(n2937[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1559_i16_3_lut.init = 16'hcaca;
    PFUMX mux_1544_i6 (.BLUT(n2772[5]), .ALUT(n4516[5]), .C0(n3615), .Z(n2890[5]));
    PFUMX mux_734_i21 (.BLUT(n1742[20]), .ALUT(n1143[20]), .C0(n25182), 
          .Z(pc_23__N_642[20]));
    LUT4 i18740_3_lut_rep_527 (.A(n25278), .B(n25284), .C(n26598), .Z(n25263)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i18740_3_lut_rep_527.init = 16'hc8c8;
    LUT4 mux_1266_i4_3_lut_rep_528 (.A(n1950[3]), .B(n1970[3]), .C(n25338), 
         .Z(n25264)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i4_3_lut_rep_528.init = 16'hcaca;
    PFUMX mux_734_i20 (.BLUT(n1742[19]), .ALUT(n1143[19]), .C0(n23898), 
          .Z(pc_23__N_642[19]));
    LUT4 i20628_2_lut_4_lut (.A(n1950[3]), .B(n1970[3]), .C(n25338), .D(instr[12]), 
         .Z(n22839)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i20628_2_lut_4_lut.init = 16'hffca;
    LUT4 instr_6__I_0_i6_2_lut_rep_503_4_lut (.A(n1950[3]), .B(n1970[3]), 
         .C(n25338), .D(n25265), .Z(n25239)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam instr_6__I_0_i6_2_lut_rep_503_4_lut.init = 16'hffca;
    LUT4 mux_1559_i15_3_lut (.A(n2703[12]), .B(n2854[14]), .C(n23220), 
         .Z(n2937[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1559_i15_3_lut.init = 16'hcaca;
    PFUMX mux_734_i19 (.BLUT(n1742[18]), .ALUT(n1143[18]), .C0(n23898), 
          .Z(pc_23__N_642[18]));
    LUT4 pc_2__bdd_3_lut_22228 (.A(\pc[6] ), .B(\pc[14] ), .C(counter_hi[3]), 
         .Z(n24660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_2__bdd_3_lut_22228.init = 16'hcaca;
    PFUMX mux_734_i18 (.BLUT(n1742[17]), .ALUT(n1143[17]), .C0(n23898), 
          .Z(pc_23__N_642[17]));
    LUT4 pc_2__bdd_3_lut_22727 (.A(\pc[2] ), .B(\pc[10] ), .C(counter_hi[3]), 
         .Z(n24661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_2__bdd_3_lut_22727.init = 16'hcaca;
    PFUMX mux_734_i17 (.BLUT(n1742[16]), .ALUT(n1143[16]), .C0(n23898), 
          .Z(pc_23__N_642[16]));
    PFUMX mux_734_i16 (.BLUT(n1742[15]), .ALUT(n1143[15]), .C0(n23897), 
          .Z(pc_23__N_642[15]));
    PFUMX mux_734_i15 (.BLUT(n1742[14]), .ALUT(n1143[14]), .C0(n23897), 
          .Z(pc_23__N_642[14]));
    PFUMX mux_734_i14 (.BLUT(n1742[13]), .ALUT(n1143[13]), .C0(n23897), 
          .Z(pc_23__N_642[13]));
    PFUMX mux_734_i13 (.BLUT(n1742[12]), .ALUT(n1143[12]), .C0(n23897), 
          .Z(pc_23__N_642[12]));
    LUT4 n24662_bdd_3_lut (.A(n24662), .B(n24659), .C(n26608), .Z(debug_branch_N_173[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24662_bdd_3_lut.init = 16'hcaca;
    PFUMX mux_734_i12 (.BLUT(n1742[11]), .ALUT(n1143[11]), .C0(n23896), 
          .Z(pc_23__N_642[11]));
    PFUMX mux_734_i11 (.BLUT(n1742[10]), .ALUT(n1143[10]), .C0(n23896), 
          .Z(pc_23__N_642[10]));
    PFUMX mux_734_i10 (.BLUT(n1742[9]), .ALUT(n1143[9]), .C0(n23896), 
          .Z(pc_23__N_642[9]));
    LUT4 i21783_2_lut_4_lut (.A(n1950[3]), .B(n1970[3]), .C(n25338), .D(n25265), 
         .Z(n20820)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i21783_2_lut_4_lut.init = 16'h35ff;
    LUT4 pc_1__bdd_3_lut_22242 (.A(\pc[5] ), .B(\pc[13] ), .C(counter_hi[3]), 
         .Z(n24686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_1__bdd_3_lut_22242.init = 16'hcaca;
    PFUMX mux_734_i9 (.BLUT(n1742[8]), .ALUT(n1143[8]), .C0(n23896), .Z(pc_23__N_642[8]));
    LUT4 i11914_2_lut_4_lut (.A(n1950[3]), .B(n1970[3]), .C(n25338), .D(n25284), 
         .Z(n2414[7])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11914_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_1559_i14_3_lut (.A(n2703[12]), .B(n2854[13]), .C(n23220), 
         .Z(n2937[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1559_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i13_3_lut (.A(n2703[12]), .B(n2854[12]), .C(n23220), 
         .Z(n2937[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1559_i13_3_lut.init = 16'hcaca;
    LUT4 pc_1__bdd_3_lut_22503 (.A(\pc[1] ), .B(\pc[9] ), .C(counter_hi[3]), 
         .Z(n24687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_1__bdd_3_lut_22503.init = 16'hcaca;
    LUT4 instr_6__I_0_127_i6_2_lut_rep_505_4_lut (.A(n1950[3]), .B(n1970[3]), 
         .C(n25338), .D(n25265), .Z(n25241)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam instr_6__I_0_127_i6_2_lut_rep_505_4_lut.init = 16'hcaff;
    PFUMX mux_734_i8 (.BLUT(n1742[7]), .ALUT(n1143[7]), .C0(n23895), .Z(pc_23__N_642[7]));
    LUT4 mux_1266_i3_3_lut_rep_529 (.A(n1950[2]), .B(n1970[2]), .C(n25338), 
         .Z(n25265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i3_3_lut_rep_529.init = 16'hcaca;
    PFUMX mux_734_i7 (.BLUT(n1742[6]), .ALUT(n1143[6]), .C0(n23895), .Z(pc_23__N_642[6]));
    PFUMX mux_734_i6 (.BLUT(n1742[5]), .ALUT(n1143[5]), .C0(n23895), .Z(pc_23__N_642[5]));
    PFUMX i22138 (.BLUT(n24488), .ALUT(n24487), .C0(n3611), .Z(n24489));
    PFUMX i21987 (.BLUT(n24229), .ALUT(n24228), .C0(n3603), .Z(n24230));
    PFUMX mux_734_i5 (.BLUT(n1742[4]), .ALUT(n1143[4]), .C0(n23895), .Z(pc_23__N_642[4]));
    PFUMX mux_734_i4 (.BLUT(n1742[3]), .ALUT(n1143[3]), .C0(n23894), .Z(pc_23__N_642[3]));
    LUT4 mux_1559_i11_4_lut (.A(n2414[9]), .B(instr[30]), .C(n3619), .D(n7734), 
         .Z(n2937[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1559_i11_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_386 (.A(n4030[2]), .B(n4030[1]), .C(n4030[0]), .D(n25178), 
         .Z(additional_mem_ops_2__N_480[2])) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_386.init = 16'ha9aa;
    PFUMX mux_734_i3 (.BLUT(n1742[2]), .ALUT(n1143[2]), .C0(n23894), .Z(pc_23__N_642[2]));
    LUT4 i20833_2_lut_rep_690 (.A(counter_hi[4]), .B(n26610), .Z(n25426)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i20833_2_lut_rep_690.init = 16'h4444;
    LUT4 pc_23__I_0_450_i269_rep_60_3_lut_4_lut (.A(counter_hi[4]), .B(counter_hi[3]), 
         .C(n209_adj_2376), .D(n22941), .Z(n22939)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam pc_23__I_0_450_i269_rep_60_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i11658_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[20] ), 
         .D(\next_pc_for_core[16] ), .Z(n225)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i11658_4_lut_4_lut.init = 16'h5140;
    LUT4 i11659_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[21] ), 
         .D(\next_pc_for_core[17] ), .Z(n226)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i11659_4_lut_4_lut.init = 16'h5140;
    LUT4 next_pc_for_core_23__bdd_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(\next_pc_for_core[19] ), .D(\next_pc_for_core[23] ), .Z(n24264)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam next_pc_for_core_23__bdd_4_lut_4_lut.init = 16'h5410;
    LUT4 c_2__N_1592_1__bdd_4_lut_4_lut (.A(n26610), .B(counter_hi[2]), 
         .C(\pc[21] ), .D(\pc[17] ), .Z(n24685)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam c_2__N_1592_1__bdd_4_lut_4_lut.init = 16'h5140;
    LUT4 c_2__N_1592_1__bdd_4_lut_22227_4_lut (.A(n26610), .B(counter_hi[2]), 
         .C(\pc[23] ), .D(\pc[19] ), .Z(n24615)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam c_2__N_1592_1__bdd_4_lut_22227_4_lut.init = 16'h5140;
    PFUMX mux_734_i2 (.BLUT(n1742[1]), .ALUT(n1143[1]), .C0(n23894), .Z(pc_23__N_642[1]));
    LUT4 i11624_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\pc[20] ), 
         .D(\pc[16] ), .Z(n225_adj_2385)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i11624_4_lut_4_lut.init = 16'h5140;
    LUT4 c_2__N_1592_1__bdd_4_lut_22240_4_lut (.A(n26610), .B(counter_hi[2]), 
         .C(\pc[22] ), .D(\pc[18] ), .Z(n24659)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam c_2__N_1592_1__bdd_4_lut_22240_4_lut.init = 16'h5140;
    LUT4 n24688_bdd_3_lut (.A(n24688), .B(n24685), .C(n26608), .Z(debug_branch_N_173[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24688_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i10_4_lut (.A(n24489), .B(instr[29]), .C(n3619), .D(n7734), 
         .Z(n2937[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1559_i10_4_lut.init = 16'hca0a;
    LUT4 instr_6__bdd_2_lut_21986_2_lut_4_lut (.A(n1950[2]), .B(n1970[2]), 
         .C(n25338), .D(n25279), .Z(n24228)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam instr_6__bdd_2_lut_21986_2_lut_4_lut.init = 16'h00ca;
    PFUMX mux_734_i1 (.BLUT(n1742[0]), .ALUT(n1143[0]), .C0(n23894), .Z(pc_23__N_642[0]));
    LUT4 i18680_2_lut_rep_492_4_lut (.A(n1950[2]), .B(n1970[2]), .C(n25338), 
         .D(instr[4]), .Z(n25228)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i18680_2_lut_rep_492_4_lut.init = 16'hca00;
    LUT4 i20626_2_lut_rep_525_4_lut (.A(n1950[2]), .B(n1970[2]), .C(n25338), 
         .D(instr[4]), .Z(n25261)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i20626_2_lut_rep_525_4_lut.init = 16'hffca;
    LUT4 mux_1266_i7_3_lut_rep_530 (.A(n1950[6]), .B(n1970[6]), .C(n25338), 
         .Z(n25266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i7_3_lut_rep_530.init = 16'hcaca;
    LUT4 instr_6__I_0_126_i7_2_lut_rep_526_4_lut (.A(n1950[6]), .B(n1970[6]), 
         .C(n25338), .D(n25267), .Z(n25262)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam instr_6__I_0_126_i7_2_lut_rep_526_4_lut.init = 16'hffca;
    LUT4 i11615_2_lut_rep_507_4_lut (.A(n1950[6]), .B(n1970[6]), .C(n25338), 
         .D(n25267), .Z(n25243)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11615_2_lut_rep_507_4_lut.init = 16'hca00;
    LUT4 i11928_2_lut_2_lut_4_lut (.A(n1950[6]), .B(n1970[6]), .C(n25338), 
         .D(n26598), .Z(n4608[6])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11928_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 instr_6__bdd_2_lut_4_lut (.A(n1950[6]), .B(n1970[6]), .C(n25338), 
         .D(n25287), .Z(n24229)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam instr_6__bdd_2_lut_4_lut.init = 16'h00ca;
    LUT4 n24567_bdd_3_lut_4_lut (.A(n25209), .B(n25290), .C(n3615), .D(n24567), 
         .Z(n24568)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n24567_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i12171_3_lut_4_lut (.A(n25221), .B(n26598), .C(n25284), .D(n25279), 
         .Z(n29)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (D)))) */ ;
    defparam i12171_3_lut_4_lut.init = 16'h001f;
    LUT4 instr_6__I_0_150_i7_2_lut_rep_498_4_lut (.A(n1950[6]), .B(n1970[6]), 
         .C(n25338), .D(n25267), .Z(n25234)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam instr_6__I_0_150_i7_2_lut_rep_498_4_lut.init = 16'hcaff;
    LUT4 i11911_2_lut_4_lut (.A(n1950[6]), .B(n1970[6]), .C(n25338), .D(n25284), 
         .Z(n2414[4])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11911_2_lut_4_lut.init = 16'hffca;
    LUT4 i3527_2_lut_rep_693 (.A(rs2[0]), .B(mem_op_increment_reg), .Z(n25429)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i3527_2_lut_rep_693.init = 16'h8888;
    LUT4 mux_1266_i6_3_lut_rep_531 (.A(n1950[5]), .B(n1970[5]), .C(n25338), 
         .Z(n25267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i6_3_lut_rep_531.init = 16'hcaca;
    LUT4 mux_1013_i11_rep_98_3_lut (.A(n1649[10]), .B(instr[31]), .C(n25209), 
         .Z(n22977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i11_rep_98_3_lut.init = 16'hcaca;
    LUT4 i3535_2_lut_rep_632_3_lut (.A(rs2[0]), .B(mem_op_increment_reg), 
         .C(rs2[1]), .Z(n25368)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i3535_2_lut_rep_632_3_lut.init = 16'h8080;
    LUT4 mux_1013_i8_rep_84_3_lut (.A(n22972), .B(instr[31]), .C(n25209), 
         .Z(n22963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i8_rep_84_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_387 (.A(n1950[5]), .B(n1970[5]), .C(n25338), 
         .D(instr[4]), .Z(n20650)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_4_lut_adj_387.init = 16'h00ca;
    LUT4 i3542_2_lut_3_lut_4_lut (.A(rs2[0]), .B(mem_op_increment_reg), 
         .C(rs2[2]), .D(rs2[1]), .Z(n5570)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i3542_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_1013_i7_rep_82_3_lut (.A(n22974), .B(instr[31]), .C(n25209), 
         .Z(n22961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i7_rep_82_3_lut.init = 16'hcaca;
    LUT4 is_system_I_0_481_2_lut_rep_694 (.A(is_system), .B(debug_instr_valid), 
         .Z(n25430)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam is_system_I_0_481_2_lut_rep_694.init = 16'h8888;
    LUT4 is_csr_I_0_573_2_lut_rep_607_4_lut_3_lut_4_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[1]), .D(alu_op[0]), .Z(n25343)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam is_csr_I_0_573_2_lut_rep_607_4_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 mux_1013_i6_rep_74_3_lut (.A(n22968), .B(instr[31]), .C(n25209), 
         .Z(n22953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i6_rep_74_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_605_2_lut_3_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[1]), .Z(n25341)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_605_2_lut_3_lut.init = 16'h8080;
    L6MUX21 i21151 (.D0(n23424), .D1(n23425), .SD(n26608), .Z(debug_rd_3__N_136[28]));
    LUT4 i1_2_lut_rep_583_3_lut_3_lut_4_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[1]), .D(alu_op[0]), .Z(n25319)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_583_3_lut_3_lut_4_lut.init = 16'h0080;
    L6MUX21 i21158 (.D0(n23431), .D1(n23432), .SD(n26608), .Z(debug_rd_3__N_136[29]));
    L6MUX21 i21165 (.D0(n23438), .D1(n23439), .SD(n26608), .Z(debug_rd_3__N_136[30]));
    L6MUX21 i21172 (.D0(n23445), .D1(n23446), .SD(n26608), .Z(debug_rd_3__N_136[31]));
    LUT4 i1_2_lut_rep_565_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut (.A(is_system), 
         .B(debug_instr_valid), .C(alu_op[1]), .D(alu_op[0]), .Z(n25301)) /* synthesis lut_function=(!(((C (D)+!C !(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_565_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h0880;
    LUT4 i18726_2_lut_3_lut_4_lut_2_lut_3_lut_3_lut_4_lut_3_lut_4_lut (.A(is_system), 
         .B(debug_instr_valid), .C(alu_op[1]), .D(alu_op[0]), .Z(n25369)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i18726_2_lut_3_lut_4_lut_2_lut_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h8880;
    LUT4 i12164_2_lut_3_lut_4_lut (.A(n22126), .B(n25175), .C(n26612), 
         .D(n25178), .Z(clk_c_enable_312)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i12164_2_lut_3_lut_4_lut.init = 16'hf040;
    LUT4 mux_1013_i5_rep_76_3_lut (.A(n22970), .B(instr[31]), .C(n25209), 
         .Z(n22955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i5_rep_76_3_lut.init = 16'hcaca;
    PFUMX pc_23__I_0_450_i209 (.BLUT(n149_adj_2377), .ALUT(n225_adj_2385), 
          .C0(n26608), .Z(n209_adj_2376)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i11677_2_lut (.A(n24230), .B(n3611), .Z(n2813[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i11677_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_696 (.A(qv_data_write_n[1]), .B(qv_data_write_n[0]), 
         .Z(n25432)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam i1_2_lut_rep_696.init = 16'h8888;
    LUT4 i1_2_lut_rep_564_3_lut (.A(qv_data_write_n[1]), .B(qv_data_write_n[0]), 
         .C(is_timer_addr), .Z(n25300)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam i1_2_lut_rep_564_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_546_3_lut_4_lut (.A(qv_data_write_n[1]), .B(qv_data_write_n[0]), 
         .C(addr[2]), .D(is_timer_addr), .Z(n25282)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam i1_2_lut_rep_546_3_lut_4_lut.init = 16'h7000;
    LUT4 i1_3_lut_4_lut_adj_388 (.A(qv_data_write_n[1]), .B(qv_data_write_n[0]), 
         .C(data_ready_sync), .D(n20805), .Z(n66)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam i1_3_lut_4_lut_adj_388.init = 16'hf8ff;
    LUT4 i1_2_lut_rep_533_3_lut_4_lut (.A(qv_data_write_n[1]), .B(qv_data_write_n[0]), 
         .C(addr[2]), .D(is_timer_addr), .Z(n25269)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam i1_2_lut_rep_533_3_lut_4_lut.init = 16'h0700;
    LUT4 i3926_2_lut_3_lut_4_lut_4_lut (.A(n25372), .B(cycle_count_wide[0]), 
         .C(cycle_count_wide[1]), .D(cy), .Z(increment_result_3__N_1642[1])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i3926_2_lut_3_lut_4_lut_4_lut.init = 16'h3cb4;
    LUT4 mux_2756_i12_3_lut (.A(instr[12]), .B(n25265), .C(n26598), .Z(n4608[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2756_i12_3_lut.init = 16'hcaca;
    LUT4 mux_2756_i13_3_lut (.A(instr[12]), .B(n25264), .C(n26598), .Z(n4608[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2756_i13_3_lut.init = 16'hcaca;
    LUT4 mux_2756_i14_3_lut (.A(instr[12]), .B(instr[4]), .C(n26598), 
         .Z(n4608[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2756_i14_3_lut.init = 16'hcaca;
    LUT4 mux_2756_i15_3_lut (.A(instr[12]), .B(n25267), .C(n26598), .Z(n4608[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2756_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1003_i2_rep_115_3_lut (.A(n2[1]), .B(n7[1]), .C(n1949), .Z(n22994)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i2_rep_115_3_lut.init = 16'hcaca;
    FD1S3IX counter_hi_3136__i3_rep_710 (.D(n17_adj_2394[1]), .CK(clk_c), 
            .CD(n25424), .Q(n26610));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3136__i3_rep_710.GSR = "DISABLED";
    LUT4 i3946_2_lut_4_lut_4_lut (.A(n25372), .B(instrret_count[0]), .C(instr_retired), 
         .D(cy_adj_2386), .Z(increment_result_3__N_1656[0])) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i3946_2_lut_4_lut_4_lut.init = 16'h369c;
    PFUMX i20794 (.BLUT(n23068), .ALUT(n226), .C0(counter_hi[4]), .Z(n23069));
    LUT4 mem_data_from_read_4__bdd_3_lut_22394_else_4_lut (.A(data_txn_len[0]), 
         .B(n25253), .C(instr_data[8]), .D(\qspi_data_buf[8] ), .Z(n25438)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mem_data_from_read_4__bdd_3_lut_22394_else_4_lut.init = 16'hf780;
    LUT4 i3948_2_lut_rep_558_4_lut_4_lut (.A(n25372), .B(instrret_count[0]), 
         .C(instr_retired), .D(cy_adj_2386), .Z(n25294)) /* synthesis lut_function=(A (B (D))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i3948_2_lut_rep_558_4_lut_4_lut.init = 16'hc840;
    LUT4 i1_3_lut_4_lut_adj_389 (.A(n25304), .B(n25161), .C(data_txn_len[1]), 
         .D(instr_active), .Z(\txn_len[1] )) /* synthesis lut_function=(!(A ((D)+!C)+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(435[34:115])
    defparam i1_3_lut_4_lut_adj_389.init = 16'h00b0;
    LUT4 mux_1266_i12_3_lut_rep_542 (.A(n1950[11]), .B(n1970[11]), .C(n25338), 
         .Z(n25278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i12_3_lut_rep_542.init = 16'hcaca;
    LUT4 mux_1003_i3_rep_113_3_lut (.A(n2[2]), .B(n7[2]), .C(n1949), .Z(n22992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i3_rep_113_3_lut.init = 16'hcaca;
    LUT4 i11926_2_lut_2_lut_4_lut (.A(n1950[11]), .B(n1970[11]), .C(n25338), 
         .D(n26598), .Z(n4608[3])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11926_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 i21759_2_lut_rep_520_4_lut (.A(n1950[11]), .B(n1970[11]), .C(n25338), 
         .D(n25287), .Z(n25256)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i21759_2_lut_rep_520_4_lut.init = 16'h35ff;
    LUT4 mux_1266_i14_3_lut_rep_543 (.A(n1950[13]), .B(n1970[13]), .C(n25338), 
         .Z(n25279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i14_3_lut_rep_543.init = 16'hcaca;
    PFUMX i22118 (.BLUT(n24451), .ALUT(n24449), .C0(n3615), .Z(n24452));
    LUT4 i21946_2_lut_rep_416 (.A(n3613), .B(n3605), .Z(n25152)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21946_2_lut_rep_416.init = 16'hbbbb;
    LUT4 mux_1517_i14_3_lut_4_lut (.A(instr[12]), .B(n25229), .C(n3613), 
         .D(n2414[9]), .Z(n2703[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1517_i14_3_lut_4_lut.init = 16'h8f80;
    LUT4 gnd_bdd_2_lut_22402_2_lut_4_lut (.A(n1950[13]), .B(n1970[13]), 
         .C(n25338), .D(n24913), .Z(n24914)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam gnd_bdd_2_lut_22402_2_lut_4_lut.init = 16'h3500;
    LUT4 mux_1517_i17_3_lut_4_lut (.A(instr[12]), .B(n25229), .C(n3613), 
         .D(n2414[16]), .Z(n2703[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1517_i17_3_lut_4_lut.init = 16'h8f80;
    LUT4 i3873_2_lut_rep_482_3_lut_4_lut_4_lut (.A(n25372), .B(alu_b_in[0]), 
         .C(n25352), .D(cy_adj_2387), .Z(n25218)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i3873_2_lut_rep_482_3_lut_4_lut_4_lut.init = 16'h3810;
    LUT4 mux_1517_i10_3_lut_4_lut (.A(instr[12]), .B(n25229), .C(n3613), 
         .D(n2047[3]), .Z(n2703[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1517_i10_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_2_lut_rep_495_4_lut (.A(n1950[13]), .B(n1970[13]), .C(n25338), 
         .D(n26598), .Z(n25231)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_2_lut_rep_495_4_lut.init = 16'h3500;
    LUT4 cy_I_0_3_lut_rep_569_4_lut_4_lut (.A(n25372), .B(cy_adj_2388), 
         .C(time_pulse_r), .D(n8527), .Z(n25305)) /* synthesis lut_function=(A (B)+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam cy_I_0_3_lut_rep_569_4_lut_4_lut.init = 16'hd8dd;
    LUT4 mux_1007_i3_3_lut (.A(n9[2]), .B(n14[2]), .C(n1969), .Z(n1649[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i3_3_lut.init = 16'hcaca;
    LUT4 equal_25_i3_2_lut_4_lut (.A(n1950[13]), .B(n1970[13]), .C(n25338), 
         .D(instr[12]), .Z(n3)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam equal_25_i3_2_lut_4_lut.init = 16'hcaff;
    L6MUX21 shift_right_317_i272 (.D0(n212), .D1(n8761), .SD(counter_hi[4]), 
            .Z(debug_branch_N_571[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    PFUMX next_pc_for_core_23__I_0_i209 (.BLUT(n149), .ALUT(n225), .C0(counter_hi[4]), 
          .Z(n209)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i1_2_lut_rep_523_4_lut (.A(n1950[13]), .B(n1970[13]), .C(n25338), 
         .D(n25284), .Z(n25259)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_523_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_494_4_lut (.A(n1950[13]), .B(n1970[13]), .C(n25338), 
         .D(n25284), .Z(n25230)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_494_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_rep_500_4_lut (.A(n1950[13]), .B(n1970[13]), .C(n25338), 
         .D(n26598), .Z(n25236)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_500_4_lut.init = 16'hca00;
    LUT4 mux_1517_i9_3_lut_4_lut (.A(instr[12]), .B(n25229), .C(n3613), 
         .D(n2047[2]), .Z(n2703[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1517_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_4_lut_adj_390 (.A(addr_out[3]), .B(n25310), .C(addr_offset[3]), 
         .D(addr_offset[2]), .Z(n21499)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(266[43:70])
    defparam i1_4_lut_adj_390.init = 16'h965a;
    LUT4 n2784_bdd_3_lut_22101_4_lut (.A(instr[31]), .B(n25258), .C(n25167), 
         .D(n24422), .Z(n24423)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n2784_bdd_3_lut_22101_4_lut.init = 16'hf808;
    LUT4 i1_4_lut_4_lut_adj_391 (.A(n25178), .B(n25175), .C(n22290), .D(n3619), 
         .Z(n21860)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_4_lut_4_lut_adj_391.init = 16'hff40;
    LUT4 i1_2_lut_rep_511_4_lut (.A(n1950[13]), .B(n1970[13]), .C(n25338), 
         .D(n26598), .Z(n25247)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_511_4_lut.init = 16'hffca;
    LUT4 mux_1522_i13_3_lut_4_lut (.A(instr[31]), .B(n25258), .C(n25167), 
         .D(n4548[5]), .Z(n2772[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1522_i13_3_lut_4_lut.init = 16'hf808;
    PFUMX shift_right_317_i212 (.BLUT(n23057), .ALUT(n8735), .C0(counter_hi[3]), 
          .Z(n212)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 mux_1522_i16_3_lut_4_lut (.A(instr[31]), .B(n25258), .C(n25167), 
         .D(n4548[8]), .Z(n2772[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1522_i16_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_1522_i14_3_lut_4_lut (.A(instr[31]), .B(n25258), .C(n25167), 
         .D(n4548[6]), .Z(n2772[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1522_i14_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_1522_i15_3_lut_4_lut (.A(instr[31]), .B(n25258), .C(n25167), 
         .D(n4548[7]), .Z(n2772[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1522_i15_3_lut_4_lut.init = 16'hf808;
    LUT4 n2784_bdd_3_lut_22121_4_lut (.A(instr[31]), .B(n25258), .C(n25167), 
         .D(n24450), .Z(n24451)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n2784_bdd_3_lut_22121_4_lut.init = 16'hf808;
    PFUMX i21149 (.BLUT(n23420), .ALUT(n23421), .C0(counter_hi[3]), .Z(n23424));
    LUT4 i21715_2_lut_4_lut (.A(n1950[13]), .B(n1970[13]), .C(n25338), 
         .D(n26597), .Z(n13701)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i21715_2_lut_4_lut.init = 16'h0035;
    LUT4 i2_2_lut_rep_502_4_lut (.A(n1950[13]), .B(n1970[13]), .C(n25338), 
         .D(n26597), .Z(n25238)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i2_2_lut_rep_502_4_lut.init = 16'h00ca;
    LUT4 i1_3_lut_4_lut_adj_392 (.A(n25304), .B(n25161), .C(n25403), .D(\addr_in[23] ), 
         .Z(spi_ram_b_select_N_2044)) /* synthesis lut_function=(A (C+!(D))+!A (B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(435[34:115])
    defparam i1_3_lut_4_lut_adj_392.init = 16'hf4ff;
    LUT4 i11817_2_lut_4_lut (.A(n1950[14]), .B(n1970[14]), .C(n25338), 
         .D(n25287), .Z(n2047[3])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11817_2_lut_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_rep_509_4_lut (.A(n1950[14]), .B(n1970[14]), .C(n25338), 
         .D(n25284), .Z(n25245)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_509_4_lut.init = 16'hca00;
    LUT4 i11586_2_lut_rep_501_4_lut (.A(n1950[14]), .B(n1970[14]), .C(n25338), 
         .D(n25284), .Z(n25237)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11586_2_lut_rep_501_4_lut.init = 16'hffca;
    LUT4 i21722_2_lut_rep_493_4_lut (.A(n1950[14]), .B(n1970[14]), .C(n25338), 
         .D(n25281), .Z(n25229)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i21722_2_lut_rep_493_4_lut.init = 16'h00ca;
    LUT4 i11816_2_lut_4_lut (.A(n1950[14]), .B(n1970[14]), .C(n25338), 
         .D(n25288), .Z(n2047[2])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11816_2_lut_4_lut.init = 16'h3500;
    LUT4 n2784_bdd_3_lut_22117_4_lut (.A(instr[31]), .B(n25258), .C(n25167), 
         .D(n24429), .Z(n24430)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n2784_bdd_3_lut_22117_4_lut.init = 16'hf808;
    LUT4 additional_mem_ops_2__N_863_0__bdd_2_lut_4_lut (.A(n1950[14]), .B(n1970[14]), 
         .C(n25338), .D(n25189), .Z(n24894)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam additional_mem_ops_2__N_863_0__bdd_2_lut_4_lut.init = 16'h00ca;
    LUT4 i11534_2_lut_4_lut (.A(n1950[14]), .B(n1970[14]), .C(n25338), 
         .D(n25289), .Z(n2047[0])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11534_2_lut_4_lut.init = 16'h3500;
    LUT4 mux_1266_i2_3_lut_rep_545 (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .Z(n25281)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i2_3_lut_rep_545.init = 16'hcaca;
    LUT4 mux_2750_i10_3_lut_4_lut (.A(instr[31]), .B(n25258), .C(n25167), 
         .D(n22990), .Z(n4548[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2750_i10_3_lut_4_lut.init = 16'hf808;
    LUT4 i11517_1_lut_rep_483_2_lut_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n26597), .Z(n25219)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11517_1_lut_rep_483_2_lut_4_lut.init = 16'h35ff;
    LUT4 mux_1007_i12_3_lut (.A(n9[11]), .B(n14[11]), .C(n1969), .Z(n1649[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i12_3_lut.init = 16'hcaca;
    LUT4 i21892_2_lut_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), .D(n26597), 
         .Z(n23379)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i21892_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_3_lut_adj_393 (.A(additional_mem_ops[1]), .B(additional_mem_ops[0]), 
         .C(additional_mem_ops[2]), .Z(any_additional_mem_ops)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(137[35:63])
    defparam i1_3_lut_adj_393.init = 16'hfefe;
    LUT4 i5352_4_lut_4_lut (.A(n25178), .B(n22008), .C(n25214), .D(instr[12]), 
         .Z(n2703[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam i5352_4_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_4_lut_adj_394 (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n25284), .Z(n22384)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_4_lut_adj_394.init = 16'hca00;
    LUT4 mux_2749_i21_3_lut_4_lut (.A(instr[31]), .B(n25258), .C(n3619), 
         .D(n2937[17]), .Z(n4516[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2749_i21_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2750_i5_4_lut_4_lut (.A(instr[31]), .B(n25258), .C(n25209), 
         .D(n3615), .Z(n4548[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2750_i5_4_lut_4_lut.init = 16'ha088;
    LUT4 i21960_2_lut_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), .D(n25284), 
         .Z(n23166)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i21960_2_lut_4_lut.init = 16'hcaff;
    LUT4 i1_2_lut_rep_513_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n26597), .Z(n25249)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_513_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_522_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n26597), .Z(n25258)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_522_4_lut.init = 16'hca00;
    LUT4 i11531_2_lut_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), .D(n25289), 
         .Z(n3636[0])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11531_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_rep_508_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n26597), .Z(n25244)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_508_4_lut.init = 16'h3500;
    LUT4 i1_3_lut_4_lut_adj_395 (.A(n25258), .B(n26612), .C(n20820), .D(n25239), 
         .Z(n21910)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_395.init = 16'h0888;
    LUT4 i166_2_lut_rep_512_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n26597), .Z(n25248)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i166_2_lut_rep_512_4_lut.init = 16'h3500;
    LUT4 gnd_bdd_2_lut_22407_2_lut_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n24941), .Z(n24942)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam gnd_bdd_2_lut_22407_2_lut_4_lut.init = 16'h3500;
    PFUMX i21150 (.BLUT(n23422), .ALUT(n23423), .C0(counter_hi[3]), .Z(n23425));
    LUT4 i11631_2_lut_2_lut_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n25290), .Z(n3636[1])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11631_2_lut_2_lut_4_lut.init = 16'h3500;
    LUT4 i11629_2_lut_2_lut_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n25287), .Z(n3636[3])) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11629_2_lut_2_lut_4_lut.init = 16'hff35;
    LUT4 i11630_2_lut_2_lut_4_lut (.A(n1950[1]), .B(n1970[1]), .C(n25338), 
         .D(n25288), .Z(n3636[2])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11630_2_lut_2_lut_4_lut.init = 16'h3500;
    LUT4 i16394_2_lut (.A(counter_hi[3]), .B(counter_hi[2]), .Z(n17_adj_2394[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i16394_2_lut.init = 16'h6666;
    LUT4 mux_1003_i12_3_lut (.A(n2[11]), .B(n7[11]), .C(n1949), .Z(n1629[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i12_3_lut.init = 16'hcaca;
    LUT4 mtimecmp_5__I_0_3_lut_4_lut (.A(addr[2]), .B(n25300), .C(data_out_slice[1]), 
         .D(mtimecmp[5]), .Z(mtimecmp_1__N_1672)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mtimecmp_5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 mtimecmp_4__I_0_3_lut_4_lut (.A(addr[2]), .B(n25300), .C(data_out_slice[0]), 
         .D(mtimecmp[4]), .Z(mtimecmp_0__N_1674)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mtimecmp_4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 mtimecmp_6__I_0_3_lut_4_lut (.A(addr[2]), .B(n25300), .C(data_out_slice[2]), 
         .D(mtimecmp[6]), .Z(mtimecmp_2__N_1670)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mtimecmp_6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_519_4_lut (.A(n1950[0]), .B(n1970[0]), .C(n25338), 
         .D(n25284), .Z(n25255)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_519_4_lut.init = 16'hca00;
    LUT4 i1_2_lut_rep_521_4_lut (.A(n1950[0]), .B(n1970[0]), .C(n25338), 
         .D(n25284), .Z(n25257)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_rep_521_4_lut.init = 16'h3500;
    LUT4 i21926_2_lut (.A(n26608), .B(n26610), .Z(n23319)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i21926_2_lut.init = 16'heeee;
    PFUMX i21156 (.BLUT(n23427), .ALUT(n23428), .C0(counter_hi[3]), .Z(n23431));
    LUT4 i21733_2_lut_rep_496_4_lut (.A(n1950[0]), .B(n1970[0]), .C(n25338), 
         .D(n25284), .Z(n25232)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i21733_2_lut_rep_496_4_lut.init = 16'h0035;
    LUT4 debug_branch_I_23_i4_3_lut (.A(debug_branch_N_571[31]), .B(timer_data[3]), 
         .C(is_timer_addr), .Z(debug_branch_N_181[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_23_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1266_i16_3_lut_rep_548 (.A(n1950[15]), .B(n1970[15]), .C(n25338), 
         .Z(n25284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i16_3_lut_rep_548.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_396 (.A(n1950[15]), .B(n1970[15]), .C(n25338), 
         .D(rst_reg_n), .Z(n21998)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_4_lut_adj_396.init = 16'hca00;
    L6MUX21 i21128 (.D0(n23399), .D1(n23400), .SD(n26610), .Z(n23403));
    LUT4 i43_3_lut_4_lut (.A(n25232), .B(n25247), .C(n25281), .D(n23), 
         .Z(n26_adj_2389)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam i43_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_1266_i11_3_lut_rep_551 (.A(n1950[10]), .B(n1970[10]), .C(n25338), 
         .Z(n25287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i11_3_lut_rep_551.init = 16'hcaca;
    LUT4 i11871_2_lut_2_lut_4_lut (.A(n1950[10]), .B(n1970[10]), .C(n25338), 
         .D(n25162), .Z(n3631[3])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11871_2_lut_2_lut_4_lut.init = 16'h00ca;
    PFUMX i54 (.BLUT(n37), .ALUT(n32), .C0(n23166), .Z(n35));
    PFUMX i22102 (.BLUT(n24430), .ALUT(n24427), .C0(n3615), .Z(n24431));
    LUT4 i1_4_lut_adj_397 (.A(was_early_branch), .B(n25144), .C(n8154), 
         .D(n25258), .Z(n7955)) /* synthesis lut_function=(A+(B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(156[34] 157[124])
    defparam i1_4_lut_adj_397.init = 16'heeae;
    LUT4 mux_1266_i10_3_lut_rep_552 (.A(n1950[9]), .B(n1970[9]), .C(n25338), 
         .Z(n25288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i10_3_lut_rep_552.init = 16'hcaca;
    LUT4 i11870_2_lut_2_lut_4_lut (.A(n1950[9]), .B(n1970[9]), .C(n25338), 
         .D(n25162), .Z(n3631[2])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11870_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_1266_i8_3_lut_rep_553 (.A(n1950[7]), .B(n1970[7]), .C(n25338), 
         .Z(n25289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i8_3_lut_rep_553.init = 16'hcaca;
    LUT4 i11573_2_lut_4_lut (.A(n1950[7]), .B(n1970[7]), .C(n25338), .D(n25162), 
         .Z(n3631[0])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11573_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_398 (.A(n1950[7]), .B(n1970[7]), .C(n25338), 
         .D(n25290), .Z(n22398)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i1_2_lut_4_lut_adj_398.init = 16'h00ca;
    PFUMX i22959 (.BLUT(n26288), .ALUT(n26287), .C0(n23900), .Z(n26289));
    LUT4 mux_1266_i9_3_lut_rep_554 (.A(n1950[8]), .B(n1970[8]), .C(n25338), 
         .Z(n25290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1266_i9_3_lut_rep_554.init = 16'hcaca;
    LUT4 i11877_2_lut_4_lut (.A(n1950[8]), .B(n1970[8]), .C(n25338), .D(n2236), 
         .Z(n2042[1])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11877_2_lut_4_lut.init = 16'hffca;
    PFUMX i21157 (.BLUT(n23429), .ALUT(n23430), .C0(counter_hi[3]), .Z(n23432));
    LUT4 i11869_2_lut_2_lut_4_lut (.A(n1950[8]), .B(n1970[8]), .C(n25338), 
         .D(n25162), .Z(n3631[1])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam i11869_2_lut_2_lut_4_lut.init = 16'h00ca;
    PFUMX i21163 (.BLUT(n23434), .ALUT(n23435), .C0(counter_hi[3]), .Z(n23438));
    PFUMX i42 (.BLUT(n10_adj_2390), .ALUT(n29), .C0(n26597), .Z(n23));
    LUT4 i1_4_lut_adj_399 (.A(no_write_in_progress), .B(data_ready_core), 
         .C(debug_instr_valid), .D(is_load), .Z(debug_rd_3__N_1306)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_4_lut_adj_399.init = 16'h8000;
    LUT4 i1_3_lut_adj_400 (.A(n7955), .B(n26598), .C(n26612), .Z(n21898)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_400.init = 16'h4040;
    PFUMX i21164 (.BLUT(n23436), .ALUT(n23437), .C0(counter_hi[3]), .Z(n23439));
    LUT4 i1_4_lut_adj_401 (.A(instr[12]), .B(n26612), .C(n25287), .D(n25279), 
         .Z(n22178)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_401.init = 16'hc088;
    PFUMX i21170 (.BLUT(n23441), .ALUT(n23442), .C0(counter_hi[3]), .Z(n23445));
    LUT4 i20665_4_lut (.A(n25169), .B(addr_offset[3]), .C(n25178), .D(addr_offset[2]), 
         .Z(n22878)) /* synthesis lut_function=(!((B (C (D))+!B !(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i20665_4_lut.init = 16'h2888;
    PFUMX i21171 (.BLUT(n23443), .ALUT(n23444), .C0(counter_hi[3]), .Z(n23446));
    LUT4 i1_4_lut_adj_402 (.A(n25266), .B(rst_reg_n), .C(n25278), .D(n25279), 
         .Z(n22238)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_402.init = 16'hc088;
    PFUMX i20764 (.BLUT(n23037), .ALUT(n23038), .C0(counter_hi[2]), .Z(n23039));
    LUT4 i20661_2_lut_3_lut_4_lut (.A(instr_addr_23__N_49[1]), .B(n25311), 
         .C(n1), .D(\pc[2] ), .Z(n22873)) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i20661_2_lut_3_lut_4_lut.init = 16'hf9f6;
    LUT4 i1_3_lut_adj_403 (.A(n25279), .B(instr[4]), .C(rst_reg_n), .Z(n22132)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_403.init = 16'h4040;
    LUT4 mux_346_i2_3_lut_4_lut (.A(instr_addr_23__N_49[1]), .B(n25311), 
         .C(debug_ret), .D(return_addr[2]), .Z(n1764[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam mux_346_i2_3_lut_4_lut.init = 16'hf606;
    PFUMX i22098 (.BLUT(n24423), .ALUT(n24420), .C0(n3615), .Z(n24424));
    L6MUX21 i22509 (.D0(n25120), .D1(n2890[2]), .SD(n3619), .Z(n25121));
    LUT4 i9307_4_lut_4_lut (.A(n25365), .B(mstatus_mpie), .C(n25372), 
         .D(mstatus_mie), .Z(csr_read_3__N_1170[3])) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i9307_4_lut_4_lut.init = 16'h4f40;
    PFUMX i21124 (.BLUT(\mem_data_from_read[1] ), .ALUT(\mem_data_from_read[5] ), 
          .C0(counter_hi[2]), .Z(n23399));
    PFUMX i22507 (.BLUT(n25119), .ALUT(n25118), .C0(n25155), .Z(n25120));
    PFUMX i21125 (.BLUT(\mem_data_from_read[9] ), .ALUT(\mem_data_from_read[13] ), 
          .C0(counter_hi[2]), .Z(n23400));
    LUT4 mux_2756_i16_3_lut (.A(instr[12]), .B(n25266), .C(n26598), .Z(n4608[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2756_i16_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_404 (.A(n25238), .B(n25245), .C(n25237), .D(n25281), 
         .Z(n4)) /* synthesis lut_function=(!((B (C (D))+!B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_404.init = 16'h0a88;
    LUT4 mux_1013_i2_3_lut (.A(n22994), .B(n1649[1]), .C(n25338), .Z(instr[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_405 (.A(clk_c_enable_69), .B(n25258), .C(n25249), 
         .D(n25236), .Z(n2242)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_405.init = 16'ha888;
    PFUMX debug_branch_I_23_i3 (.BLUT(n8759), .ALUT(debug_branch_N_571[30]), 
          .C0(n23106), .Z(debug_branch_N_181[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i1_4_lut_adj_406 (.A(clk_c_enable_69), .B(n25258), .C(n20), .D(n25), 
         .Z(n2244)) /* synthesis lut_function=(A (B+!(C+(D)))) */ ;
    defparam i1_4_lut_adj_406.init = 16'h888a;
    LUT4 i21882_2_lut_3_lut_4_lut (.A(is_store), .B(clk_c_enable_54), .C(mem_op[1]), 
         .D(rst_reg_n), .Z(data_write_n_1__N_100[1])) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i21882_2_lut_3_lut_4_lut.init = 16'hf7ff;
    LUT4 i11460_2_lut_3_lut_4_lut (.A(is_store), .B(clk_c_enable_54), .C(mem_op[0]), 
         .D(rst_reg_n), .Z(data_write_n_1__N_100[0])) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i11460_2_lut_3_lut_4_lut.init = 16'hf7ff;
    LUT4 i1_4_lut_adj_407 (.A(n25284), .B(instr[12]), .C(n25227), .D(n25212), 
         .Z(n20641)) /* synthesis lut_function=(!((B (C+(D))+!B !((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_407.init = 16'h220a;
    FD1S3IX counter_hi_3136__i4_rep_708 (.D(n17_adj_2394[2]), .CK(clk_c), 
            .CD(n25424), .Q(n26608));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3136__i4_rep_708.GSR = "DISABLED";
    LUT4 next_instr_write_offset_3__I_0_i2_2_lut_rep_536_3_lut_4_lut (.A(n25336), 
         .B(instr_addr_23__N_49[0]), .C(\pc[2] ), .D(instr_addr_23__N_49[1]), 
         .Z(n25272)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam next_instr_write_offset_3__I_0_i2_2_lut_rep_536_3_lut_4_lut.init = 16'h8778;
    PFUMX debug_branch_I_23_i1 (.BLUT(n8755), .ALUT(debug_branch_N_571[28]), 
          .C0(n23106), .Z(debug_branch_N_181[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i1_3_lut_4_lut_adj_408 (.A(n25336), .B(instr_addr_23__N_49[0]), 
         .C(\instr_write_offset[3] ), .D(instr_addr_23__N_49[1]), .Z(n21868)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i1_3_lut_4_lut_adj_408.init = 16'h78f0;
    LUT4 i1_4_lut_adj_409 (.A(instr[12]), .B(n26612), .C(n25288), .D(n25279), 
         .Z(n22214)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_409.init = 16'hc088;
    LUT4 i1_4_lut_adj_410 (.A(instr[12]), .B(n26612), .C(n25290), .D(n25279), 
         .Z(n22226)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_410.init = 16'hc088;
    LUT4 i1_4_lut_4_lut_adj_411 (.A(n25178), .B(n22038), .C(n6), .D(n25171), 
         .Z(n22044)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_411.init = 16'h4000;
    LUT4 i1_4_lut_4_lut_adj_412 (.A(n25178), .B(n22062), .C(n6), .D(n25171), 
         .Z(n22068)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_412.init = 16'h4000;
    LUT4 i1_2_lut_adj_413 (.A(is_jal_de), .B(n26612), .Z(n21696)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_413.init = 16'h8888;
    LUT4 i1_3_lut_adj_414 (.A(n25179), .B(n7955), .C(n26612), .Z(n22334)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_adj_414.init = 16'h1010;
    LUT4 n24875_bdd_3_lut (.A(n24875), .B(instr[31]), .C(n25209), .Z(n24876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24875_bdd_3_lut.init = 16'hcaca;
    LUT4 n13739_bdd_3_lut_22414 (.A(n1649[14]), .B(n1629[14]), .C(n25338), 
         .Z(n24875)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n13739_bdd_3_lut_22414.init = 16'hacac;
    LUT4 mux_1256_i6_3_lut (.A(n14[5]), .B(n2[5]), .C(n1949), .Z(n1950[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i6_3_lut.init = 16'hcaca;
    LUT4 mux_1260_i6_3_lut (.A(n7[5]), .B(n9[5]), .C(n1969), .Z(n1970[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i6_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_415 (.A(n25177), .B(n8), .C(n25182), .D(n21696), 
         .Z(was_early_branch_N_759)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_415.init = 16'h0200;
    PFUMX i6505 (.BLUT(n23065), .ALUT(n23066), .C0(n25337), .Z(n8761));
    LUT4 i16_4_lut_adj_416 (.A(n21860), .B(clk_c_enable_38), .C(rst_reg_n), 
         .D(n25156), .Z(clk_c_enable_392)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i16_4_lut_adj_416.init = 16'hcfca;
    LUT4 i1_4_lut_adj_417 (.A(n25179), .B(n35), .C(n22286), .D(n26), 
         .Z(n22290)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_417.init = 16'h5040;
    LUT4 i1_3_lut_adj_418 (.A(n25279), .B(n25016), .C(n28), .Z(n26)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_adj_418.init = 16'hecec;
    LUT4 i2_4_lut (.A(n25258), .B(clk_c_enable_69), .C(n25249), .D(n25245), 
         .Z(n3619)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'hc888;
    LUT4 i1_4_lut_adj_419 (.A(instr[12]), .B(n26612), .C(n25289), .D(n25279), 
         .Z(n22202)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_419.init = 16'hc088;
    LUT4 mux_346_i1_3_lut_4_lut (.A(n25336), .B(instr_addr_23__N_49[0]), 
         .C(debug_ret), .D(return_addr[1]), .Z(n1764[0])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam mux_346_i1_3_lut_4_lut.init = 16'hf606;
    LUT4 i38_3_lut (.A(n26597), .B(n25281), .C(n24_adj_2391), .Z(n22)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;
    defparam i38_3_lut.init = 16'h9898;
    LUT4 next_instr_write_offset_3__I_0_i1_2_lut_3_lut (.A(n25336), .B(instr_addr_23__N_49[0]), 
         .C(\pc[1] ), .Z(n1)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam next_instr_write_offset_3__I_0_i1_2_lut_3_lut.init = 16'h9696;
    LUT4 i21866_4_lut (.A(n25182), .B(rst_reg_n), .C(n20952), .D(n21966), 
         .Z(clk_c_enable_218)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i21866_4_lut.init = 16'h3337;
    LUT4 mux_1256_i7_3_lut (.A(n14[6]), .B(n2[6]), .C(n1949), .Z(n1950[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i7_3_lut.init = 16'hcaca;
    PFUMX i20784 (.BLUT(\mem_data_from_read[24] ), .ALUT(\mem_data_from_read[28] ), 
          .C0(counter_hi[2]), .Z(n23059));
    LUT4 mux_1260_i7_3_lut (.A(n7[6]), .B(n9[6]), .C(n1969), .Z(n1970[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1559_i12_3_lut_4_lut (.A(n25155), .B(n25152), .C(n2854[11]), 
         .D(n2414[9]), .Z(n2937[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1559_i12_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i21685_3_lut_4_lut (.A(n25278), .B(n25153), .C(n3611), .D(n21230), 
         .Z(n2813[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21685_3_lut_4_lut.init = 16'hf808;
    PFUMX i20787 (.BLUT(\mem_data_from_read[26] ), .ALUT(\mem_data_from_read[30] ), 
          .C0(counter_hi[2]), .Z(n23062));
    LUT4 mux_1256_i3_3_lut (.A(n14[2]), .B(n2[2]), .C(n1949), .Z(n1950[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i3_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_420 (.A(n25279), .B(n25267), .C(n26612), .Z(n22146)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_420.init = 16'h4040;
    LUT4 mux_1540_i1_4_lut (.A(n22004), .B(n7955), .C(n3613), .D(n22160), 
         .Z(n22933)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1540_i1_4_lut.init = 16'h3a0a;
    LUT4 mux_1260_i3_3_lut (.A(n7[2]), .B(n9[2]), .C(n1969), .Z(n1970[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1007_i5_rep_91_3_lut (.A(n9[4]), .B(n14[4]), .C(n1969), .Z(n22970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i5_rep_91_3_lut.init = 16'hcaca;
    LUT4 mux_1003_i5_rep_80_3_lut (.A(n2[4]), .B(n7[4]), .C(n1949), .Z(n22959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i5_rep_80_3_lut.init = 16'hcaca;
    LUT4 is_jalr_N_1103_bdd_4_lut_22479 (.A(n25227), .B(n26597), .C(n25281), 
         .D(n25212), .Z(n24913)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A ((C)+!B))) */ ;
    defparam is_jalr_N_1103_bdd_4_lut_22479.init = 16'h0c2c;
    LUT4 mux_1256_i4_3_lut (.A(n14[3]), .B(n2[3]), .C(n1949), .Z(n1950[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1256_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1260_i4_3_lut (.A(n7[3]), .B(n9[3]), .C(n1969), .Z(n1970[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1260_i4_3_lut.init = 16'hcaca;
    PFUMX i29 (.BLUT(n11), .ALUT(n13), .C0(n26598), .Z(n16_adj_2392));
    LUT4 mux_1007_i6_rep_89_3_lut (.A(n9[5]), .B(n14[5]), .C(n1969), .Z(n22968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i6_rep_89_3_lut.init = 16'hcaca;
    LUT4 mux_1003_i6_rep_78_3_lut (.A(n2[5]), .B(n7[5]), .C(n1949), .Z(n22957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i6_rep_78_3_lut.init = 16'hcaca;
    LUT4 mux_1007_i7_rep_95_3_lut (.A(n9[6]), .B(n14[6]), .C(n1969), .Z(n22974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i7_rep_95_3_lut.init = 16'hcaca;
    LUT4 mux_1003_i7_rep_85_3_lut (.A(n2[6]), .B(n7[6]), .C(n1949), .Z(n22964)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i7_rep_85_3_lut.init = 16'hcaca;
    LUT4 mux_1007_i8_rep_93_3_lut (.A(n9[7]), .B(n14[7]), .C(n1969), .Z(n22972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i8_rep_93_3_lut.init = 16'hcaca;
    LUT4 mux_1003_i8_rep_87_3_lut (.A(n2[7]), .B(n7[7]), .C(n1949), .Z(n22966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i8_rep_87_3_lut.init = 16'hcaca;
    LUT4 mux_1007_i11_3_lut (.A(n9[10]), .B(n14[10]), .C(n1969), .Z(n1649[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i11_3_lut.init = 16'hcaca;
    PFUMX i22453 (.BLUT(n25028), .ALUT(n25027), .C0(mem_data_ready), .Z(n25029));
    LUT4 mux_1003_i11_rep_99_3_lut (.A(n2[10]), .B(n7[10]), .C(n1949), 
         .Z(n22978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i11_rep_99_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_421 (.A(n25178), .B(n22074), .C(n6), .D(n25171), 
         .Z(n22080)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_421.init = 16'h4000;
    LUT4 mux_1007_i4_3_lut (.A(n9[3]), .B(n14[3]), .C(n1969), .Z(n1649[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1003_i4_3_lut (.A(n2[3]), .B(n7[3]), .C(n1949), .Z(n1629[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1007_i9_3_lut (.A(n9[8]), .B(n14[8]), .C(n1969), .Z(n1649[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1003_i9_3_lut (.A(n2[8]), .B(n7[8]), .C(n1949), .Z(n1629[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i9_3_lut.init = 16'hcaca;
    LUT4 mem_data_from_read_6__bdd_4_lut (.A(counter_hi[3]), .B(\data_from_read[6] ), 
         .C(\data_from_read[2] ), .D(counter_hi[2]), .Z(n24927)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam mem_data_from_read_6__bdd_4_lut.init = 16'he4f0;
    LUT4 n24930_bdd_3_lut_22634 (.A(n24930), .B(n25443), .C(counter_hi[3]), 
         .Z(n24931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24930_bdd_3_lut_22634.init = 16'hcaca;
    PFUMX i22442 (.BLUT(n25015), .ALUT(n25014), .C0(n23899), .Z(n25016));
    LUT4 mem_data_from_read_4__bdd_4_lut (.A(counter_hi[3]), .B(\data_from_read[0] ), 
         .C(\data_from_read[2] ), .D(counter_hi[2]), .Z(n24933)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam mem_data_from_read_4__bdd_4_lut.init = 16'hf0e4;
    LUT4 mux_1517_i11_4_lut (.A(n25290), .B(n25206), .C(n3613), .D(n26598), 
         .Z(n2703[10])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1517_i11_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_rep_426_4_lut (.A(n25178), .B(n21944), .C(n25164), .D(n10_c), 
         .Z(n25162)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_rep_426_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_422 (.A(n20952), .B(n25163), .C(instr_fetch_restart_N_678), 
         .D(n25304), .Z(start_instr)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(435[34:115])
    defparam i1_4_lut_adj_422.init = 16'h0040;
    LUT4 i3997_2_lut_rep_555_4_lut_4_lut (.A(n25372), .B(mtime_out[0]), 
         .C(n25329), .D(cy_adj_2388), .Z(n25291)) /* synthesis lut_function=(A (B (D))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i3997_2_lut_rep_555_4_lut_4_lut.init = 16'hc840;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n25372), .B(alu_a_in[0]), .C(n25352), 
         .D(cy_adj_2387), .Z(n22558)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h369c;
    LUT4 i1_rep_10_4_lut (.A(is_ret_de), .B(n25177), .C(n8), .D(n20807), 
         .Z(n20952)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[18] 227[12])
    defparam i1_rep_10_4_lut.init = 16'h0800;
    LUT4 n24936_bdd_3_lut (.A(n24936), .B(n25440), .C(counter_hi[3]), 
         .Z(n24937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24936_bdd_3_lut.init = 16'hcaca;
    LUT4 i21681_3_lut_4_lut (.A(n3613), .B(n3605), .C(n2703[8]), .D(n2414[8]), 
         .Z(n2854[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i21681_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_3_lut_adj_423 (.A(n35), .B(n26_adj_2389), .C(n22254), .Z(n22258)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_423.init = 16'h8080;
    PFUMX i22541 (.BLUT(n25467), .ALUT(n25468), .C0(n25338), .Z(instr[12]));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n25372), .B(n25333), .C(n25293), 
         .D(n25316), .Z(clk_c_enable_111)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hfdfc;
    PFUMX i22435 (.BLUT(n25005), .ALUT(n25004), .C0(n25281), .Z(n22_adj_2374));
    LUT4 i1_2_lut_rep_535_3_lut_4_lut_4_lut (.A(n25372), .B(n25333), .C(interrupt_core), 
         .D(n25344), .Z(n25271)) /* synthesis lut_function=(A (B)+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_2_lut_rep_535_3_lut_4_lut_4_lut.init = 16'hdddc;
    LUT4 tmp_data_in_3__I_99_i4_4_lut_4_lut_4_lut (.A(n25372), .B(data_rs1[3]), 
         .C(interrupt_core), .D(n25344), .Z(tmp_data_in_3__N_1245[3])) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam tmp_data_in_3__I_99_i4_4_lut_4_lut_4_lut.init = 16'h505c;
    PFUMX i22535 (.BLUT(n25456), .ALUT(n25457), .C0(n25418), .Z(n25458));
    LUT4 mux_1007_i10_3_lut (.A(n9[9]), .B(n14[9]), .C(n1969), .Z(n1649[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1007_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1013_i15_3_lut (.A(n1629[14]), .B(n1649[14]), .C(n25338), 
         .Z(instr[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1013_i15_3_lut.init = 16'hcaca;
    PFUMX i22531 (.BLUT(n25450), .ALUT(n25451), .C0(n25338), .Z(instr[4]));
    LUT4 mux_1003_i10_3_lut (.A(n2[9]), .B(n7[9]), .C(n1949), .Z(n1629[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(443[113:125])
    defparam mux_1003_i10_3_lut.init = 16'hcaca;
    PFUMX mux_1013_i14 (.BLUT(n1629[13]), .ALUT(n1649[13]), .C0(n25338), 
          .Z(instr[29]));
    LUT4 i12059_4_lut_4_lut (.A(n25372), .B(\imm[1] ), .C(mcause[2]), 
         .D(mstatus_mte), .Z(n7775)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i12059_4_lut_4_lut.init = 16'h5140;
    PFUMX mux_1013_i13 (.BLUT(n1629[12]), .ALUT(n1649[12]), .C0(n25338), 
          .Z(instr[28]));
    PFUMX i22428 (.BLUT(n24998), .ALUT(n24997), .C0(n25370), .Z(n24999));
    tinyQV_time i_timer (.clk_c(clk_c), .n25424(n25424), .mtimecmp_1__N_1672(mtimecmp_1__N_1672), 
            .mtimecmp_3__N_1666(mtimecmp_3__N_1666), .mtimecmp_0__N_1674(mtimecmp_0__N_1674), 
            .time_pulse_r(time_pulse_r), .clk_c_enable_205(clk_c_enable_205), 
            .n25329(n25329), .\mtimecmp[6] (mtimecmp[6]), .\mtimecmp[7] (mtimecmp[7]), 
            .\addr[2] (addr[2]), .timer_data({timer_data}), .\mtime_out[0] (mtime_out[0]), 
            .\mtimecmp[4] (mtimecmp[4]), .\mtimecmp[5] (mtimecmp[5]), .clk_c_enable_206(clk_c_enable_206), 
            .mtimecmp_2__N_1670(mtimecmp_2__N_1670), .timer_interrupt(timer_interrupt), 
            .n8527(n8527), .cy(cy_adj_2388), .rst_reg_n(rst_reg_n), .n26597(n26597), 
            .n25281(n25281), .\instr_len_2__N_307[1] (instr_len_2__N_307[1]), 
            .n26612(n26612), .no_write_in_progress(no_write_in_progress), 
            .is_store(is_store), .n25350(n25350), .n25178(n25178), .n25175(n25175), 
            .n22126(n22126), .clk_c_enable_84(clk_c_enable_84), .n25365(n25365), 
            .clk_c_enable_328(clk_c_enable_328), .clk_c_enable_54(clk_c_enable_54), 
            .n20762(n20762), .n25372(n25372), .clk_c_enable_324(clk_c_enable_324), 
            .clk_c_enable_352(clk_c_enable_352), .n11558(n11558), .clk_c_enable_344(clk_c_enable_344), 
            .\instr_addr_23__N_49[1] (instr_addr_23__N_49[1]), .\instr_addr_23__N_49[0] (instr_addr_23__N_49[0]), 
            .n22016(n22016), .n25422(n25422), .n5(n5_adj_2393), .clk_c_enable_309(clk_c_enable_309), 
            .n22022(n22022), .\reg_access[3][2] (\reg_access[3] [2]), .clk_c_enable_332(clk_c_enable_332), 
            .\instr_data[0] (instr_data[0]), .\instr_data_0__15__N_369[0] (instr_data_0__15__N_369[0]), 
            .\reg_access[4][3] (\reg_access[4] [3]), .clk_c_enable_348(clk_c_enable_348), 
            .\instr_data[1] (instr_data[1]), .\instr_data_0__15__N_369[49] (instr_data_0__15__N_369[49]), 
            .\cycle_count_wide[3] (cycle_count_wide[3]), .n25246(n25246), 
            .clk_c_enable_170(clk_c_enable_170), .n25432(n25432), .is_timer_addr(is_timer_addr), 
            .n25291(n25291), .n20805(n20805), .data_ready_sync(data_ready_sync), 
            .clk_c_enable_314(clk_c_enable_314), .n25305(n25305), .\data_out_slice[2] (data_out_slice[2]), 
            .n25269(n25269), .\data_out_slice[1] (data_out_slice[1]), .\data_out_slice[0] (data_out_slice[0]), 
            .n25277(n25277)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(450[17] 461[6])
    tinyqv_decoder i_decoder (.n24956(n24956), .n25281(n25281), .n26597(n26597), 
            .is_alu_imm_de(is_alu_imm_de), .n25258(n25258), .n35(n35), 
            .n26612(n26612), .clk_c_enable_38(clk_c_enable_38), .n3611(n3611), 
            .n24919(n24919), .n25284(n25284), .n24894(n24894), .n25227(n25227), 
            .n13701(n13701), .is_ret_de(is_ret_de), .n22839(n22839), .n25262(n25262), 
            .n25261(n25261), .n22398(n22398), .n25288(n25288), .n26598(n26598), 
            .n25287(n25287), .n22384(n22384), .n25265(n25265), .n25267(n25267), 
            .\instr[4] (instr[4]), .n25264(n25264), .n20820(n20820), .n25266(n25266), 
            .n20650(n20650), .n3597(n3597), .\additional_mem_ops[2] (additional_mem_ops[2]), 
            .n4031(n4030[2]), .n26(n26), .n3613(n3613), .clk_c_enable_69(clk_c_enable_69), 
            .n23341(n23341), .n25155(n25155), .n16(n16_adj_2392), .rst_reg_n(rst_reg_n), 
            .n22(n22), .n3589(n3589), .n25153(n25153), .n19(n19), .n3605(n3605), 
            .n25279(n25279), .n25231(n25231), .n25278(n25278), .n25247(n25247), 
            .n25249(n25249), .n21978(n21978), .\instr[12] (instr[12]), 
            .n25256(n25256), .n24939(n24939), .n25290(n25290), .n25260(n25260), 
            .n24940(n24940), .\alu_op_3__N_901[2] (alu_op_3__N_901[2]), 
            .n25234(n25234), .\instr[26] (instr[26]), .n25239(n25239), 
            .n22086(n22086), .n25202(n25202), .n25257(n25257), .is_store_de(is_store_de), 
            .n2438(n2414[8]), .n25214(n25214), .\instr[30] (instr[30]), 
            .n3(n3), .n28(n28), .n25259(n25259), .n25212(n25212), .n25241(n25241), 
            .n25243(n25243), .n25209(n25209), .n25216(n25216), .n10(n10_adj_2390), 
            .n24(n24_adj_2391), .n25210(n25210), .n12(n12), .n26596(n26596), 
            .n25211(n25211), .n25189(n25189), .n22202(n22202), .n7955(n7955), 
            .n26_adj_4(n26_adj_2389), .n22208(n22208), .\instr[31] (instr[31]), 
            .n4532(n4516[15]), .\alu_op_3__N_1068[2] (alu_op_3__N_1068[2]), 
            .n22146(n22146), .n22152(n22152), .\instr[27] (instr[27]), 
            .n157(n155[2]), .n25221(n25221), .n13814(n13814), .n25248(n25248), 
            .\mem_op_de[2] (mem_op_de[2]), .n25226(n25226), .n2797(n2772[7]), 
            .n25196(n25196), .n22867(n22867), .\instr[20] (instr[20]), 
            .n25167(n25167), .n21594(n21594), .n26289(n26289), .n27(n27), 
            .n25245(n25245), .n25244(n25244), .is_branch_de(is_branch_de), 
            .n25208(n25208), .n25338(n25338), .n3615(n3615), .n23255(n23255), 
            .\instr[16] (instr[16]), .n2055(n2052[1]), .n27_adj_5(n27_adj_2381), 
            .n22470(n22470), .n25207(n25207), .n7734(n7734), .n25203(n25203), 
            .n22286(n22286), .\instr[25] (instr[25]), .n2799(n2772[5]), 
            .n25166(n25166), .n4533(n4516[14]), .n1655(n1649[10]), .n25289(n25289), 
            .n22976(n22976), .mem_op_increment_reg_de(mem_op_increment_reg_de), 
            .n25014(n25014), .n7375(n7375), .n25225(n25225), .n6647(n6647), 
            .n25222(n25222), .n22_adj_6(n22_adj_2374), .n2240(n2240), 
            .n15(n15_adj_2383), .n23899(n23899), .alu_op_de({alu_op_de}), 
            .n4534(n4516[13]), .n4535(n4516[12]), .n15_adj_7(n15_adj_2380), 
            .n23900(n23900), .n4531(n4516[16]), .n25228(n25228), .n2437(n2414[9]), 
            .is_alu_reg_de(is_alu_reg_de), .n22226(n22226), .n22232(n22232), 
            .is_system_de(is_system_de), .is_jalr_N_1101(is_jalr_N_1101), 
            .is_jalr_de(is_jalr_de), .n4547(n4516[0]), .n4542(n4516[5]), 
            .n4540(n4516[7]), .n3619(n3619), .n23245(n23245), .n8(n8_adj_2384), 
            .n23379(n23379), .is_load_de(is_load_de), .n4543(n4516[4]), 
            .n20720(n20720), .is_lui_N_1096(is_lui_N_1096), .is_lui_de(is_lui_de), 
            .n25190(n25190), .n2430(n2414[16]), .is_auipc_de(is_auipc_de), 
            .\mem_op_de[1] (mem_op_de[1]), .n2242(n2242), .\instr[17] (instr[17]), 
            .n2049(n2047[2]), .n2077(n2075[2]), .n22126(n22126), .n25182(n25182), 
            .n25177(n25177), .n10_adj_8(n10_c), .n15_adj_9(n15_adj_2382), 
            .n22254(n22254), .n22238(n22238), .n22244(n22244), .n25178(n25178), 
            .n25171(n25171), .n25158(n25158), .n3603(n3603), .n21998(n21998), 
            .n22004(n22004), .n22178(n22178), .n22184(n22184), .n4(n4), 
            .n22120(n22120), .is_jal_de(is_jal_de), .n2658(n2627[1]), 
            .n22132(n22132), .n22138(n22138), .n25156(n25156), .n22276(n22276), 
            .n22214(n22214), .n22220(n22220)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    tinyqv_core i_core (.clk_c(clk_c), .n25273(n25273), .clk_c_enable_27(clk_c_enable_27), 
            .\mie[0] (mie[0]), .n92({n92}), .instr_retired(instr_retired), 
            .instr_complete_N_1378(instr_complete_N_1378), .n25424(n25424), 
            .cmp(cmp), .\imm[11] (\imm[11] ), .instr_complete_N_1382(instr_complete_N_1382), 
            .\next_fsm_state_3__N_2230[3] (\next_fsm_state_3__N_2230[3] ), 
            .cy(cy_adj_2387), .mstatus_mte(mstatus_mte), .clk_c_enable_111(clk_c_enable_111), 
            .mstatus_mpie(mstatus_mpie), .clk_c_enable_170(clk_c_enable_170), 
            .\addr_out[11] (addr_out[11]), .\addr_out[12] (addr_out[12]), 
            .\addr_out[13] (addr_out[13]), .\addr_out[14] (addr_out[14]), 
            .\addr_out[15] (addr_out[15]), .counter_hi({counter_hi}), .\addr_out[16] (addr_out[16]), 
            .\addr_out[17] (addr_out[17]), .\addr_out[18] (addr_out[18]), 
            .\addr_out[19] (addr_out[19]), .n25372(n25372), .n25365(n25365), 
            .\addr_out[20] (addr_out[20]), .\addr_out[21] (addr_out[21]), 
            .\addr_out[22] (addr_out[22]), .\imm[6] (\imm[6] ), .\addr_out[23] (addr_out[23]), 
            .\alu_op[1] (alu_op[1]), .debug_instr_valid(debug_instr_valid), 
            .is_system(is_system), .\alu_op[0] (alu_op[0]), .n25310(n25310), 
            .n5(n5), .clk_c_enable_205(clk_c_enable_205), .n25344(n25344), 
            .\imm[1] (\imm[1] ), .cycle_count_wide({Open_31, Open_32, 
            Open_33, cycle_count_wide[3], Open_34, cycle_count_wide[1:0]}), 
            .\imm[0] (imm[0]), .\next_pc_for_core[22] (\next_pc_for_core[22] ), 
            .\next_pc_for_core[18] (\next_pc_for_core[18] ), .\mie[8] (mie[8]), 
            .data_rs1({Open_35, Open_36, Open_37, data_rs1[0]}), .n25179(n25179), 
            .n25175(n25175), .n22208(n22208), .n25178(n25178), .n21248(n21248), 
            .n22098(n22098), .n3615(n3615), .timer_interrupt(timer_interrupt), 
            .n26608(n26608), .n22172(n22172), .n2037(n2034[1]), .n22258(n22258), 
            .n2835(n2813[10]), .n22867(n22867), .n7955(n7955), .n24916(n24916), 
            .n22272(n22272), .n22152(n22152), .n21113(n21113), .\alu_op_in[2] (alu_op_in[2]), 
            .n25430(n25430), .n22254(n22254), .n26(n26_adj_2389), .n24486(n24486), 
            .n22184(n22184), .n21260(n21260), .n22244(n22244), .n21230(n21230), 
            .n22138(n22138), .n21121(n21121), .n22004(n22004), .n25182(n25182), 
            .n25177(n25177), .n22008(n22008), .n22324(n22324), .n21303(n21303), 
            .n22298(n22298), .n21297(n21297), .n22120(n22120), .n2236(n2236), 
            .n22220(n22220), .n21242(n21242), .n25216(n25216), .n21910(n21910), 
            .n21916(n21916), .n22933(n22933), .n22852(n22852), .n22086(n22086), 
            .n25191(n25191), .n22092(n22092), .n22276(n22276), .n12(n12), 
            .n22282(n22282), .n21898(n21898), .n21212(n21212), .n22232(n22232), 
            .n21236(n21236), .n23322(n23322), .\cycle[0] (\cycle[0] ), 
            .\addr_out[3] (addr_out[3]), .n11558(n11558), .\ui_in_sync[1] (\ui_in_sync[1] ), 
            .n1092(n1092), .n25343(n25343), .n26610(n26610), .any_additional_mem_ops(any_additional_mem_ops), 
            .clk_c_enable_206(clk_c_enable_206), .n25349(n25349), .interrupt_core(interrupt_core), 
            .clk_c_enable_209(clk_c_enable_209), .is_load(is_load), .n54(n54), 
            .n20739(n20739), .clk_c_enable_393(clk_c_enable_393), .n21402(n21402), 
            .n4455({n4455}), .n1768({n1768}), .pc_2__N_663({pc_2__N_663}), 
            .load_done(load_done), .n6638(n6638), .n1767(n1764[0]), .\instr_write_offset_3__N_665[0] (instr_write_offset_3__N_665[0]), 
            .n1766(n1764[1]), .\instr_write_offset_3__N_665[1] (instr_write_offset_3__N_665[1]), 
            .n25181(n25181), .mem_op({mem_op}), .n5031(n5029[2]), .\addr_out[6] (addr_out[6]), 
            .debug_rd({debug_rd}), .debug_rd_3__N_1306(debug_rd_3__N_1306), 
            .\addr_out[7] (addr_out[7]), .n25369(n25369), .\imm[2] (\imm[2] ), 
            .n25410(n25410), .accum({accum}), .d_3__N_1599({d_3__N_1599}), 
            .\imm[7] (\imm[7] ), .\imm[8] (\imm[8] ), .\imm[10] (\imm[10] ), 
            .\imm[9] (\imm[9] ), .n24938(n24938), .\debug_branch_N_181[0] (debug_branch_N_181[0]), 
            .\addr_out[4] (addr_out[4]), .\mul_out[1] (\mul_out[1] ), .n25421(n25421), 
            .data_rs2({data_rs2}), .\debug_rd_3__N_136[28] (debug_rd_3__N_136[28]), 
            .alu_b_in({Open_38, Open_39, Open_40, alu_b_in[0]}), .n25316(n25316), 
            .\addr_out[8] (addr_out[8]), .\mul_out[3] (\mul_out[3] ), .\mcause[2] (mcause[2]), 
            .\alu_b_in[1] (alu_b_in[1]), .\alu_a_in[1] (alu_a_in[1]), .n5047({n5047}), 
            .\alu_a_in[0] (alu_a_in[0]), .n6657(n6657), .was_early_branch(was_early_branch), 
            .instr_fetch_restart_N_678(instr_fetch_restart_N_678), .data_out_3__N_1116(data_out_3__N_1116), 
            .\data_out_slice[1] (data_out_slice[1]), .n22354(n22354), .mstatus_mie(mstatus_mie), 
            .n21750(n21750), .n22028(n22028), .n22030(n22030), .n25180(n25180), 
            .rst_reg_n(rst_reg_n), .n14111(n14111), .n20807(n20807), .\next_pc_offset[3] (next_pc_offset[3]), 
            .n21864(n21864), .n25422(n25422), .n5_adj_1(n5_adj_2393), 
            .clk_c_enable_54(clk_c_enable_54), .\addr_out[10] (addr_out[10]), 
            .\debug_branch_N_173[28] (debug_branch_N_173[28]), .n22941(n22941), 
            .\addr_out[0] (addr_out[0]), .n25411(n25411), .n25333(n25333), 
            .n25359(n25359), .\next_pc_for_core[15] (\next_pc_for_core[15] ), 
            .\next_pc_for_core[11] (\next_pc_for_core[11] ), .load_top_bit(load_top_bit), 
            .\debug_branch_N_181[3] (debug_branch_N_181[3]), .n25352(n25352), 
            .cy_adj_2(cy_adj_2386), .data_ready_sync(data_ready_sync), .n25197(n25197), 
            .data_ready_core(data_ready_core), .n24186(n24186), .cy_adj_3(cy), 
            .\addr_out[5] (addr_out[5]), .\instrret_count[0] (instrret_count[0]), 
            .n23011(n23011), .n25408(n25408), .\debug_branch_N_173[30] (debug_branch_N_173[30]), 
            .n25402(n25402), .n25350(n25350), .clk_c_enable_336(clk_c_enable_336), 
            .n18(n17_adj_2394[2]), .clk_c_enable_197(clk_c_enable_197), 
            .n23898(n23898), .n23897(n23897), .n23896(n23896), .n23895(n23895), 
            .n23894(n23894), .\imm[4] (\imm[4] ), .\addr_out[26] (addr_out[26]), 
            .n25307(n25307), .\addr_out[25] (addr_out[25]), .\addr_out[24] (addr_out[24]), 
            .\alu_op[3] (alu_op[3]), .is_alu_imm(is_alu_imm), .is_alu_reg(is_alu_reg), 
            .is_auipc(is_auipc), .\debug_branch_N_173[29] (debug_branch_N_173[29]), 
            .is_jal(is_jal), .n25426(n25426), .\debug_rd_3__N_136[29] (debug_rd_3__N_136[29]), 
            .n4996(n4994[2]), .n24264(n24264), .is_jalr(is_jalr), .n25412(n25412), 
            .n23395(n23395), .is_lui(is_lui), .is_store(is_store), .\data_out_slice[0] (data_out_slice[0]), 
            .\debug_branch_N_571[29] (debug_branch_N_571[29]), .\timer_data[1] (timer_data[1]), 
            .is_timer_addr(is_timer_addr), .\imm[5] (\imm[5] ), .\imm[3] (\imm[3] ), 
            .is_branch(is_branch), .n25277(n25277), .\data_rs1[3] (data_rs1[3]), 
            .n23111(n23111), .n25375(n25375), .n22798(n22798), .n25387(n25387), 
            .\debug_rd_3__N_136[31] (debug_rd_3__N_136[31]), .\tmp_data_in_3__N_1245[3] (tmp_data_in_3__N_1245[3]), 
            .n25319(n25319), .\debug_rd_3__N_136[30] (debug_rd_3__N_136[30]), 
            .\addr_out[9] (addr_out[9]), .\debug_branch_N_173[31] (debug_branch_N_173[31]), 
            .n25301(n25301), .\debug_rd_3__N_1298[0] (debug_rd_3__N_1298[0]), 
            .n25293(n25293), .n25282(n25282), .\mtimecmp[7] (mtimecmp[7]), 
            .mtimecmp_3__N_1666(mtimecmp_3__N_1666), .\data_out_slice[2] (data_out_slice[2]), 
            .n24932(n24932), .\debug_branch_N_181[2] (debug_branch_N_181[2]), 
            .no_write_in_progress(no_write_in_progress), .n25348(n25348), 
            .n25326(n25326), .n23069(n23069), .\addr_out[1] (addr_out[1]), 
            .n22944(n22944), .\debug_branch_N_571[31] (debug_branch_N_571[31]), 
            .n23073(n23073), .\debug_branch_N_177[31] (debug_branch_N_177[31]), 
            .\mul_out[2] (\mul_out[2] ), .n23067(n23067), .\debug_branch_N_177[29] (debug_branch_N_177[29]), 
            .\next_pc_for_core[14] (\next_pc_for_core[14] ), .\next_pc_for_core[10] (\next_pc_for_core[10] ), 
            .n66(n66), .n12257(n12257), .\addr_offset[2] (addr_offset[2]), 
            .n701(n699[0]), .n23070(n23070), .\debug_branch_N_177[30] (debug_branch_N_177[30]), 
            .n25341(n25341), .n25271(n25271), .n22939(n22939), .n23012(n23012), 
            .n25475(n25475), .\csr_read_3__N_1170[3] (csr_read_3__N_1170[3]), 
            .\next_accum[6] (\next_accum[6] ), .\next_accum[7] (\next_accum[7] ), 
            .\next_accum[8] (\next_accum[8] ), .\next_accum[9] (\next_accum[9] ), 
            .\next_accum[10] (\next_accum[10] ), .\next_accum[11] (\next_accum[11] ), 
            .\next_accum[12] (\next_accum[12] ), .\next_accum[13] (\next_accum[13] ), 
            .\next_accum[14] (\next_accum[14] ), .\next_accum[15] (\next_accum[15] ), 
            .GND_net(GND_net), .VCC_net(VCC_net), .\next_accum[16] (\next_accum[16] ), 
            .\next_accum[17] (\next_accum[17] ), .\next_accum[18] (\next_accum[18] ), 
            .\next_accum[19] (\next_accum[19] ), .\next_accum[5] (\next_accum[5] ), 
            .\next_accum[4] (\next_accum[4] ), .rs2({rs2}), .rs1({rs1}), 
            .rd({rd}), .return_addr({return_addr}), .\reg_access[4][3] (\reg_access[4] [3]), 
            .\reg_access[3][2] (\reg_access[3] [2]), .\instr[12] (instr[12]), 
            .n3645(n3641[0]), .\increment_result_3__N_1656[0] (increment_result_3__N_1656[0]), 
            .n25294(n25294), .\increment_result_3__N_1642[1] (increment_result_3__N_1642[1]), 
            .n25246(n25246), .n22558(n22558), .n25218(n25218), .n21812(n21812)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(322[72] 368[6])
    
endmodule
//
// Verilog Description of module tinyQV_time
//

module tinyQV_time (clk_c, n25424, mtimecmp_1__N_1672, mtimecmp_3__N_1666, 
            mtimecmp_0__N_1674, time_pulse_r, clk_c_enable_205, n25329, 
            \mtimecmp[6] , \mtimecmp[7] , \addr[2] , timer_data, \mtime_out[0] , 
            \mtimecmp[4] , \mtimecmp[5] , clk_c_enable_206, mtimecmp_2__N_1670, 
            timer_interrupt, n8527, cy, rst_reg_n, n26597, n25281, 
            \instr_len_2__N_307[1] , n26612, no_write_in_progress, is_store, 
            n25350, n25178, n25175, n22126, clk_c_enable_84, n25365, 
            clk_c_enable_328, clk_c_enable_54, n20762, n25372, clk_c_enable_324, 
            clk_c_enable_352, n11558, clk_c_enable_344, \instr_addr_23__N_49[1] , 
            \instr_addr_23__N_49[0] , n22016, n25422, n5, clk_c_enable_309, 
            n22022, \reg_access[3][2] , clk_c_enable_332, \instr_data[0] , 
            \instr_data_0__15__N_369[0] , \reg_access[4][3] , clk_c_enable_348, 
            \instr_data[1] , \instr_data_0__15__N_369[49] , \cycle_count_wide[3] , 
            n25246, clk_c_enable_170, n25432, is_timer_addr, n25291, 
            n20805, data_ready_sync, clk_c_enable_314, n25305, \data_out_slice[2] , 
            n25269, \data_out_slice[1] , \data_out_slice[0] , n25277) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output n25424;
    input mtimecmp_1__N_1672;
    input mtimecmp_3__N_1666;
    input mtimecmp_0__N_1674;
    output time_pulse_r;
    input clk_c_enable_205;
    output n25329;
    output \mtimecmp[6] ;
    output \mtimecmp[7] ;
    input \addr[2] ;
    output [3:0]timer_data;
    output \mtime_out[0] ;
    output \mtimecmp[4] ;
    output \mtimecmp[5] ;
    input clk_c_enable_206;
    input mtimecmp_2__N_1670;
    output timer_interrupt;
    input n8527;
    output cy;
    input rst_reg_n;
    input n26597;
    input n25281;
    output \instr_len_2__N_307[1] ;
    input n26612;
    input no_write_in_progress;
    input is_store;
    output n25350;
    input n25178;
    input n25175;
    input n22126;
    output clk_c_enable_84;
    input n25365;
    output clk_c_enable_328;
    input clk_c_enable_54;
    output n20762;
    input n25372;
    output clk_c_enable_324;
    output clk_c_enable_352;
    input n11558;
    output clk_c_enable_344;
    input \instr_addr_23__N_49[1] ;
    input \instr_addr_23__N_49[0] ;
    output n22016;
    input n25422;
    input n5;
    output clk_c_enable_309;
    output n22022;
    input \reg_access[3][2] ;
    output clk_c_enable_332;
    input \instr_data[0] ;
    output \instr_data_0__15__N_369[0] ;
    input \reg_access[4][3] ;
    output clk_c_enable_348;
    input \instr_data[1] ;
    output \instr_data_0__15__N_369[49] ;
    input \cycle_count_wide[3] ;
    input n25246;
    output clk_c_enable_170;
    input n25432;
    input is_timer_addr;
    input n25291;
    input n20805;
    input data_ready_sync;
    output clk_c_enable_314;
    input n25305;
    input \data_out_slice[2] ;
    input n25269;
    input \data_out_slice[1] ;
    input \data_out_slice[0] ;
    input n25277;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [31:0]mtimecmp;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(30[16:24])
    wire [3:0]mtime_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(29[16:25])
    
    wire n4, n25447, cy_c;
    wire [4:0]comparison;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[16:26])
    
    wire timer_interrupt_N_1685, n6, n2, n25448;
    
    FD1S3IX mtimecmp_1__91 (.D(mtimecmp_1__N_1672), .CK(clk_c), .CD(n25424), 
            .Q(mtimecmp[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_1__91.GSR = "DISABLED";
    FD1S3IX mtimecmp_3__89 (.D(mtimecmp_3__N_1666), .CK(clk_c), .CD(n25424), 
            .Q(mtimecmp[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_3__89.GSR = "DISABLED";
    FD1S3IX mtimecmp_0__92 (.D(mtimecmp_0__N_1674), .CK(clk_c), .CD(n25424), 
            .Q(mtimecmp[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_0__92.GSR = "DISABLED";
    FD1S3IX time_pulse_r_95 (.D(n25329), .CK(clk_c), .CD(clk_c_enable_205), 
            .Q(time_pulse_r)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(82[12] 85[8])
    defparam time_pulse_r_95.GSR = "DISABLED";
    LUT4 i11682_4_lut_else_4_lut (.A(mtime_out[3]), .B(n4), .C(\mtimecmp[6] ), 
         .D(\mtimecmp[7] ), .Z(n25447)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A (B (C+(D))+!B !(C (D))))) */ ;
    defparam i11682_4_lut_else_4_lut.init = 16'h1824;
    LUT4 mtime_out_3__I_0_96_i3_3_lut (.A(mtime_out[2]), .B(\mtimecmp[6] ), 
         .C(\addr[2] ), .Z(timer_data[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i3_3_lut.init = 16'hcaca;
    LUT4 mtime_out_3__I_0_96_i1_3_lut (.A(\mtime_out[0] ), .B(\mtimecmp[4] ), 
         .C(\addr[2] ), .Z(timer_data[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i1_3_lut.init = 16'hcaca;
    FD1S3AX mtimecmp_30__62 (.D(mtimecmp[2]), .CK(clk_c), .Q(mtimecmp[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_30__62.GSR = "DISABLED";
    FD1S3AX mtimecmp_29__63 (.D(mtimecmp[1]), .CK(clk_c), .Q(mtimecmp[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_29__63.GSR = "DISABLED";
    FD1S3AX mtimecmp_28__64 (.D(mtimecmp[0]), .CK(clk_c), .Q(mtimecmp[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_28__64.GSR = "DISABLED";
    FD1S3AX mtimecmp_27__65 (.D(mtimecmp[31]), .CK(clk_c), .Q(mtimecmp[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_27__65.GSR = "DISABLED";
    FD1S3AX mtimecmp_26__66 (.D(mtimecmp[30]), .CK(clk_c), .Q(mtimecmp[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_26__66.GSR = "DISABLED";
    FD1S3AX mtimecmp_25__67 (.D(mtimecmp[29]), .CK(clk_c), .Q(mtimecmp[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_25__67.GSR = "DISABLED";
    FD1S3AX mtimecmp_24__68 (.D(mtimecmp[28]), .CK(clk_c), .Q(mtimecmp[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_24__68.GSR = "DISABLED";
    FD1S3AX mtimecmp_23__69 (.D(mtimecmp[27]), .CK(clk_c), .Q(mtimecmp[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_23__69.GSR = "DISABLED";
    FD1S3AX mtimecmp_22__70 (.D(mtimecmp[26]), .CK(clk_c), .Q(mtimecmp[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_22__70.GSR = "DISABLED";
    FD1S3AX mtimecmp_21__71 (.D(mtimecmp[25]), .CK(clk_c), .Q(mtimecmp[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_21__71.GSR = "DISABLED";
    FD1S3AX mtimecmp_20__72 (.D(mtimecmp[24]), .CK(clk_c), .Q(mtimecmp[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_20__72.GSR = "DISABLED";
    FD1S3AX mtimecmp_19__73 (.D(mtimecmp[23]), .CK(clk_c), .Q(mtimecmp[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_19__73.GSR = "DISABLED";
    FD1S3AX mtimecmp_18__74 (.D(mtimecmp[22]), .CK(clk_c), .Q(mtimecmp[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_18__74.GSR = "DISABLED";
    FD1S3AX mtimecmp_17__75 (.D(mtimecmp[21]), .CK(clk_c), .Q(mtimecmp[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_17__75.GSR = "DISABLED";
    FD1S3AX mtimecmp_16__76 (.D(mtimecmp[20]), .CK(clk_c), .Q(mtimecmp[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_16__76.GSR = "DISABLED";
    FD1S3AX mtimecmp_15__77 (.D(mtimecmp[19]), .CK(clk_c), .Q(mtimecmp[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_15__77.GSR = "DISABLED";
    FD1S3AX mtimecmp_14__78 (.D(mtimecmp[18]), .CK(clk_c), .Q(mtimecmp[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_14__78.GSR = "DISABLED";
    FD1S3AX mtimecmp_13__79 (.D(mtimecmp[17]), .CK(clk_c), .Q(mtimecmp[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_13__79.GSR = "DISABLED";
    FD1S3AX mtimecmp_12__80 (.D(mtimecmp[16]), .CK(clk_c), .Q(mtimecmp[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_12__80.GSR = "DISABLED";
    FD1S3AX mtimecmp_11__81 (.D(mtimecmp[15]), .CK(clk_c), .Q(mtimecmp[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_11__81.GSR = "DISABLED";
    FD1S3AX mtimecmp_10__82 (.D(mtimecmp[14]), .CK(clk_c), .Q(mtimecmp[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_10__82.GSR = "DISABLED";
    FD1S3AX mtimecmp_9__83 (.D(mtimecmp[13]), .CK(clk_c), .Q(mtimecmp[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_9__83.GSR = "DISABLED";
    FD1S3AX mtimecmp_8__84 (.D(mtimecmp[12]), .CK(clk_c), .Q(mtimecmp[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_8__84.GSR = "DISABLED";
    FD1S3AX mtimecmp_7__85 (.D(mtimecmp[11]), .CK(clk_c), .Q(\mtimecmp[7] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_7__85.GSR = "DISABLED";
    FD1S3AX mtimecmp_6__86 (.D(mtimecmp[10]), .CK(clk_c), .Q(\mtimecmp[6] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_6__86.GSR = "DISABLED";
    FD1S3AX mtimecmp_5__87 (.D(mtimecmp[9]), .CK(clk_c), .Q(\mtimecmp[5] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_5__87.GSR = "DISABLED";
    FD1S3AX mtimecmp_4__88 (.D(mtimecmp[8]), .CK(clk_c), .Q(\mtimecmp[4] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_4__88.GSR = "DISABLED";
    FD1S3JX cy_93 (.D(comparison[4]), .CK(clk_c), .PD(clk_c_enable_206), 
            .Q(cy_c)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(74[12] 76[8])
    defparam cy_93.GSR = "DISABLED";
    FD1S3AX mtimecmp_31__61 (.D(mtimecmp[3]), .CK(clk_c), .Q(mtimecmp[31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_31__61.GSR = "DISABLED";
    FD1S3IX mtimecmp_2__90 (.D(mtimecmp_2__N_1670), .CK(clk_c), .CD(n25424), 
            .Q(mtimecmp[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_2__90.GSR = "DISABLED";
    FD1P3AX timer_interrupt_94 (.D(timer_interrupt_N_1685), .SP(clk_c_enable_206), 
            .CK(clk_c), .Q(timer_interrupt)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(78[12] 80[8])
    defparam timer_interrupt_94.GSR = "DISABLED";
    LUT4 mtime_out_3__I_0_96_i2_3_lut (.A(mtime_out[1]), .B(\mtimecmp[5] ), 
         .C(\addr[2] ), .Z(timer_data[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i2_3_lut.init = 16'hcaca;
    LUT4 i3793_3_lut (.A(mtime_out[3]), .B(\mtimecmp[7] ), .C(n6), .Z(comparison[4])) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i3793_3_lut.init = 16'hb2b2;
    LUT4 i3786_3_lut (.A(mtime_out[2]), .B(\mtimecmp[6] ), .C(n4), .Z(n6)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i3786_3_lut.init = 16'hb2b2;
    LUT4 i3779_3_lut (.A(mtime_out[1]), .B(\mtimecmp[5] ), .C(n2), .Z(n4)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i3779_3_lut.init = 16'hb2b2;
    LUT4 i3772_3_lut (.A(\mtime_out[0] ), .B(\mtimecmp[4] ), .C(cy_c), 
         .Z(n2)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i3772_3_lut.init = 16'hb2b2;
    LUT4 mtime_out_3__I_0_96_i4_3_lut (.A(mtime_out[3]), .B(\mtimecmp[7] ), 
         .C(\addr[2] ), .Z(timer_data[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i4_3_lut.init = 16'hcaca;
    LUT4 i11682_4_lut_then_4_lut (.A(mtime_out[3]), .B(n4), .C(\mtimecmp[6] ), 
         .D(\mtimecmp[7] ), .Z(n25448)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;
    defparam i11682_4_lut_then_4_lut.init = 16'h8241;
    LUT4 time_pulse_I_0_2_lut_rep_593 (.A(n8527), .B(time_pulse_r), .Z(n25329)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(37[14:39])
    defparam time_pulse_I_0_2_lut_rep_593.init = 16'hdddd;
    PFUMX i22529 (.BLUT(n25447), .ALUT(n25448), .C0(mtime_out[2]), .Z(timer_interrupt_N_1685));
    tinyqv_counter i_mtime (.clk_c(clk_c), .n25424(n25424), .cy(cy), .mtime_out({mtime_out[3:1], 
            \mtime_out[0] }), .rst_reg_n(rst_reg_n), .n26597(n26597), 
            .n25281(n25281), .\instr_len_2__N_307[1] (\instr_len_2__N_307[1] ), 
            .n26612(n26612), .no_write_in_progress(no_write_in_progress), 
            .is_store(is_store), .n25350(n25350), .n25178(n25178), .n25175(n25175), 
            .n22126(n22126), .clk_c_enable_84(clk_c_enable_84), .n25365(n25365), 
            .clk_c_enable_328(clk_c_enable_328), .clk_c_enable_54(clk_c_enable_54), 
            .n20762(n20762), .n25372(n25372), .clk_c_enable_324(clk_c_enable_324), 
            .clk_c_enable_206(clk_c_enable_206), .clk_c_enable_352(clk_c_enable_352), 
            .n11558(n11558), .clk_c_enable_344(clk_c_enable_344), .\instr_addr_23__N_49[1] (\instr_addr_23__N_49[1] ), 
            .\instr_addr_23__N_49[0] (\instr_addr_23__N_49[0] ), .n22016(n22016), 
            .n25422(n25422), .n5(n5), .clk_c_enable_309(clk_c_enable_309), 
            .n22022(n22022), .\reg_access[3][2] (\reg_access[3][2] ), .clk_c_enable_332(clk_c_enable_332), 
            .\instr_data[0] (\instr_data[0] ), .\instr_data_0__15__N_369[0] (\instr_data_0__15__N_369[0] ), 
            .\reg_access[4][3] (\reg_access[4][3] ), .clk_c_enable_348(clk_c_enable_348), 
            .\instr_data[1] (\instr_data[1] ), .\instr_data_0__15__N_369[49] (\instr_data_0__15__N_369[49] ), 
            .\cycle_count_wide[3] (\cycle_count_wide[3] ), .n25246(n25246), 
            .clk_c_enable_170(clk_c_enable_170), .\addr[2] (\addr[2] ), 
            .n25432(n25432), .is_timer_addr(is_timer_addr), .n25291(n25291), 
            .n20805(n20805), .data_ready_sync(data_ready_sync), .clk_c_enable_314(clk_c_enable_314), 
            .n25305(n25305), .\data_out_slice[2] (\data_out_slice[2] ), 
            .n25269(n25269), .\data_out_slice[1] (\data_out_slice[1] ), 
            .\data_out_slice[0] (\data_out_slice[0] ), .n25277(n25277)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(34[20] 42[6])
    
endmodule
//
// Verilog Description of module tinyqv_counter
//

module tinyqv_counter (clk_c, n25424, cy, mtime_out, rst_reg_n, n26597, 
            n25281, \instr_len_2__N_307[1] , n26612, no_write_in_progress, 
            is_store, n25350, n25178, n25175, n22126, clk_c_enable_84, 
            n25365, clk_c_enable_328, clk_c_enable_54, n20762, n25372, 
            clk_c_enable_324, clk_c_enable_206, clk_c_enable_352, n11558, 
            clk_c_enable_344, \instr_addr_23__N_49[1] , \instr_addr_23__N_49[0] , 
            n22016, n25422, n5, clk_c_enable_309, n22022, \reg_access[3][2] , 
            clk_c_enable_332, \instr_data[0] , \instr_data_0__15__N_369[0] , 
            \reg_access[4][3] , clk_c_enable_348, \instr_data[1] , \instr_data_0__15__N_369[49] , 
            \cycle_count_wide[3] , n25246, clk_c_enable_170, \addr[2] , 
            n25432, is_timer_addr, n25291, n20805, data_ready_sync, 
            clk_c_enable_314, n25305, \data_out_slice[2] , n25269, \data_out_slice[1] , 
            \data_out_slice[0] , n25277) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output n25424;
    output cy;
    output [3:0]mtime_out;
    input rst_reg_n;
    input n26597;
    input n25281;
    output \instr_len_2__N_307[1] ;
    input n26612;
    input no_write_in_progress;
    input is_store;
    output n25350;
    input n25178;
    input n25175;
    input n22126;
    output clk_c_enable_84;
    input n25365;
    output clk_c_enable_328;
    input clk_c_enable_54;
    output n20762;
    input n25372;
    output clk_c_enable_324;
    input clk_c_enable_206;
    output clk_c_enable_352;
    input n11558;
    output clk_c_enable_344;
    input \instr_addr_23__N_49[1] ;
    input \instr_addr_23__N_49[0] ;
    output n22016;
    input n25422;
    input n5;
    output clk_c_enable_309;
    output n22022;
    input \reg_access[3][2] ;
    output clk_c_enable_332;
    input \instr_data[0] ;
    output \instr_data_0__15__N_369[0] ;
    input \reg_access[4][3] ;
    output clk_c_enable_348;
    input \instr_data[1] ;
    output \instr_data_0__15__N_369[49] ;
    input \cycle_count_wide[3] ;
    input n25246;
    output clk_c_enable_170;
    input \addr[2] ;
    input n25432;
    input is_timer_addr;
    input n25291;
    input n20805;
    input data_ready_sync;
    output clk_c_enable_314;
    input n25305;
    input \data_out_slice[2] ;
    input n25269;
    input \data_out_slice[1] ;
    input \data_out_slice[0] ;
    input n25277;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    wire [4:0]increment_result;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[16:32])
    
    wire n7696;
    wire [4:0]increment_result_3__N_1656;
    
    wire n25268, n25235;
    
    FD1S3IX register_2__48 (.D(increment_result[2]), .CK(clk_c), .CD(n25424), 
            .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result[1]), .CK(clk_c), .CD(n25424), 
            .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(increment_result[0]), .CK(clk_c), .CD(n25424), 
            .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3IX cy_51 (.D(increment_result_3__N_1656[4]), .CK(clk_c), .CD(n7696), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(register[10])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(register[9])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(register[8])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(mtime_out[3])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(register[10]), .CK(clk_c), .Q(mtime_out[2])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(register[9]), .CK(clk_c), .Q(mtime_out[1])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(register[8]), .CK(clk_c), .Q(mtime_out[0])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result[3]), .CK(clk_c), .CD(n25424), 
            .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 rstn_I_0_1_lut_rep_688 (.A(rst_reg_n), .Z(n25424)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam rstn_I_0_1_lut_rep_688.init = 16'h5555;
    LUT4 i11666_2_lut_3_lut_3_lut (.A(rst_reg_n), .B(n26597), .C(n25281), 
         .Z(\instr_len_2__N_307[1] )) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i11666_2_lut_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i3213_3_lut_rep_614_3_lut (.A(n26612), .B(no_write_in_progress), 
         .C(is_store), .Z(n25350)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3213_3_lut_rep_614_3_lut.init = 16'hd5d5;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(n25178), .C(n25175), 
         .D(n22126), .Z(clk_c_enable_84)) /* synthesis lut_function=(!(A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h5575;
    LUT4 i21875_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n25365), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_328)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i21875_2_lut_4_lut_4_lut.init = 16'h3111;
    LUT4 i1_2_lut_3_lut_3_lut (.A(rst_reg_n), .B(clk_c_enable_54), .C(is_store), 
         .Z(n20762)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i21724_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n25372), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_324)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i21724_2_lut_4_lut_4_lut.init = 16'h3111;
    LUT4 i12230_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(clk_c_enable_206), 
         .C(no_write_in_progress), .D(is_store), .Z(clk_c_enable_352)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i12230_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i21868_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n11558), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_344)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i21868_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i1_2_lut_3_lut_3_lut_adj_317 (.A(n26612), .B(\instr_addr_23__N_49[1] ), 
         .C(\instr_addr_23__N_49[0] ), .Z(n22016)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_3_lut_adj_317.init = 16'hf7f7;
    LUT4 i1_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n25422), .C(n5), .D(clk_c_enable_206), 
         .Z(clk_c_enable_309)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_2_lut_3_lut_3_lut_adj_318 (.A(n26612), .B(\instr_addr_23__N_49[0] ), 
         .C(\instr_addr_23__N_49[1] ), .Z(n22022)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_3_lut_adj_318.init = 16'hfdfd;
    LUT4 i21873_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(\reg_access[3][2] ), 
         .C(no_write_in_progress), .D(is_store), .Z(clk_c_enable_332)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i21873_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i11491_2_lut_2_lut (.A(rst_reg_n), .B(\instr_data[0] ), .Z(\instr_data_0__15__N_369[0] )) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i11491_2_lut_2_lut.init = 16'hdddd;
    LUT4 i21867_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(\reg_access[4][3] ), 
         .C(no_write_in_progress), .D(is_store), .Z(clk_c_enable_348)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i21867_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i11628_2_lut_2_lut (.A(rst_reg_n), .B(\instr_data[1] ), .Z(\instr_data_0__15__N_369[49] )) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i11628_2_lut_2_lut.init = 16'hdddd;
    LUT4 i3239_4_lut_4_lut (.A(n26612), .B(\cycle_count_wide[3] ), .C(n25246), 
         .D(clk_c_enable_206), .Z(clk_c_enable_170)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3239_4_lut_4_lut.init = 16'hd555;
    LUT4 i5466_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(\addr[2] ), .C(n25432), 
         .D(is_timer_addr), .Z(n7696)) /* synthesis lut_function=(!(A (B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i5466_2_lut_3_lut_4_lut_4_lut.init = 16'h5755;
    LUT4 i4019_2_lut_3_lut_4_lut (.A(mtime_out[1]), .B(n25291), .C(mtime_out[3]), 
         .D(mtime_out[2]), .Z(increment_result_3__N_1656[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4019_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut (.A(n20762), .B(n20805), .C(data_ready_sync), .D(clk_c_enable_206), 
         .Z(clk_c_enable_314)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_4_lut.init = 16'hfbbb;
    LUT4 i4005_2_lut_rep_532_3_lut (.A(mtime_out[0]), .B(n25305), .C(mtime_out[1]), 
         .Z(n25268)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4005_2_lut_rep_532_3_lut.init = 16'h8080;
    LUT4 i4012_2_lut_rep_499_3_lut_4_lut (.A(mtime_out[0]), .B(n25305), 
         .C(mtime_out[2]), .D(mtime_out[1]), .Z(n25235)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4012_2_lut_rep_499_3_lut_4_lut.init = 16'h8000;
    LUT4 increment_result_3__I_143_i3_4_lut (.A(mtime_out[2]), .B(\data_out_slice[2] ), 
         .C(n25269), .D(n25268), .Z(increment_result[2])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_143_i3_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_143_i2_4_lut (.A(mtime_out[1]), .B(\data_out_slice[1] ), 
         .C(n25269), .D(n25291), .Z(increment_result[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_143_i2_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_143_i1_4_lut (.A(mtime_out[0]), .B(\data_out_slice[0] ), 
         .C(n25269), .D(n25305), .Z(increment_result[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_143_i1_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_143_i4_4_lut (.A(mtime_out[3]), .B(n25277), 
         .C(n25269), .D(n25235), .Z(increment_result[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_143_i4_4_lut.init = 16'hc5ca;
    
endmodule
//
// Verilog Description of module tinyqv_decoder
//

module tinyqv_decoder (n24956, n25281, n26597, is_alu_imm_de, n25258, 
            n35, n26612, clk_c_enable_38, n3611, n24919, n25284, 
            n24894, n25227, n13701, is_ret_de, n22839, n25262, n25261, 
            n22398, n25288, n26598, n25287, n22384, n25265, n25267, 
            \instr[4] , n25264, n20820, n25266, n20650, n3597, \additional_mem_ops[2] , 
            n4031, n26, n3613, clk_c_enable_69, n23341, n25155, 
            n16, rst_reg_n, n22, n3589, n25153, n19, n3605, n25279, 
            n25231, n25278, n25247, n25249, n21978, \instr[12] , 
            n25256, n24939, n25290, n25260, n24940, \alu_op_3__N_901[2] , 
            n25234, \instr[26] , n25239, n22086, n25202, n25257, 
            is_store_de, n2438, n25214, \instr[30] , n3, n28, n25259, 
            n25212, n25241, n25243, n25209, n25216, n10, n24, 
            n25210, n12, n26596, n25211, n25189, n22202, n7955, 
            n26_adj_4, n22208, \instr[31] , n4532, \alu_op_3__N_1068[2] , 
            n22146, n22152, \instr[27] , n157, n25221, n13814, n25248, 
            \mem_op_de[2] , n25226, n2797, n25196, n22867, \instr[20] , 
            n25167, n21594, n26289, n27, n25245, n25244, is_branch_de, 
            n25208, n25338, n3615, n23255, \instr[16] , n2055, n27_adj_5, 
            n22470, n25207, n7734, n25203, n22286, \instr[25] , 
            n2799, n25166, n4533, n1655, n25289, n22976, mem_op_increment_reg_de, 
            n25014, n7375, n25225, n6647, n25222, n22_adj_6, n2240, 
            n15, n23899, alu_op_de, n4534, n4535, n15_adj_7, n23900, 
            n4531, n25228, n2437, is_alu_reg_de, n22226, n22232, 
            is_system_de, is_jalr_N_1101, is_jalr_de, n4547, n4542, 
            n4540, n3619, n23245, n8, n23379, is_load_de, n4543, 
            n20720, is_lui_N_1096, is_lui_de, n25190, n2430, is_auipc_de, 
            \mem_op_de[1] , n2242, \instr[17] , n2049, n2077, n22126, 
            n25182, n25177, n10_adj_8, n15_adj_9, n22254, n22238, 
            n22244, n25178, n25171, n25158, n3603, n21998, n22004, 
            n22178, n22184, n4, n22120, is_jal_de, n2658, n22132, 
            n22138, n25156, n22276, n22214, n22220) /* synthesis syn_module_defined=1 */ ;
    input n24956;
    input n25281;
    input n26597;
    output is_alu_imm_de;
    input n25258;
    input n35;
    input n26612;
    input clk_c_enable_38;
    output n3611;
    input n24919;
    input n25284;
    input n24894;
    output n25227;
    input n13701;
    output is_ret_de;
    input n22839;
    input n25262;
    input n25261;
    input n22398;
    input n25288;
    input n26598;
    input n25287;
    input n22384;
    input n25265;
    input n25267;
    input \instr[4] ;
    input n25264;
    input n20820;
    input n25266;
    input n20650;
    output n3597;
    input \additional_mem_ops[2] ;
    output n4031;
    input n26;
    output n3613;
    input clk_c_enable_69;
    output n23341;
    output n25155;
    input n16;
    input rst_reg_n;
    input n22;
    input n3589;
    output n25153;
    input n19;
    output n3605;
    input n25279;
    input n25231;
    input n25278;
    input n25247;
    input n25249;
    output n21978;
    input \instr[12] ;
    input n25256;
    output n24939;
    input n25290;
    output n25260;
    output n24940;
    input \alu_op_3__N_901[2] ;
    input n25234;
    input \instr[26] ;
    input n25239;
    output n22086;
    output n25202;
    input n25257;
    output is_store_de;
    output n2438;
    output n25214;
    input \instr[30] ;
    input n3;
    output n28;
    input n25259;
    output n25212;
    input n25241;
    input n25243;
    output n25209;
    output n25216;
    output n10;
    output n24;
    output n25210;
    output n12;
    output n26596;
    output n25211;
    output n25189;
    input n22202;
    input n7955;
    input n26_adj_4;
    output n22208;
    input \instr[31] ;
    output n4532;
    output \alu_op_3__N_1068[2] ;
    input n22146;
    output n22152;
    input \instr[27] ;
    output n157;
    output n25221;
    output n13814;
    input n25248;
    output \mem_op_de[2] ;
    output n25226;
    output n2797;
    output n25196;
    output n22867;
    input \instr[20] ;
    input n25167;
    output n21594;
    input n26289;
    output n27;
    input n25245;
    input n25244;
    output is_branch_de;
    output n25208;
    input n25338;
    input n3615;
    output n23255;
    input \instr[16] ;
    output n2055;
    input n27_adj_5;
    output n22470;
    output n25207;
    output n7734;
    output n25203;
    output n22286;
    input \instr[25] ;
    output n2799;
    output n25166;
    output n4533;
    input n1655;
    input n25289;
    output n22976;
    output mem_op_increment_reg_de;
    output n25014;
    output n7375;
    input n25225;
    output n6647;
    output n25222;
    input n22_adj_6;
    output n2240;
    output n15;
    input n23899;
    output [3:0]alu_op_de;
    output n4534;
    output n4535;
    input n15_adj_7;
    input n23900;
    output n4531;
    input n25228;
    output n2437;
    output is_alu_reg_de;
    input n22226;
    output n22232;
    output is_system_de;
    input is_jalr_N_1101;
    output is_jalr_de;
    output n4547;
    output n4542;
    output n4540;
    input n3619;
    output n23245;
    input n8;
    input n23379;
    output is_load_de;
    output n4543;
    output n20720;
    input is_lui_N_1096;
    output is_lui_de;
    output n25190;
    output n2430;
    output is_auipc_de;
    output \mem_op_de[1] ;
    input n2242;
    input \instr[17] ;
    input n2049;
    output n2077;
    input n22126;
    input n25182;
    input n25177;
    output n10_adj_8;
    input n15_adj_9;
    output n22254;
    input n22238;
    output n22244;
    input n25178;
    input n25171;
    output n25158;
    output n3603;
    input n21998;
    output n22004;
    input n22178;
    output n22184;
    input n4;
    output n22120;
    output is_jal_de;
    output n2658;
    input n22132;
    output n22138;
    output n25156;
    output n22276;
    input n22214;
    output n22220;
    
    
    wire n24957, n24958, n24922, n24921, n24918, n24920, n24893, 
        n25205, n24895, n22408, n22392, n25037, n25038, n25049;
    wire [2:0]additional_mem_ops_2__N_860;
    
    wire n26604, n7, n19_adj_2359, n25201, n25223, n14350, n6997, 
        n21444, n25193, n25199, n3_c, n21498, n14012, n25198;
    wire [3:0]alu_op_3__N_901;
    
    wire n26605, n25966;
    wire [3:0]n155;
    
    wire n30, n30_adj_2361, n30_adj_2362, n22476, imm_31__N_900, n25213, 
        n22588, alu_op_3__N_911, n21609, n26603, n20555, mem_op_2__N_1115, 
        n13744, n22580, n25961;
    wire [3:0]n328;
    
    wire n25224, n15_c, n15_adj_2364, n15_adj_2365, n25215, n6645, 
        n7369, n22516, n7373, n25050, n15_adj_2367;
    
    PFUMX i22412 (.BLUT(n24957), .ALUT(n24956), .C0(n25281), .Z(n24958));
    PFUMX i22386 (.BLUT(n24922), .ALUT(n24921), .C0(n26597), .Z(is_alu_imm_de));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n25258), .B(n35), .C(n26612), 
         .D(clk_c_enable_38), .Z(n3611)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h4000;
    PFUMX i22383 (.BLUT(n24919), .ALUT(n24918), .C0(n25284), .Z(n24920));
    PFUMX i22370 (.BLUT(n24894), .ALUT(n24893), .C0(n25205), .Z(n24895));
    LUT4 i1_4_lut (.A(n22408), .B(n22392), .C(n25227), .D(n13701), .Z(is_ret_de)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_290 (.A(n22839), .B(n25262), .C(n25261), .D(n22398), 
         .Z(n22408)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_290.init = 16'h0100;
    LUT4 i1_4_lut_adj_291 (.A(n25288), .B(n26598), .C(n25287), .D(n22384), 
         .Z(n22392)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_291.init = 16'h0100;
    LUT4 instr_3__bdd_3_lut (.A(n25265), .B(n25267), .C(\instr[4] ), .Z(n25037)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam instr_3__bdd_3_lut.init = 16'hf7f7;
    LUT4 instr_3__bdd_4_lut (.A(n25264), .B(n25265), .C(n25267), .D(\instr[4] ), 
         .Z(n25038)) /* synthesis lut_function=(A+(B (C+!(D))+!B (D))) */ ;
    defparam instr_3__bdd_4_lut.init = 16'hfbee;
    LUT4 n4_bdd_4_lut_22464 (.A(n20820), .B(n25266), .C(n25267), .D(\instr[4] ), 
         .Z(n25049)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam n4_bdd_4_lut_22464.init = 16'h0040;
    LUT4 i1_4_lut_adj_292 (.A(n25264), .B(n20650), .C(n25265), .D(n25266), 
         .Z(n3597)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_292.init = 16'h0400;
    LUT4 mux_55_i3_4_lut_4_lut (.A(n25258), .B(clk_c_enable_38), .C(additional_mem_ops_2__N_860[2]), 
         .D(\additional_mem_ops[2] ), .Z(n4031)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;
    defparam mux_55_i3_4_lut_4_lut.init = 16'h7340;
    LUT4 i21913_2_lut_3_lut_4_lut_4_lut (.A(n25258), .B(n26), .C(n3613), 
         .D(clk_c_enable_69), .Z(n23341)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i21913_2_lut_3_lut_4_lut_4_lut.init = 16'hfbff;
    LUT4 i1_2_lut_rep_419_3_lut_4_lut_4_lut (.A(n25258), .B(n26), .C(n26612), 
         .D(clk_c_enable_38), .Z(n25155)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_rep_419_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_293 (.A(n25258), .B(n16), .C(rst_reg_n), 
         .D(clk_c_enable_38), .Z(n3613)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_293.init = 16'h4000;
    LUT4 i6973_2_lut_rep_417_3_lut_4_lut_4_lut (.A(n25258), .B(n22), .C(n3589), 
         .D(clk_c_enable_69), .Z(n25153)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i6973_2_lut_rep_417_3_lut_4_lut_4_lut.init = 16'hfbff;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_294 (.A(n25258), .B(n19), .C(rst_reg_n), 
         .D(clk_c_enable_38), .Z(n3605)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_294.init = 16'h4000;
    LUT4 i22786_then_4_lut (.A(n25258), .B(n25281), .C(n26598), .D(n25279), 
         .Z(n26604)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam i22786_then_4_lut.init = 16'h4470;
    LUT4 instr_1__I_0_139_i7_4_lut (.A(n25231), .B(n25278), .C(n25284), 
         .D(n25247), .Z(n7)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam instr_1__I_0_139_i7_4_lut.init = 16'h0a3a;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n25258), .B(n25249), .C(rst_reg_n), 
         .D(n25284), .Z(n21978)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h1000;
    LUT4 n928_bdd_3_lut_22399_4_lut (.A(\instr[12] ), .B(n25256), .C(n25279), 
         .D(n26598), .Z(n24939)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam n928_bdd_3_lut_22399_4_lut.init = 16'h0002;
    LUT4 n928_bdd_3_lut_4_lut (.A(n25290), .B(n25260), .C(n25279), .D(n26598), 
         .Z(n24940)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(182[25:44])
    defparam n928_bdd_3_lut_4_lut.init = 16'h2000;
    LUT4 i12128_4_lut (.A(n19_adj_2359), .B(n25201), .C(n26597), .D(n25223), 
         .Z(n14350)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i12128_4_lut.init = 16'hcac0;
    LUT4 i1_3_lut (.A(n6997), .B(\alu_op_3__N_901[2] ), .C(n26597), .Z(n21444)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i25_2_lut_rep_457_3_lut_4_lut (.A(\instr[4] ), .B(n25234), .C(\instr[26] ), 
         .D(n25239), .Z(n25193)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(67[27:51])
    defparam i25_2_lut_rep_457_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_4_lut_adj_295 (.A(n25199), .B(n3_c), .C(n25287), .D(n25205), 
         .Z(n21498)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i1_4_lut_adj_295.init = 16'h5044;
    LUT4 i1_3_lut_rep_491 (.A(n25278), .B(n25260), .C(n25290), .Z(n25227)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_3_lut_rep_491.init = 16'hfefe;
    LUT4 i1_2_lut_2_lut_4_lut (.A(n25278), .B(n25260), .C(n25290), .D(n25258), 
         .Z(n22086)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_2_lut_4_lut.init = 16'h00fe;
    LUT4 is_store_I_0_4_lut (.A(n14012), .B(n25202), .C(n25258), .D(n25257), 
         .Z(is_store_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam is_store_I_0_4_lut.init = 16'h3a30;
    LUT4 i11792_4_lut (.A(n25281), .B(n26598), .C(n25279), .D(n25278), 
         .Z(n14012)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i11792_4_lut.init = 16'hcdcc;
    LUT4 mux_1484_i9_3_lut_4_lut_4_lut (.A(\instr[4] ), .B(n25265), .C(n25284), 
         .D(n25264), .Z(n2438)) /* synthesis lut_function=(A (B+((D)+!C))+!A (C (D))) */ ;
    defparam mux_1484_i9_3_lut_4_lut_4_lut.init = 16'hfa8a;
    LUT4 i21801_2_lut_rep_478_3_lut (.A(\instr[4] ), .B(n25265), .C(n25264), 
         .Z(n25214)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i21801_2_lut_rep_478_3_lut.init = 16'h0808;
    LUT4 mux_29_i2_4_lut (.A(n26598), .B(n25193), .C(n25198), .D(n25279), 
         .Z(alu_op_3__N_901[1])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[18] 85[91])
    defparam mux_29_i2_4_lut.init = 16'hfaca;
    LUT4 i4441_4_lut (.A(\instr[12] ), .B(n25279), .C(n25193), .D(n25198), 
         .Z(alu_op_3__N_901[0])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[18] 85[91])
    defparam i4441_4_lut.init = 16'hcacc;
    LUT4 n25965_bdd_3_lut_4_lut (.A(n26598), .B(n25258), .C(n25284), .D(n26605), 
         .Z(n25966)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam n25965_bdd_3_lut_4_lut.init = 16'h2f20;
    LUT4 i11664_4_lut (.A(\instr[30] ), .B(n25193), .C(n25267), .D(n3), 
         .Z(n155[3])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(85[18:91])
    defparam i11664_4_lut.init = 16'hecee;
    LUT4 i12040_2_lut_3_lut_4_lut (.A(n26598), .B(n26597), .C(n25279), 
         .D(n25284), .Z(n30)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i12040_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i21811_2_lut_rep_487_3_lut (.A(n26598), .B(n26597), .C(n25284), 
         .Z(n25223)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i21811_2_lut_rep_487_3_lut.init = 16'h1010;
    LUT4 i49_3_lut_3_lut (.A(n26598), .B(n26597), .C(n25281), .Z(n28)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i49_3_lut_3_lut.init = 16'h1c1c;
    LUT4 i12038_2_lut_3_lut_4_lut (.A(n26598), .B(n26597), .C(n25290), 
         .D(n25259), .Z(n30_adj_2361)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i12038_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i12036_2_lut_3_lut_4_lut (.A(n26598), .B(n26597), .C(n25288), 
         .D(n25259), .Z(n30_adj_2362)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i12036_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i20704_3_lut_rep_476_4_lut (.A(n25264), .B(n25265), .C(\instr[4] ), 
         .D(n25262), .Z(n25212)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20704_3_lut_rep_476_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut (.A(n25264), .B(n25265), .C(\instr[12] ), .Z(n22476)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_466_3_lut_4_lut (.A(n25267), .B(n25266), .C(n25239), 
         .D(\instr[4] ), .Z(n25202)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(67[27:51])
    defparam i1_2_lut_rep_466_3_lut_4_lut.init = 16'hfffd;
    LUT4 instr_6__I_0_127_i10_2_lut_3_lut_4_lut (.A(n25267), .B(n25266), 
         .C(n25241), .D(\instr[4] ), .Z(imm_31__N_900)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(67[27:51])
    defparam instr_6__I_0_127_i10_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i21747_2_lut_rep_465_3_lut_4_lut (.A(n25267), .B(n25266), .C(n25239), 
         .D(\instr[4] ), .Z(n25201)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(67[27:51])
    defparam i21747_2_lut_rep_465_3_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_477_3_lut (.A(n25267), .B(n25266), .C(\instr[4] ), 
         .Z(n25213)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(67[27:51])
    defparam i1_2_lut_rep_477_3_lut.init = 16'hfdfd;
    LUT4 instr_6__I_0_157_i9_2_lut_rep_462_3_lut_4_lut (.A(n25265), .B(n25264), 
         .C(n25243), .D(\instr[4] ), .Z(n25198)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(72[27:51])
    defparam instr_6__I_0_157_i9_2_lut_rep_462_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_3_lut_4_lut (.A(n25265), .B(n25264), .C(\instr[4] ), .D(n25281), 
         .Z(n22588)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(72[27:51])
    defparam i1_3_lut_4_lut.init = 16'h1000;
    LUT4 instr_6__I_0_130_i10_2_lut_3_lut_4_lut (.A(n25265), .B(n25264), 
         .C(n25243), .D(\instr[4] ), .Z(alu_op_3__N_911)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam instr_6__I_0_130_i10_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_3_lut_rep_473_4_lut (.A(n25265), .B(n25264), .C(n25266), .D(\instr[4] ), 
         .Z(n25209)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i1_3_lut_rep_473_4_lut.init = 16'hfdff;
    LUT4 i1_2_lut_rep_480_3_lut (.A(n25267), .B(n25266), .C(\instr[4] ), 
         .Z(n25216)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(218[25] 223[32])
    defparam i1_2_lut_rep_480_3_lut.init = 16'hf7f7;
    LUT4 n20725_bdd_2_lut_3_lut (.A(n26598), .B(n25284), .C(n25279), .Z(n24957)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n20725_bdd_2_lut_3_lut.init = 16'h7070;
    LUT4 i2_2_lut_3_lut (.A(n26598), .B(n25284), .C(n25279), .Z(n10)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n26598), .B(n25284), .C(n25279), 
         .D(n25258), .Z(n21609)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i22786_else_4_lut (.A(n25258), .B(n25281), .C(n26598), .D(n25279), 
         .Z(n26603)) /* synthesis lut_function=(!(A (B+(D))+!A !(B (C+(D))+!B !(D)))) */ ;
    defparam i22786_else_4_lut.init = 16'h4473;
    LUT4 i37_3_lut_3_lut (.A(n26598), .B(n25284), .C(n25279), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;
    defparam i37_3_lut_3_lut.init = 16'h7a7a;
    LUT4 i2_2_lut_3_lut_3_lut_4_lut (.A(n26598), .B(n25279), .C(n25210), 
         .D(n25258), .Z(n12)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i2_2_lut_3_lut_3_lut_4_lut.init = 16'hf0fe;
    LUT4 is_alu_imm_N_1098_bdd_2_lut_22385_3_lut_4_lut (.A(n26598), .B(n25279), 
         .C(n25256), .D(\instr[12] ), .Z(n24918)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam is_alu_imm_N_1098_bdd_2_lut_22385_3_lut_4_lut.init = 16'h1110;
    LUT4 is_alu_imm_N_1098_bdd_2_lut_3_lut (.A(n26598), .B(n25279), .C(n25284), 
         .Z(n24922)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam is_alu_imm_N_1098_bdd_2_lut_3_lut.init = 16'h0101;
    LUT4 i169_2_lut_rep_704 (.A(n25281), .B(n26597), .C(n25279), .Z(n26596)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i169_2_lut_rep_704.init = 16'h7070;
    LUT4 i21827_2_lut_3_lut (.A(n26598), .B(n25279), .C(n25284), .Z(n20555)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i21827_2_lut_3_lut.init = 16'h0101;
    LUT4 i21749_2_lut_rep_475_3_lut_4_lut (.A(n26598), .B(n25279), .C(n25284), 
         .D(n26597), .Z(n25211)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i21749_2_lut_rep_475_3_lut_4_lut.init = 16'h0001;
    LUT4 i528_4_lut_rep_453 (.A(n25279), .B(mem_op_2__N_1115), .C(n13744), 
         .D(\instr[12] ), .Z(n25189)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(93[13] 98[16])
    defparam i528_4_lut_rep_453.init = 16'h3b33;
    LUT4 i1_2_lut_4_lut (.A(n25279), .B(mem_op_2__N_1115), .C(n13744), 
         .D(\instr[12] ), .Z(n3_c)) /* synthesis lut_function=(A (B (C (D)))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(93[13] 98[16])
    defparam i1_2_lut_4_lut.init = 16'hc400;
    LUT4 i1_4_lut_4_lut (.A(n25258), .B(n22202), .C(n7955), .D(n26_adj_4), 
         .Z(n22208)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h0400;
    LUT4 mux_2749_i16_3_lut_3_lut (.A(n25209), .B(n25284), .C(\instr[31] ), 
         .Z(n4532)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2749_i16_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n25267), .B(n25266), .C(n25256), .D(\instr[12] ), 
         .Z(\alu_op_3__N_1068[2] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    PFUMX i23145 (.BLUT(n26603), .ALUT(n26604), .C0(mem_op_2__N_1115), 
          .Z(n26605));
    LUT4 i1_2_lut_3_lut_adj_296 (.A(n25267), .B(n25266), .C(\instr[12] ), 
         .Z(n22580)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam i1_2_lut_3_lut_adj_296.init = 16'hfefe;
    LUT4 i1_4_lut_4_lut_adj_297 (.A(n25258), .B(n22146), .C(n7955), .D(n26_adj_4), 
         .Z(n22152)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_297.init = 16'h0400;
    LUT4 mux_28_i3_3_lut_4_lut (.A(\instr[26] ), .B(n25201), .C(\instr[27] ), 
         .D(n26598), .Z(n157)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[22:45])
    defparam mux_28_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 n25283_bdd_4_lut_22957_4_lut (.A(n25281), .B(n26597), .C(n25279), 
         .D(mem_op_2__N_1115), .Z(n25961)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam n25283_bdd_4_lut_22957_4_lut.init = 16'h808a;
    LUT4 i532_2_lut_rep_485_3_lut (.A(n25287), .B(n25278), .C(\instr[12] ), 
         .Z(n25221)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i532_2_lut_rep_485_3_lut.init = 16'h8080;
    LUT4 i11595_2_lut_3_lut_4_lut (.A(n25287), .B(n25278), .C(n26597), 
         .D(\instr[12] ), .Z(n13814)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i11595_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_298 (.A(n25199), .B(n24895), .C(n25249), .D(n25248), 
         .Z(\mem_op_de[2] )) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_298.init = 16'h0004;
    LUT4 i11841_3_lut_3_lut_4_lut (.A(n25287), .B(n25278), .C(n328[0]), 
         .D(n25224), .Z(n15_c)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;
    defparam i11841_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 i12042_4_lut_4_lut_4_lut (.A(n25287), .B(n25278), .C(n328[1]), 
         .D(n25224), .Z(n15_adj_2364)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!B))) */ ;
    defparam i12042_4_lut_4_lut_4_lut.init = 16'h00c4;
    LUT4 i11902_2_lut_3_lut_4_lut (.A(n25287), .B(n25278), .C(n25224), 
         .D(\instr[12] ), .Z(n15_adj_2365)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i11902_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_490_3_lut_4_lut (.A(n25284), .B(n26597), .C(n25279), 
         .D(n26598), .Z(n25226)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i1_2_lut_rep_490_3_lut_4_lut.init = 16'h2000;
    LUT4 i5264_3_lut_4_lut (.A(n25281), .B(n26597), .C(\instr[27] ), .D(n25290), 
         .Z(n2797)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5264_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_460_2_lut_3_lut (.A(n25281), .B(n26597), .C(n26612), 
         .Z(n25196)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_2_lut_rep_460_2_lut_3_lut.init = 16'h7070;
    LUT4 i20655_2_lut_3_lut (.A(n25281), .B(n26597), .C(n26598), .Z(n22867)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i20655_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i4685_2_lut_rep_463_2_lut_3_lut_4_lut (.A(n25281), .B(n26597), 
         .C(n25279), .D(n26598), .Z(n25199)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i4685_2_lut_rep_463_2_lut_3_lut_4_lut.init = 16'h7770;
    LUT4 i1_3_lut_3_lut_4_lut (.A(n25281), .B(n26597), .C(\instr[20] ), 
         .D(n25167), .Z(n21594)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_adj_299 (.A(n25281), .B(n26597), .C(n26289), .Z(n27)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_2_lut_3_lut_adj_299.init = 16'hf8f8;
    LUT4 is_branch_I_0_4_lut (.A(n25245), .B(n25198), .C(n25258), .D(n25244), 
         .Z(is_branch_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam is_branch_I_0_4_lut.init = 16'h3a30;
    LUT4 i1_2_lut_rep_472_3_lut (.A(n25281), .B(n26597), .C(n26612), .Z(n25208)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_2_lut_rep_472_3_lut.init = 16'h8080;
    LUT4 i21941_3_lut_4_lut (.A(n25281), .B(n26597), .C(n25338), .D(n3615), 
         .Z(n23255)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i21941_3_lut_4_lut.init = 16'hff08;
    LUT4 i11609_2_lut_3_lut (.A(n25281), .B(n26597), .C(\instr[16] ), 
         .Z(n2055)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i11609_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_3_lut_4_lut_adj_300 (.A(n25281), .B(n26597), .C(n27_adj_5), 
         .D(n25284), .Z(n22470)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !((D)+!C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_3_lut_4_lut_adj_300.init = 16'h88f8;
    LUT4 i12002_2_lut_rep_471_3_lut (.A(n25281), .B(n26597), .C(\instr[31] ), 
         .Z(n25207)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i12002_2_lut_rep_471_3_lut.init = 16'h8080;
    LUT4 i5503_3_lut_4_lut (.A(n25281), .B(n26597), .C(n3615), .D(n25209), 
         .Z(n7734)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5503_3_lut_4_lut.init = 16'hf808;
    LUT4 i168_2_lut_rep_467_2_lut_3_lut (.A(n25281), .B(n26597), .C(n26598), 
         .Z(n25203)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i168_2_lut_rep_467_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut_adj_301 (.A(n25281), .B(n26597), .C(n26612), 
         .D(n7955), .Z(n22286)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_2_lut_3_lut_3_lut_4_lut_adj_301.init = 16'h0070;
    LUT4 i167_2_lut_rep_469_2_lut_3_lut (.A(n25281), .B(n26597), .C(n25284), 
         .Z(n25205)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i167_2_lut_rep_469_2_lut_3_lut.init = 16'h7070;
    LUT4 n24920_bdd_3_lut_4_lut (.A(n25239), .B(n25215), .C(n25281), .D(n24920), 
         .Z(n24921)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;
    defparam n24920_bdd_3_lut_4_lut.init = 16'h1f10;
    LUT4 i5260_3_lut_4_lut (.A(n25281), .B(n26597), .C(\instr[25] ), .D(\instr[12] ), 
         .Z(n2799)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5260_3_lut_4_lut.init = 16'hf780;
    LUT4 i5256_rep_430_4_lut (.A(n25281), .B(n26597), .C(n25167), .D(n3597), 
         .Z(n25166)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5256_rep_430_4_lut.init = 16'h08f8;
    LUT4 mux_2749_i15_3_lut_3_lut (.A(n25209), .B(n26598), .C(\instr[31] ), 
         .Z(n4533)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2749_i15_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_1013_i11_rep_97_3_lut_3_lut_4_lut (.A(n25281), .B(n26597), 
         .C(n1655), .D(n25289), .Z(n22976)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam mux_1013_i11_rep_97_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 i11538_2_lut_2_lut_3_lut (.A(n25281), .B(n26597), .C(mem_op_2__N_1115), 
         .Z(mem_op_increment_reg_de)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i11538_2_lut_2_lut_3_lut.init = 16'hf7f7;
    LUT4 n15_bdd_3_lut_3_lut (.A(n26597), .B(n25284), .C(n26598), .Z(n25014)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam n15_bdd_3_lut_3_lut.init = 16'h1414;
    LUT4 i4446_4_lut_4_lut (.A(n26597), .B(n6997), .C(n20555), .D(alu_op_3__N_901[0]), 
         .Z(n6645)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i4446_4_lut_4_lut.init = 16'hd850;
    LUT4 i5139_4_lut_4_lut (.A(n26597), .B(n6997), .C(n30), .D(alu_op_3__N_901[1]), 
         .Z(n7369)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5139_4_lut_4_lut.init = 16'hd850;
    LUT4 i21596_3_lut_4_lut_4_lut (.A(n26597), .B(n30_adj_2361), .C(n25189), 
         .D(n26598), .Z(n7375)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i21596_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 i5143_4_lut_4_lut (.A(n26597), .B(n155[3]), .C(n30), .D(n22516), 
         .Z(n7373)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5143_4_lut_4_lut.init = 16'hd850;
    LUT4 i1_3_lut_rep_488_4_lut_4_lut (.A(n26597), .B(n25284), .C(n25279), 
         .D(n26598), .Z(n25224)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_3_lut_rep_488_4_lut_4_lut.init = 16'hfff7;
    LUT4 i4448_4_lut_4_lut (.A(n26597), .B(n25225), .C(n25289), .D(n25189), 
         .Z(n6647)) /* synthesis lut_function=(A (D)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i4448_4_lut_4_lut.init = 16'hea40;
    LUT4 i1_3_lut_rep_524 (.A(n25289), .B(n25287), .C(n25288), .Z(n25260)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(182[25:44])
    defparam i1_3_lut_rep_524.init = 16'hfefe;
    LUT4 i1_2_lut_rep_486_4_lut (.A(n25289), .B(n25287), .C(n25288), .D(n25290), 
         .Z(n25222)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(182[25:44])
    defparam i1_2_lut_rep_486_4_lut.init = 16'hfeff;
    LUT4 i1_3_lut_rep_474_4_lut (.A(\instr[4] ), .B(n25265), .C(n25264), 
         .D(n25262), .Z(n25210)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_rep_474_4_lut.init = 16'hfffe;
    LUT4 n4_bdd_4_lut_4_lut_4_lut (.A(n25281), .B(n25279), .C(n26597), 
         .D(n26598), .Z(n25050)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam n4_bdd_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_479_3_lut (.A(n25267), .B(n25266), .C(\instr[4] ), 
         .Z(n25215)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(65[27:51])
    defparam i1_2_lut_rep_479_3_lut.init = 16'hefef;
    LUT4 i12039_4_lut_4_lut (.A(n25224), .B(n22580), .C(n25287), .D(n25278), 
         .Z(n15_adj_2367)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C)))) */ ;
    defparam i12039_4_lut_4_lut.init = 16'h1050;
    LUT4 i2_2_lut_3_lut_4_lut_4_lut (.A(n25258), .B(n22_adj_6), .C(n26612), 
         .D(clk_c_enable_38), .Z(n2240)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i2_2_lut_3_lut_4_lut_4_lut.init = 16'h4000;
    PFUMX instr_1__I_0_133_Mux_0_i15 (.BLUT(n21498), .ALUT(n21609), .C0(n25248), 
          .Z(n15)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    PFUMX i5140 (.BLUT(n15_adj_2364), .ALUT(n7369), .C0(n23899), .Z(alu_op_de[1]));
    PFUMX i4447 (.BLUT(n15_c), .ALUT(n6645), .C0(n23899), .Z(alu_op_de[0]));
    LUT4 mux_2749_i14_3_lut_3_lut (.A(n25209), .B(n25279), .C(\instr[31] ), 
         .Z(n4534)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2749_i14_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_2749_i13_3_lut_3_lut (.A(n25209), .B(\instr[12] ), .C(\instr[31] ), 
         .Z(n4535)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2749_i13_3_lut_3_lut.init = 16'he4e4;
    PFUMX i5142 (.BLUT(n15_adj_7), .ALUT(n21444), .C0(n23900), .Z(alu_op_de[2]));
    LUT4 mux_2749_i17_3_lut_3_lut (.A(n25209), .B(\instr[16] ), .C(\instr[31] ), 
         .Z(n4531)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam mux_2749_i17_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_1484_i11_rep_72_3_lut_4_lut (.A(n25264), .B(n25228), .C(n25284), 
         .D(\instr[12] ), .Z(n2437)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(205[25] 214[32])
    defparam mux_1484_i11_rep_72_3_lut_4_lut.init = 16'hefe0;
    PFUMX i5144 (.BLUT(n15_adj_2367), .ALUT(n7373), .C0(n23900), .Z(alu_op_de[3]));
    PFUMX i12129 (.BLUT(n15_adj_2365), .ALUT(n14350), .C0(n23899), .Z(is_alu_reg_de));
    LUT4 i1_4_lut_4_lut_adj_302 (.A(n25258), .B(n22226), .C(n7955), .D(n26_adj_4), 
         .Z(n22232)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_302.init = 16'h0400;
    LUT4 i24_4_lut (.A(n24958), .B(n22588), .C(n26597), .D(n25243), 
         .Z(is_system_de)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i24_4_lut.init = 16'hca0a;
    PFUMX is_jalr_I_0 (.BLUT(is_jalr_N_1101), .ALUT(alu_op_3__N_911), .C0(n25258), 
          .Z(is_jalr_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 i11611_2_lut_4_lut (.A(\instr[4] ), .B(n25241), .C(n25266), .D(n25289), 
         .Z(n4547)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i11611_2_lut_4_lut.init = 16'hfd00;
    LUT4 i11887_2_lut_4_lut (.A(\instr[4] ), .B(n25241), .C(n25266), .D(\instr[25] ), 
         .Z(n4542)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i11887_2_lut_4_lut.init = 16'hfd00;
    LUT4 i11889_2_lut_4_lut (.A(\instr[4] ), .B(n25241), .C(n25266), .D(\instr[27] ), 
         .Z(n4540)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i11889_2_lut_4_lut.init = 16'hfd00;
    LUT4 i21943_2_lut_3_lut_4_lut_4_lut (.A(n25258), .B(n26), .C(n3619), 
         .D(clk_c_enable_69), .Z(n23245)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i21943_2_lut_3_lut_4_lut_4_lut.init = 16'hfbff;
    PFUMX i21 (.BLUT(n7), .ALUT(n8), .C0(n23379), .Z(is_load_de));
    LUT4 i11886_2_lut_4_lut (.A(\instr[4] ), .B(n25241), .C(n25266), .D(n25278), 
         .Z(n4543)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;
    defparam i11886_2_lut_4_lut.init = 16'hfd00;
    LUT4 i11808_2_lut_4_lut (.A(n25261), .B(n25262), .C(n25264), .D(n25279), 
         .Z(n19_adj_2359)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(72[27:51])
    defparam i11808_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_303 (.A(n25262), .B(n25239), .C(\instr[4] ), 
         .D(n25281), .Z(n20720)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_4_lut_adj_303.init = 16'h0100;
    LUT4 i11525_2_lut_3_lut_4_lut (.A(\instr[4] ), .B(n25234), .C(n25210), 
         .D(n25239), .Z(n13744)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i11525_2_lut_3_lut_4_lut.init = 16'hf0e0;
    PFUMX is_lui_I_0 (.BLUT(is_lui_N_1096), .ALUT(imm_31__N_900), .C0(n25258), 
          .Z(is_lui_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 i11702_2_lut_rep_454_3_lut_4_lut (.A(\instr[4] ), .B(n25234), .C(n25209), 
         .D(n25239), .Z(n25190)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i11702_2_lut_rep_454_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_61_i2_3_lut_4_lut (.A(n25264), .B(n25228), .C(\instr[12] ), 
         .D(n25266), .Z(n328[1])) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_61_i2_3_lut_4_lut.init = 16'hbfb0;
    LUT4 mux_61_i1_3_lut_4_lut (.A(n25264), .B(n25228), .C(\instr[12] ), 
         .D(n25243), .Z(n328[0])) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_61_i1_3_lut_4_lut.init = 16'hbfb0;
    LUT4 mux_1484_i17_3_lut_4_lut (.A(n25264), .B(n25228), .C(n25284), 
         .D(\instr[12] ), .Z(n2430)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_1484_i17_3_lut_4_lut.init = 16'h4f40;
    LUT4 i1_3_lut_4_lut_adj_304 (.A(\instr[4] ), .B(n25262), .C(n25258), 
         .D(n25241), .Z(is_auipc_de)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(65[27:51])
    defparam i1_3_lut_4_lut_adj_304.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_305 (.A(\instr[4] ), .B(n25243), .C(n6997), 
         .D(n25239), .Z(n22516)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(70[27:51])
    defparam i1_2_lut_3_lut_4_lut_adj_305.init = 16'hf0b0;
    PFUMX i22788 (.BLUT(n25966), .ALUT(n25961), .C0(n26597), .Z(\mem_op_de[1] ));
    LUT4 mux_1313_i3_4_lut_4_lut (.A(n25258), .B(n2242), .C(\instr[17] ), 
         .D(n2049), .Z(n2077)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;
    defparam mux_1313_i3_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i2_2_lut_3_lut_4_lut_4_lut_adj_306 (.A(n25258), .B(n22126), .C(n25182), 
         .D(n25177), .Z(n10_adj_8)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i2_2_lut_3_lut_4_lut_4_lut_adj_306.init = 16'h1110;
    PFUMX instr_1__I_0_138_Mux_2_i31 (.BLUT(n15_adj_9), .ALUT(n30_adj_2362), 
          .C0(n23900), .Z(additional_mem_ops_2__N_860[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 i1_4_lut_4_lut_adj_307 (.A(n25258), .B(n26612), .C(\instr[12] ), 
         .D(n7955), .Z(n22254)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_307.init = 16'h0040;
    LUT4 i1_4_lut_adj_308 (.A(n25279), .B(n25213), .C(n26598), .D(n22476), 
         .Z(mem_op_2__N_1115)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_308.init = 16'hffdf;
    LUT4 i1_4_lut_4_lut_adj_309 (.A(n25258), .B(n22238), .C(n7955), .D(n26_adj_4), 
         .Z(n22244)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_309.init = 16'h0400;
    LUT4 additional_mem_ops_2__N_863_0__bdd_3_lut (.A(n25278), .B(n25287), 
         .C(n25266), .Z(n24893)) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam additional_mem_ops_2__N_863_0__bdd_3_lut.init = 16'h1515;
    LUT4 i1_2_lut_rep_422_3_lut_4_lut_4_lut (.A(n25258), .B(n26612), .C(n25178), 
         .D(n25171), .Z(n25158)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_422_3_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_310 (.A(n25258), .B(n26_adj_4), 
         .C(n26612), .D(clk_c_enable_38), .Z(n3603)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_310.init = 16'h4000;
    LUT4 i1_4_lut_4_lut_adj_311 (.A(n25258), .B(n21998), .C(n7955), .D(n19), 
         .Z(n22004)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_311.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_312 (.A(n25258), .B(n22178), .C(n7955), .D(n26_adj_4), 
         .Z(n22184)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_312.init = 16'h0400;
    LUT4 i1_3_lut_4_lut_4_lut_adj_313 (.A(n25258), .B(n7955), .C(n4), 
         .D(rst_reg_n), .Z(n22120)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_313.init = 16'h1000;
    PFUMX i22465 (.BLUT(n25050), .ALUT(n25049), .C0(n25258), .Z(is_jal_de));
    PFUMX i22456 (.BLUT(n25038), .ALUT(n25037), .C0(n25266), .Z(n6997));
    LUT4 i11933_2_lut_3_lut_4_lut_4_lut (.A(n25258), .B(n22), .C(n3589), 
         .D(clk_c_enable_69), .Z(n2658)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i11933_2_lut_3_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_314 (.A(n25258), .B(n22132), .C(n7955), .D(n26_adj_4), 
         .Z(n22138)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_314.init = 16'h0400;
    LUT4 i1_2_lut_rep_420_3_lut_4_lut_4_lut (.A(n25258), .B(n22), .C(n26612), 
         .D(clk_c_enable_38), .Z(n25156)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_rep_420_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i1_3_lut_4_lut_4_lut_adj_315 (.A(n25258), .B(n25248), .C(n25249), 
         .D(n25284), .Z(n22276)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_315.init = 16'h1000;
    LUT4 i1_4_lut_4_lut_adj_316 (.A(n25258), .B(n22214), .C(n7955), .D(n26_adj_4), 
         .Z(n22220)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_316.init = 16'h0400;
    
endmodule
//
// Verilog Description of module tinyqv_core
//

module tinyqv_core (clk_c, n25273, clk_c_enable_27, \mie[0] , n92, 
            instr_retired, instr_complete_N_1378, n25424, cmp, \imm[11] , 
            instr_complete_N_1382, \next_fsm_state_3__N_2230[3] , cy, 
            mstatus_mte, clk_c_enable_111, mstatus_mpie, clk_c_enable_170, 
            \addr_out[11] , \addr_out[12] , \addr_out[13] , \addr_out[14] , 
            \addr_out[15] , counter_hi, \addr_out[16] , \addr_out[17] , 
            \addr_out[18] , \addr_out[19] , n25372, n25365, \addr_out[20] , 
            \addr_out[21] , \addr_out[22] , \imm[6] , \addr_out[23] , 
            \alu_op[1] , debug_instr_valid, is_system, \alu_op[0] , 
            n25310, n5, clk_c_enable_205, n25344, \imm[1] , cycle_count_wide, 
            \imm[0] , \next_pc_for_core[22] , \next_pc_for_core[18] , 
            \mie[8] , data_rs1, n25179, n25175, n22208, n25178, 
            n21248, n22098, n3615, timer_interrupt, n26608, n22172, 
            n2037, n22258, n2835, n22867, n7955, n24916, n22272, 
            n22152, n21113, \alu_op_in[2] , n25430, n22254, n26, 
            n24486, n22184, n21260, n22244, n21230, n22138, n21121, 
            n22004, n25182, n25177, n22008, n22324, n21303, n22298, 
            n21297, n22120, n2236, n22220, n21242, n25216, n21910, 
            n21916, n22933, n22852, n22086, n25191, n22092, n22276, 
            n12, n22282, n21898, n21212, n22232, n21236, n23322, 
            \cycle[0] , \addr_out[3] , n11558, \ui_in_sync[1] , n1092, 
            n25343, n26610, any_additional_mem_ops, clk_c_enable_206, 
            n25349, interrupt_core, clk_c_enable_209, is_load, n54, 
            n20739, clk_c_enable_393, n21402, n4455, n1768, pc_2__N_663, 
            load_done, n6638, n1767, \instr_write_offset_3__N_665[0] , 
            n1766, \instr_write_offset_3__N_665[1] , n25181, mem_op, 
            n5031, \addr_out[6] , debug_rd, debug_rd_3__N_1306, \addr_out[7] , 
            n25369, \imm[2] , n25410, accum, d_3__N_1599, \imm[7] , 
            \imm[8] , \imm[10] , \imm[9] , n24938, \debug_branch_N_181[0] , 
            \addr_out[4] , \mul_out[1] , n25421, data_rs2, \debug_rd_3__N_136[28] , 
            alu_b_in, n25316, \addr_out[8] , \mul_out[3] , \mcause[2] , 
            \alu_b_in[1] , \alu_a_in[1] , n5047, \alu_a_in[0] , n6657, 
            was_early_branch, instr_fetch_restart_N_678, data_out_3__N_1116, 
            \data_out_slice[1] , n22354, mstatus_mie, n21750, n22028, 
            n22030, n25180, rst_reg_n, n14111, n20807, \next_pc_offset[3] , 
            n21864, n25422, n5_adj_1, clk_c_enable_54, \addr_out[10] , 
            \debug_branch_N_173[28] , n22941, \addr_out[0] , n25411, 
            n25333, n25359, \next_pc_for_core[15] , \next_pc_for_core[11] , 
            load_top_bit, \debug_branch_N_181[3] , n25352, cy_adj_2, 
            data_ready_sync, n25197, data_ready_core, n24186, cy_adj_3, 
            \addr_out[5] , \instrret_count[0] , n23011, n25408, \debug_branch_N_173[30] , 
            n25402, n25350, clk_c_enable_336, n18, clk_c_enable_197, 
            n23898, n23897, n23896, n23895, n23894, \imm[4] , \addr_out[26] , 
            n25307, \addr_out[25] , \addr_out[24] , \alu_op[3] , is_alu_imm, 
            is_alu_reg, is_auipc, \debug_branch_N_173[29] , is_jal, 
            n25426, \debug_rd_3__N_136[29] , n4996, n24264, is_jalr, 
            n25412, n23395, is_lui, is_store, \data_out_slice[0] , 
            \debug_branch_N_571[29] , \timer_data[1] , is_timer_addr, 
            \imm[5] , \imm[3] , is_branch, n25277, \data_rs1[3] , 
            n23111, n25375, n22798, n25387, \debug_rd_3__N_136[31] , 
            \tmp_data_in_3__N_1245[3] , n25319, \debug_rd_3__N_136[30] , 
            \addr_out[9] , \debug_branch_N_173[31] , n25301, \debug_rd_3__N_1298[0] , 
            n25293, n25282, \mtimecmp[7] , mtimecmp_3__N_1666, \data_out_slice[2] , 
            n24932, \debug_branch_N_181[2] , no_write_in_progress, n25348, 
            n25326, n23069, \addr_out[1] , n22944, \debug_branch_N_571[31] , 
            n23073, \debug_branch_N_177[31] , \mul_out[2] , n23067, 
            \debug_branch_N_177[29] , \next_pc_for_core[14] , \next_pc_for_core[10] , 
            n66, n12257, \addr_offset[2] , n701, n23070, \debug_branch_N_177[30] , 
            n25341, n25271, n22939, n23012, n25475, \csr_read_3__N_1170[3] , 
            \next_accum[6] , \next_accum[7] , \next_accum[8] , \next_accum[9] , 
            \next_accum[10] , \next_accum[11] , \next_accum[12] , \next_accum[13] , 
            \next_accum[14] , \next_accum[15] , GND_net, VCC_net, \next_accum[16] , 
            \next_accum[17] , \next_accum[18] , \next_accum[19] , \next_accum[5] , 
            \next_accum[4] , rs2, rs1, rd, return_addr, \reg_access[4][3] , 
            \reg_access[3][2] , \instr[12] , n3645, \increment_result_3__N_1656[0] , 
            n25294, \increment_result_3__N_1642[1] , n25246, n22558, 
            n25218, n21812) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output n25273;
    input clk_c_enable_27;
    output \mie[0] ;
    input [3:0]n92;
    output instr_retired;
    output instr_complete_N_1378;
    input n25424;
    output cmp;
    input \imm[11] ;
    input instr_complete_N_1382;
    input \next_fsm_state_3__N_2230[3] ;
    output cy;
    output mstatus_mte;
    input clk_c_enable_111;
    output mstatus_mpie;
    input clk_c_enable_170;
    output \addr_out[11] ;
    output \addr_out[12] ;
    output \addr_out[13] ;
    output \addr_out[14] ;
    output \addr_out[15] ;
    input [4:2]counter_hi;
    output \addr_out[16] ;
    output \addr_out[17] ;
    output \addr_out[18] ;
    output \addr_out[19] ;
    output n25372;
    output n25365;
    output \addr_out[20] ;
    output \addr_out[21] ;
    output \addr_out[22] ;
    input \imm[6] ;
    output \addr_out[23] ;
    input \alu_op[1] ;
    input debug_instr_valid;
    input is_system;
    input \alu_op[0] ;
    output n25310;
    input n5;
    output clk_c_enable_205;
    output n25344;
    input \imm[1] ;
    output [6:0]cycle_count_wide;
    input \imm[0] ;
    input \next_pc_for_core[22] ;
    input \next_pc_for_core[18] ;
    output \mie[8] ;
    output [3:0]data_rs1;
    output n25179;
    output n25175;
    input n22208;
    output n25178;
    output n21248;
    input n22098;
    output n3615;
    input timer_interrupt;
    input n26608;
    input n22172;
    output n2037;
    input n22258;
    output n2835;
    input n22867;
    input n7955;
    input n24916;
    output n22272;
    input n22152;
    output n21113;
    input \alu_op_in[2] ;
    input n25430;
    input n22254;
    input n26;
    output n24486;
    input n22184;
    output n21260;
    input n22244;
    output n21230;
    input n22138;
    output n21121;
    input n22004;
    output n25182;
    output n25177;
    output n22008;
    input n22324;
    output n21303;
    input n22298;
    output n21297;
    input n22120;
    output n2236;
    input n22220;
    output n21242;
    input n25216;
    input n21910;
    output n21916;
    input n22933;
    output n22852;
    input n22086;
    input n25191;
    output n22092;
    input n22276;
    input n12;
    output n22282;
    input n21898;
    output n21212;
    input n22232;
    output n21236;
    input n23322;
    output \cycle[0] ;
    output \addr_out[3] ;
    input n11558;
    input \ui_in_sync[1] ;
    output n1092;
    input n25343;
    input n26610;
    input any_additional_mem_ops;
    output clk_c_enable_206;
    input n25349;
    input interrupt_core;
    output clk_c_enable_209;
    input is_load;
    output n54;
    input n20739;
    output clk_c_enable_393;
    output n21402;
    input [1:0]n4455;
    input [1:0]n1768;
    output [1:0]pc_2__N_663;
    output load_done;
    input n6638;
    input n1767;
    output \instr_write_offset_3__N_665[0] ;
    input n1766;
    output \instr_write_offset_3__N_665[1] ;
    output n25181;
    input [2:0]mem_op;
    input n5031;
    output \addr_out[6] ;
    output [3:0]debug_rd;
    input debug_rd_3__N_1306;
    output \addr_out[7] ;
    input n25369;
    input \imm[2] ;
    output n25410;
    output [15:0]accum;
    output [19:0]d_3__N_1599;
    input \imm[7] ;
    input \imm[8] ;
    input \imm[10] ;
    input \imm[9] ;
    input n24938;
    input \debug_branch_N_181[0] ;
    output \addr_out[4] ;
    input \mul_out[1] ;
    output n25421;
    output [3:0]data_rs2;
    input \debug_rd_3__N_136[28] ;
    output [3:0]alu_b_in;
    output n25316;
    output \addr_out[8] ;
    input \mul_out[3] ;
    output \mcause[2] ;
    output \alu_b_in[1] ;
    output \alu_a_in[1] ;
    output [3:0]n5047;
    output \alu_a_in[0] ;
    output n6657;
    input was_early_branch;
    output instr_fetch_restart_N_678;
    output data_out_3__N_1116;
    output \data_out_slice[1] ;
    output n22354;
    output mstatus_mie;
    output n21750;
    input n22028;
    output n22030;
    output n25180;
    input rst_reg_n;
    output n14111;
    output n20807;
    input \next_pc_offset[3] ;
    output n21864;
    input n25422;
    output n5_adj_1;
    output clk_c_enable_54;
    output \addr_out[10] ;
    input \debug_branch_N_173[28] ;
    input n22941;
    output \addr_out[0] ;
    input n25411;
    output n25333;
    output n25359;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[11] ;
    output load_top_bit;
    input \debug_branch_N_181[3] ;
    output n25352;
    output cy_adj_2;
    input data_ready_sync;
    input n25197;
    output data_ready_core;
    input n24186;
    output cy_adj_3;
    output \addr_out[5] ;
    output \instrret_count[0] ;
    output n23011;
    output n25408;
    input \debug_branch_N_173[30] ;
    output n25402;
    input n25350;
    output clk_c_enable_336;
    output n18;
    output clk_c_enable_197;
    output n23898;
    output n23897;
    output n23896;
    output n23895;
    output n23894;
    input \imm[4] ;
    output \addr_out[26] ;
    output n25307;
    output \addr_out[25] ;
    output \addr_out[24] ;
    input \alu_op[3] ;
    input is_alu_imm;
    input is_alu_reg;
    input is_auipc;
    input \debug_branch_N_173[29] ;
    input is_jal;
    input n25426;
    input \debug_rd_3__N_136[29] ;
    output n4996;
    input n24264;
    input is_jalr;
    output n25412;
    output n23395;
    input is_lui;
    input is_store;
    output \data_out_slice[0] ;
    input \debug_branch_N_571[29] ;
    input \timer_data[1] ;
    input is_timer_addr;
    input \imm[5] ;
    input \imm[3] ;
    input is_branch;
    output n25277;
    output \data_rs1[3] ;
    input n23111;
    input n25375;
    input n22798;
    input n25387;
    input \debug_rd_3__N_136[31] ;
    input \tmp_data_in_3__N_1245[3] ;
    input n25319;
    input \debug_rd_3__N_136[30] ;
    output \addr_out[9] ;
    input \debug_branch_N_173[31] ;
    input n25301;
    input \debug_rd_3__N_1298[0] ;
    output n25293;
    input n25282;
    input \mtimecmp[7] ;
    output mtimecmp_3__N_1666;
    output \data_out_slice[2] ;
    input n24932;
    input \debug_branch_N_181[2] ;
    input no_write_in_progress;
    input n25348;
    input n25326;
    input n23069;
    output \addr_out[1] ;
    input n22944;
    input \debug_branch_N_571[31] ;
    input n23073;
    input \debug_branch_N_177[31] ;
    input \mul_out[2] ;
    input n23067;
    input \debug_branch_N_177[29] ;
    input \next_pc_for_core[14] ;
    input \next_pc_for_core[10] ;
    input n66;
    output n12257;
    input \addr_offset[2] ;
    output n701;
    input n23070;
    input \debug_branch_N_177[30] ;
    input n25341;
    input n25271;
    input n22939;
    input n23012;
    output n25475;
    input \csr_read_3__N_1170[3] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input GND_net;
    input VCC_net;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[5] ;
    input \next_accum[4] ;
    input [3:0]rs2;
    input [3:0]rs1;
    input [3:0]rd;
    output [23:1]return_addr;
    output \reg_access[4][3] ;
    output \reg_access[3][2] ;
    input \instr[12] ;
    output n3645;
    input \increment_result_3__N_1656[0] ;
    input n25294;
    input \increment_result_3__N_1642[1] ;
    output n25246;
    input n22558;
    input n25218;
    input n21812;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [16:0]mie;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(323[16:19])
    
    wire clk_c_enable_190, n793, n20023;
    wire [17:16]mip_reg;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(321[17:24])
    wire [1:0]n979;
    
    wire n795;
    wire [31:0]tmp_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(88[16:24])
    
    wire clk_c_enable_255, n9319;
    wire [3:0]tmp_data_in_3__N_1245;
    wire [5:0]shift_amt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[16:25])
    
    wire clk_c_enable_161, n13946;
    wire [2:0]time_hi;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(292[15:22])
    wire [2:0]n1;
    wire [1:0]cycle;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(58[15:20])
    
    wire clk_c_enable_94, n19489, cmp_out;
    wire [23:0]mepc;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(68[16:20])
    
    wire clk_c_enable_396, n20586, n21576, n46, instr_complete_N_1383, 
        debug_rd_3__N_1132, instr_complete_N_1381;
    wire [5:0]mcause;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(325[15:21])
    
    wire clk_c_enable_279;
    wire [5:0]n611;
    wire [1:0]last_interrupt_req;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(417[15:33])
    
    wire clk_c_enable_280, cy_out, mstatus_mte_N_1434, n24884, n24882, 
        debug_rd_3__N_1131, debug_reg_wen;
    wire [4:0]shift_amt_adj_2358;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(124[15:24])
    
    wire clk_c_enable_158, clk_c_enable_162, n5400;
    wire [2:0]n498;
    
    wire n25390, n20692, n24865, n24863, n25366, n24866;
    wire [3:0]csr_read_3__N_1190;
    
    wire n22604;
    wire [3:0]csr_read_3__N_1186;
    
    wire n24577, n24576, n4404;
    wire [3:0]csr_read_3__N_1178;
    
    wire n25389;
    wire [3:0]n5013;
    
    wire n25460, n25459, n3, n25351, is_double_fault_r, n5287, n25474, 
        n25473, n23010, n25652, clk_c_enable_176, n20019, clk_c_enable_180, 
        n925, n926, n20033, n928, clk_c_enable_184, n892, n893, 
        n20031, n895, n25655;
    wire [3:0]debug_rd_3__N_1127;
    wire [3:0]debug_rd_3__N_1123;
    
    wire n652;
    wire [3:0]n653;
    
    wire n19, n24219, clk_c_enable_189, n859, n860, n20029, n862, 
        n20021, n24218;
    wire [3:0]data_rs1_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(83[16:24])
    
    wire n24266;
    wire [3:0]n234;
    
    wire n25849;
    wire [3:0]n191;
    
    wire n24268, n15, n25847, n25846;
    wire [1:0]n948;
    
    wire n25461;
    wire [1:0]n822;
    
    wire n25435, n21786, n25436, n25292, n25327, n25378, n24220, 
        n21036, n5094, n23334, n25296, n24221, n25388, n14329, 
        n22674, n17061, n20855, n24222;
    wire [3:0]time_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(299[16:26])
    
    wire n23368;
    wire [3:0]n5041;
    
    wire n23001, n9321;
    wire [3:0]n658;
    
    wire n8461, n22770;
    wire [3:0]debug_rd_3__N_1298;
    
    wire n24280, n24281;
    wire [3:0]n5003;
    
    wire n20677;
    wire [3:0]n5035;
    
    wire n20561, n25404;
    wire [3:0]n196;
    wire [3:0]alu_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(110[16:23])
    
    wire n25405, n18_c, n21, n16, n22698, n23306;
    wire [3:0]debug_rd_3__N_1302;
    
    wire n24694, n24693, n24695;
    wire [3:0]tmp_data_in_3__N_1313;
    wire [3:0]tmp_data_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(242[15:26])
    
    wire alu_b_in_3__N_1235, n25323;
    wire [3:0]alu_b_in_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[16:24])
    wire [3:0]alu_a_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[16:24])
    wire [3:0]n4411;
    
    wire n24569, n24571;
    wire [3:0]debug_rd_3__N_1290;
    
    wire n21695, instr_complete_N_1387, instr_complete_N_1385, n23081, 
        n5040, n20584, n8500, interrupt_pending_N_1402;
    wire [6:0]cycle_count_wide_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(279[16:32])
    
    wire n23078, n25428;
    wire [3:0]shift_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(132[16:25])
    
    wire n23385, n23094, n21778, clk_c_enable_320, mstatus_mie_N_1438, 
        n24265, clk_c_enable_359, n14438, n25318, n25308;
    wire [3:0]instrret_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(301[16:30])
    wire [4:0]increment_result_3__N_1642;
    
    wire n24258, n25298, n24257, n8_adj_2353, n24259, n25376, n82, 
        n5_adj_2354, n21446, n25425, n40, n22590;
    wire [3:0]csr_read_3__N_1182;
    wire [3:0]debug_rd_3__N_1294;
    
    wire instr_complete_N_1379, n13853, n8720;
    wire [3:0]n4994;
    
    wire n6452, n13929, n25254, n25250, n25251, n25367, n25274, 
        n25357, n25358, n23325, n25413, n24279, n22937, n14477, 
        n25309, n25270, n22602, n24278, n12484, n8_adj_2356, instr_complete_N_1380, 
        n25295, n39, n20, n22935, n33, n8448;
    wire [3:0]csr_read_3__N_1174;
    
    wire load_top_bit_next_N_1462, n25315, n25306;
    wire [2:0]n4495;
    
    wire n22450, n20_adj_2357, n23077, n25653, n24883;
    wire [65:0]dr_3__N_1595;
    
    wire n24864, n22927, n25850, n25848;
    wire [3:0]mul_out_3__N_1241;
    
    wire n23080, n22782, n22776, n23076, n23079, n25654;
    
    FD1P3IX mie__i2 (.D(n793), .SP(clk_c_enable_190), .CD(n25273), .CK(clk_c), 
            .Q(mie[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i2.GSR = "DISABLED";
    FD1P3IX mie__i1 (.D(n20023), .SP(clk_c_enable_190), .CD(n25273), .CK(clk_c), 
            .Q(mie[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i1.GSR = "DISABLED";
    FD1P3IX mip_reg__i17 (.D(n979[1]), .SP(clk_c_enable_27), .CD(n25273), 
            .CK(clk_c), .Q(mip_reg[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mip_reg__i17.GSR = "DISABLED";
    FD1P3IX mip_reg__i16 (.D(n979[0]), .SP(clk_c_enable_27), .CD(n25273), 
            .CK(clk_c), .Q(mip_reg[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mip_reg__i16.GSR = "DISABLED";
    FD1P3IX mie__i0 (.D(n795), .SP(clk_c_enable_190), .CD(n25273), .CK(clk_c), 
            .Q(\mie[0] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i0.GSR = "DISABLED";
    FD1P3IX tmp_data_i0_i29 (.D(tmp_data_in_3__N_1245[1]), .SP(clk_c_enable_255), 
            .CD(n9319), .CK(clk_c), .Q(tmp_data[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i29.GSR = "DISABLED";
    FD1P3AX shift_amt__i1 (.D(n92[0]), .SP(clk_c_enable_161), .CK(clk_c), 
            .Q(shift_amt[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i1.GSR = "DISABLED";
    FD1P3IX tmp_data_i0_i28 (.D(tmp_data_in_3__N_1245[0]), .SP(clk_c_enable_255), 
            .CD(n9319), .CK(clk_c), .Q(tmp_data[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i28.GSR = "DISABLED";
    FD1S3IX instr_retired_518 (.D(instr_complete_N_1378), .CK(clk_c), .CD(n13946), 
            .Q(instr_retired)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(303[12] 305[8])
    defparam instr_retired_518.GSR = "DISABLED";
    FD1S3IX time_hi__i0 (.D(n1[0]), .CK(clk_c), .CD(n25424), .Q(time_hi[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i0.GSR = "DISABLED";
    FD1P3IX cycle__i1 (.D(n19489), .SP(clk_c_enable_94), .CD(n25424), 
            .CK(clk_c), .Q(cycle[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam cycle__i1.GSR = "DISABLED";
    FD1S3AX cmp_511 (.D(cmp_out), .CK(clk_c), .Q(cmp)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(117[12] 120[8])
    defparam cmp_511.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i0 (.D(tmp_data[4]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i0.GSR = "DISABLED";
    FD1P3AX mepc_i0_i0 (.D(mepc[4]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i0.GSR = "DISABLED";
    PFUMX i66 (.BLUT(n20586), .ALUT(n21576), .C0(\imm[11] ), .Z(n46));
    PFUMX instr_complete_I_108 (.BLUT(instr_complete_N_1382), .ALUT(instr_complete_N_1383), 
          .C0(debug_rd_3__N_1132), .Z(instr_complete_N_1381)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    FD1P3IX mcause__i0 (.D(n611[0]), .SP(clk_c_enable_279), .CD(n25424), 
            .CK(clk_c), .Q(mcause[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i0.GSR = "DISABLED";
    FD1P3AX last_interrupt_req_i0_i0 (.D(\next_fsm_state_3__N_2230[3] ), .SP(clk_c_enable_280), 
            .CK(clk_c), .Q(last_interrupt_req[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam last_interrupt_req_i0_i0.GSR = "DISABLED";
    FD1S3AX cy_510 (.D(cy_out), .CK(clk_c), .Q(cy)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(117[12] 120[8])
    defparam cy_510.GSR = "DISABLED";
    FD1P3BX mstatus_mte_523 (.D(mstatus_mte_N_1434), .SP(clk_c_enable_111), 
            .CK(clk_c), .PD(n25424), .Q(mstatus_mte)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(384[18] 390[12])
    defparam mstatus_mte_523.GSR = "DISABLED";
    PFUMX i22364 (.BLUT(n24884), .ALUT(n24882), .C0(debug_rd_3__N_1131), 
          .Z(debug_reg_wen));
    FD1P3AX shift_amt__i5 (.D(n92[0]), .SP(clk_c_enable_158), .CK(clk_c), 
            .Q(shift_amt_adj_2358[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i5.GSR = "DISABLED";
    FD1P3AX shift_amt__i4 (.D(n92[3]), .SP(clk_c_enable_161), .CK(clk_c), 
            .Q(shift_amt_adj_2358[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i4.GSR = "DISABLED";
    FD1P3AX shift_amt__i3 (.D(n92[2]), .SP(clk_c_enable_161), .CK(clk_c), 
            .Q(shift_amt_adj_2358[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i3.GSR = "DISABLED";
    FD1P3AX shift_amt__i2 (.D(n92[1]), .SP(clk_c_enable_161), .CK(clk_c), 
            .Q(shift_amt[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i2.GSR = "DISABLED";
    FD1P3AX mstatus_mpie_525 (.D(n5400), .SP(clk_c_enable_162), .CK(clk_c), 
            .Q(mstatus_mpie)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam mstatus_mpie_525.GSR = "DISABLED";
    FD1P3IX time_hi__i2 (.D(n498[2]), .SP(clk_c_enable_170), .CD(n25424), 
            .CK(clk_c), .Q(time_hi[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i2.GSR = "DISABLED";
    LUT4 tmp_data_31__I_0_542_i12_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[11]), 
         .D(tmp_data[15]), .Z(\addr_out[11] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i13_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[12]), 
         .D(tmp_data[16]), .Z(\addr_out[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i14_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[13]), 
         .D(tmp_data[17]), .Z(\addr_out[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX i22352 (.BLUT(n24865), .ALUT(n24863), .C0(n25366), .Z(n24866));
    LUT4 tmp_data_31__I_0_542_i15_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[14]), 
         .D(tmp_data[18]), .Z(\addr_out[14] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i16_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[15]), 
         .D(tmp_data[19]), .Z(\addr_out[15] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .D(mip_reg[16]), .Z(csr_read_3__N_1190[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_4_lut_adj_206 (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .D(mip_reg[17]), .Z(csr_read_3__N_1190[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut_4_lut_adj_206.init = 16'h0400;
    LUT4 tmp_data_31__I_0_542_i17_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[16]), 
         .D(tmp_data[20]), .Z(\addr_out[16] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i18_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[17]), 
         .D(tmp_data[21]), .Z(\addr_out[17] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i19_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[18]), 
         .D(tmp_data[22]), .Z(\addr_out[18] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i20_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[19]), 
         .D(tmp_data[23]), .Z(\addr_out[19] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 csr_read_3__I_103_i4_4_lut (.A(mcause[3]), .B(n22604), .C(n25372), 
         .D(n25365), .Z(csr_read_3__N_1186[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(490[33] 493[57])
    defparam csr_read_3__I_103_i4_4_lut.init = 16'hca0a;
    LUT4 tmp_data_31__I_0_542_i21_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[20]), 
         .D(tmp_data[24]), .Z(\addr_out[20] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i22_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[21]), 
         .D(tmp_data[25]), .Z(\addr_out[21] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i23_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[22]), 
         .D(tmp_data[26]), .Z(\addr_out[22] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i23_3_lut_4_lut.init = 16'hf780;
    FD1P3IX time_hi__i1 (.D(n498[1]), .SP(clk_c_enable_170), .CD(n25424), 
            .CK(clk_c), .Q(time_hi[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i1.GSR = "DISABLED";
    LUT4 n24577_bdd_4_lut (.A(n24577), .B(n24576), .C(counter_hi[2]), 
         .D(n4404), .Z(csr_read_3__N_1178[1])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n24577_bdd_4_lut.init = 16'hca00;
    LUT4 mux_3095_i3_4_lut (.A(n25389), .B(mepc[2]), .C(\imm[6] ), .D(clk_c_enable_396), 
         .Z(n5013[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3095_i3_4_lut.init = 16'hca0a;
    LUT4 tmp_data_31__I_0_542_i24_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[23]), 
         .D(tmp_data[27]), .Z(\addr_out[23] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 i10270_4_lut_then_4_lut (.A(\alu_op[1] ), .B(debug_instr_valid), 
         .C(is_system), .D(\alu_op[0] ), .Z(n25460)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(78[10:20])
    defparam i10270_4_lut_then_4_lut.init = 16'h0080;
    LUT4 i10270_4_lut_else_4_lut (.A(\alu_op[1] ), .B(debug_instr_valid), 
         .C(is_system), .D(mip_reg[17]), .Z(n25459)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(78[10:20])
    defparam i10270_4_lut_else_4_lut.init = 16'h8000;
    LUT4 tmp_data_31__I_0_542_i3_3_lut_rep_574_4_lut (.A(n25390), .B(n20692), 
         .C(mepc[2]), .D(tmp_data[6]), .Z(n25310)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i3_3_lut_rep_574_4_lut.init = 16'hf780;
    LUT4 i11568_2_lut_4_lut (.A(n3), .B(n5), .C(n25351), .D(n4404), 
         .Z(csr_read_3__N_1178[0])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i11568_2_lut_4_lut.init = 16'hca00;
    FD1P3IX is_double_fault_r_520 (.D(n25344), .SP(clk_c_enable_205), .CD(n5287), 
            .CK(clk_c), .Q(is_double_fault_r)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(361[12] 364[8])
    defparam is_double_fault_r_520.GSR = "DISABLED";
    LUT4 i11744_4_lut_then_4_lut (.A(\imm[1] ), .B(mcause[4]), .C(counter_hi[4]), 
         .D(counter_hi[3]), .Z(n25474)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i11744_4_lut_then_4_lut.init = 16'h0008;
    LUT4 i11744_4_lut_else_4_lut (.A(mcause[0]), .B(\imm[1] ), .C(counter_hi[4]), 
         .D(counter_hi[3]), .Z(n25473)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i11744_4_lut_else_4_lut.init = 16'h0008;
    LUT4 i20735_3_lut (.A(cycle_count_wide[0]), .B(cycle_count_wide[3]), 
         .C(\imm[0] ), .Z(n23010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20735_3_lut.init = 16'hcaca;
    LUT4 next_pc_for_core_22__bdd_4_lut_23106 (.A(\next_pc_for_core[22] ), 
         .B(\next_pc_for_core[18] ), .C(counter_hi[3]), .D(counter_hi[2]), 
         .Z(n25652)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam next_pc_for_core_22__bdd_4_lut_23106.init = 16'h0a0c;
    FD1P3IX mie__i16 (.D(n20019), .SP(clk_c_enable_176), .CD(n25273), 
            .CK(clk_c), .Q(mie[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i16.GSR = "DISABLED";
    FD1P3IX mie__i15 (.D(n925), .SP(clk_c_enable_180), .CD(n25273), .CK(clk_c), 
            .Q(mie[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i15.GSR = "DISABLED";
    FD1P3IX mie__i14 (.D(n926), .SP(clk_c_enable_180), .CD(n25273), .CK(clk_c), 
            .Q(mie[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i14.GSR = "DISABLED";
    FD1P3IX mie__i13 (.D(n20033), .SP(clk_c_enable_180), .CD(n25273), 
            .CK(clk_c), .Q(mie[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i13.GSR = "DISABLED";
    FD1P3IX mie__i12 (.D(n928), .SP(clk_c_enable_180), .CD(n25273), .CK(clk_c), 
            .Q(mie[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i12.GSR = "DISABLED";
    FD1P3IX mie__i11 (.D(n892), .SP(clk_c_enable_184), .CD(n25273), .CK(clk_c), 
            .Q(mie[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i11.GSR = "DISABLED";
    FD1P3IX mie__i10 (.D(n893), .SP(clk_c_enable_184), .CD(n25273), .CK(clk_c), 
            .Q(mie[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i10.GSR = "DISABLED";
    FD1P3IX mie__i9 (.D(n20031), .SP(clk_c_enable_184), .CD(n25273), .CK(clk_c), 
            .Q(mie[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i9.GSR = "DISABLED";
    FD1P3IX mie__i8 (.D(n895), .SP(clk_c_enable_184), .CD(n25273), .CK(clk_c), 
            .Q(\mie[8] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i8.GSR = "DISABLED";
    LUT4 n25655_bdd_3_lut_22638 (.A(n25655), .B(debug_rd_3__N_1127[2]), 
         .C(debug_rd_3__N_1131), .Z(debug_rd_3__N_1123[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25655_bdd_3_lut_22638.init = 16'hcaca;
    LUT4 mux_251_i1_3_lut (.A(mepc[0]), .B(data_rs1[0]), .C(n652), .Z(n653[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i1_3_lut.init = 16'hcaca;
    LUT4 n19_bdd_4_lut_21980 (.A(n19), .B(mie[16]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n24219)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A !((C+(D))+!B)) */ ;
    defparam n19_bdd_4_lut_21980.init = 16'haa0c;
    FD1P3IX mie__i7 (.D(n859), .SP(clk_c_enable_189), .CD(n25273), .CK(clk_c), 
            .Q(mie[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i7.GSR = "DISABLED";
    FD1P3IX mie__i6 (.D(n860), .SP(clk_c_enable_189), .CD(n25273), .CK(clk_c), 
            .Q(mie[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i6.GSR = "DISABLED";
    FD1P3IX mie__i5 (.D(n20029), .SP(clk_c_enable_189), .CD(n25273), .CK(clk_c), 
            .Q(mie[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i5.GSR = "DISABLED";
    FD1P3IX mie__i4 (.D(n862), .SP(clk_c_enable_189), .CD(n25273), .CK(clk_c), 
            .Q(mie[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i4.GSR = "DISABLED";
    FD1P3IX mie__i3 (.D(n20021), .SP(clk_c_enable_190), .CD(n25273), .CK(clk_c), 
            .Q(mie[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i3.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_4_lut (.A(n25179), .B(n25175), .C(n22208), .D(n25178), 
         .Z(n21248)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_207 (.A(n25179), .B(n25175), .C(n22098), 
         .D(n25178), .Z(n3615)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_207.init = 16'h0040;
    LUT4 imm_6__bdd_4_lut_22422 (.A(counter_hi[2]), .B(timer_interrupt), 
         .C(counter_hi[3]), .D(n26608), .Z(n24218)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam imm_6__bdd_4_lut_22422.init = 16'h0008;
    LUT4 i2753_4_lut_4_lut_4_lut (.A(n25179), .B(n25175), .C(n22172), 
         .D(n25178), .Z(n2037)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i2753_4_lut_4_lut_4_lut.init = 16'hffbf;
    LUT4 i1_4_lut_4_lut_4_lut_adj_208 (.A(n25179), .B(n25175), .C(n22258), 
         .D(n25178), .Z(n2835)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_208.init = 16'h0040;
    LUT4 i1_4_lut_4_lut (.A(n25179), .B(n22867), .C(n7955), .D(n24916), 
         .Z(n22272)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_4_lut_4_lut_adj_209 (.A(n25179), .B(n25175), .C(n22152), 
         .D(n25178), .Z(n21113)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_209.init = 16'h0040;
    LUT4 i1_4_lut (.A(\alu_op_in[2] ), .B(n25430), .C(\alu_op[1] ), .D(\alu_op[0] ), 
         .Z(n20692)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut.init = 16'h0004;
    LUT4 n10_bdd_4_lut_4_lut (.A(n25179), .B(n22254), .C(n26), .D(n25175), 
         .Z(n24486)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam n10_bdd_4_lut_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_4_lut_4_lut_adj_210 (.A(n25179), .B(n25175), .C(n22184), 
         .D(n25178), .Z(n21260)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_210.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_211 (.A(n25179), .B(n25175), .C(n22244), 
         .D(n25178), .Z(n21230)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_211.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_212 (.A(n25179), .B(n25175), .C(n22138), 
         .D(n25178), .Z(n21121)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_212.init = 16'h0040;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n25179), .B(n22004), .C(n25182), .D(n25177), 
         .Z(n22008)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 i1_4_lut_4_lut_4_lut_adj_213 (.A(n25179), .B(n25175), .C(n22324), 
         .D(n25178), .Z(n21303)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_213.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_214 (.A(n25179), .B(n25175), .C(n22298), 
         .D(n25178), .Z(n21297)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_214.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_215 (.A(n25179), .B(n25175), .C(n22120), 
         .D(n25178), .Z(n2236)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_215.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_216 (.A(n25179), .B(n25175), .C(n22220), 
         .D(n25178), .Z(n21242)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_216.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_217 (.A(n25179), .B(n25216), .C(n21910), .D(n7955), 
         .Z(n21916)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_217.init = 16'h0010;
    LUT4 i20640_4_lut_4_lut_4_lut (.A(n25179), .B(n25175), .C(n22933), 
         .D(n25178), .Z(n22852)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i20640_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_218 (.A(n25179), .B(n22086), .C(n25191), .D(n7955), 
         .Z(n22092)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_218.init = 16'h0040;
    LUT4 mux_251_i3_3_lut (.A(mepc[2]), .B(data_rs1_c[2]), .C(n652), .Z(n653[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i3_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_219 (.A(n25179), .B(n22276), .C(n12), .D(n7955), 
         .Z(n22282)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_219.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_220 (.A(n25179), .B(n25175), .C(n21898), 
         .D(n25178), .Z(n21212)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_220.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_221 (.A(n25179), .B(n25175), .C(n22232), 
         .D(n25178), .Z(n21236)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_221.init = 16'h0040;
    LUT4 mux_251_i2_3_lut (.A(mepc[1]), .B(data_rs1_c[1]), .C(n652), .Z(n653[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i2_3_lut.init = 16'hcaca;
    LUT4 n24266_bdd_3_lut (.A(n24266), .B(n234[3]), .C(n23322), .Z(n25849)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n24266_bdd_3_lut.init = 16'hacac;
    LUT4 n192_bdd_4_lut (.A(n191[3]), .B(n24268), .C(n15), .D(n25366), 
         .Z(n25847)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(((D)+!C)+!B)) */ ;
    defparam n192_bdd_4_lut.init = 16'ha0c0;
    LUT4 n192_bdd_3_lut (.A(cycle[1]), .B(\cycle[0] ), .C(tmp_data[3]), 
         .Z(n25846)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam n192_bdd_3_lut.init = 16'h4040;
    LUT4 tmp_data_31__I_0_542_i4_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[3]), 
         .D(tmp_data[7]), .Z(\addr_out[3] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i11876_4_lut (.A(mip_reg[17]), .B(n11558), .C(\ui_in_sync[1] ), 
         .D(last_interrupt_req[1]), .Z(n948[1])) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(447[18] 459[12])
    defparam i11876_4_lut.init = 16'h88c8;
    LUT4 i11875_4_lut (.A(n25461), .B(n1092), .C(data_rs1_c[1]), .D(n25343), 
         .Z(n822[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(434[22] 438[16])
    defparam i11875_4_lut.init = 16'hc088;
    LUT4 i1_2_lut_rep_699 (.A(n26610), .B(n26608), .Z(n25435)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_699.init = 16'heeee;
    LUT4 i2_rep_443 (.A(any_additional_mem_ops), .B(clk_c_enable_206), .C(instr_complete_N_1378), 
         .D(n21786), .Z(n25179)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i2_rep_443.init = 16'h4000;
    LUT4 i1_2_lut_rep_442_4_lut (.A(n25349), .B(instr_complete_N_1378), 
         .C(clk_c_enable_206), .D(any_additional_mem_ops), .Z(n25178)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_rep_442_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_556_3_lut_3_lut_4_lut (.A(n25436), .B(n20692), .C(interrupt_core), 
         .D(n25349), .Z(n25292)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_556_3_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_1_lut_rep_437_2_lut_4_lut (.A(n25349), .B(instr_complete_N_1378), 
         .C(clk_c_enable_206), .D(any_additional_mem_ops), .Z(clk_c_enable_209)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_1_lut_rep_437_2_lut_4_lut.init = 16'hbfff;
    LUT4 i21880_2_lut_4_lut (.A(n25349), .B(instr_complete_N_1378), .C(n25327), 
         .D(is_load), .Z(n54)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i21880_2_lut_4_lut.init = 16'h40ff;
    LUT4 i1_2_lut_4_lut (.A(n25349), .B(instr_complete_N_1378), .C(n25327), 
         .D(n20739), .Z(clk_c_enable_393)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_4_lut.init = 16'hff40;
    LUT4 interrupt_core_I_7_2_lut_rep_441_4_lut (.A(n25349), .B(instr_complete_N_1378), 
         .C(n25327), .D(n21402), .Z(n25177)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam interrupt_core_I_7_2_lut_rep_441_4_lut.init = 16'h40ff;
    LUT4 mux_233_i2_3_lut_4_lut (.A(n25436), .B(n20692), .C(interrupt_core), 
         .D(n25378), .Z(n611[1])) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_233_i2_3_lut_4_lut.init = 16'hf404;
    LUT4 i1_3_lut_4_lut (.A(instr_complete_N_1378), .B(clk_c_enable_206), 
         .C(cycle[1]), .D(\cycle[0] ), .Z(n19489)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_4_lut.init = 16'h0770;
    LUT4 n19_bdd_4_lut_22814 (.A(mie[11]), .B(mie[3]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n24220)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !((C+!(D))+!B)) */ ;
    defparam n19_bdd_4_lut_22814.init = 16'hac00;
    LUT4 mux_352_i1_3_lut_4_lut (.A(clk_c_enable_206), .B(n21036), .C(n4455[0]), 
         .D(n1768[0]), .Z(pc_2__N_663[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_352_i1_3_lut_4_lut.init = 16'hf780;
    FD1P3AX load_done_515 (.D(n6638), .SP(clk_c_enable_205), .CK(clk_c), 
            .Q(load_done)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(232[12] 235[8])
    defparam load_done_515.GSR = "DISABLED";
    LUT4 mux_351_i1_3_lut_4_lut (.A(clk_c_enable_206), .B(n21036), .C(n4455[0]), 
         .D(n1767), .Z(\instr_write_offset_3__N_665[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_351_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i21916_2_lut_3_lut_4_lut (.A(n25436), .B(n20692), .C(n5094), 
         .D(interrupt_core), .Z(n23334)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i21916_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 i11878_2_lut_rep_560_3_lut_3_lut_4_lut (.A(n25436), .B(n20692), 
         .C(interrupt_core), .D(n25372), .Z(n25296)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam i11878_2_lut_rep_560_3_lut_3_lut_4_lut.init = 16'h00f4;
    LUT4 i7055_2_lut_3_lut_4_lut (.A(n25436), .B(n20692), .C(clk_c_enable_255), 
         .D(interrupt_core), .Z(n9319)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i7055_2_lut_3_lut_4_lut.init = 16'hf040;
    LUT4 mux_352_i2_3_lut_4_lut (.A(clk_c_enable_206), .B(n21036), .C(n4455[1]), 
         .D(n1768[1]), .Z(pc_2__N_663[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_352_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_351_i2_3_lut_4_lut (.A(clk_c_enable_206), .B(n21036), .C(n4455[1]), 
         .D(n1766), .Z(\instr_write_offset_3__N_665[1] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_351_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 interrupt_core_I_6_2_lut_rep_439_3_lut_4_lut (.A(clk_c_enable_206), 
         .B(n21036), .C(n25181), .D(n21402), .Z(n25175)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (C+!(D))) */ ;
    defparam interrupt_core_I_6_2_lut_rep_439_3_lut_4_lut.init = 16'hf8ff;
    PFUMX i21981 (.BLUT(n24220), .ALUT(n24219), .C0(counter_hi[2]), .Z(n24221));
    LUT4 i12249_3_lut_4_lut (.A(n26608), .B(n25388), .C(mem_op[0]), .D(n25365), 
         .Z(n14329)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(149[15:31])
    defparam i12249_3_lut_4_lut.init = 16'hbfb0;
    LUT4 i11582_4_lut (.A(mip_reg[16]), .B(n11558), .C(\next_fsm_state_3__N_2230[3] ), 
         .D(last_interrupt_req[0]), .Z(n948[0])) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(447[18] 459[12])
    defparam i11582_4_lut.init = 16'h88c8;
    LUT4 i11577_4_lut (.A(n22674), .B(n1092), .C(n17061), .D(n20855), 
         .Z(n822[0])) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(434[22] 438[16])
    defparam i11577_4_lut.init = 16'hc8c0;
    LUT4 n24221_bdd_3_lut_22821 (.A(n24221), .B(n24218), .C(\imm[6] ), 
         .Z(n24222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24221_bdd_3_lut_22821.init = 16'hcaca;
    PFUMX mux_3107_i3 (.BLUT(time_count[2]), .ALUT(n5031), .C0(n23368), 
          .Z(n5041[2]));
    LUT4 i20726_3_lut (.A(cycle_count_wide[1]), .B(time_count[1]), .C(\imm[0] ), 
         .Z(n23001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20726_3_lut.init = 16'hcaca;
    LUT4 tmp_data_31__I_0_542_i7_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[6]), 
         .D(tmp_data[10]), .Z(\addr_out[6] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i7_3_lut_4_lut.init = 16'hf780;
    FD1P3AX tmp_data_i0_i1 (.D(tmp_data[5]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i1.GSR = "DISABLED";
    FD1P3IX mepc_i0_i23 (.D(n658[3]), .SP(clk_c_enable_396), .CD(n9321), 
            .CK(clk_c), .Q(mepc[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i23.GSR = "DISABLED";
    LUT4 i18_3_lut (.A(mie[7]), .B(mie[15]), .C(counter_hi[3]), .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(139[15:25])
    defparam i18_3_lut.init = 16'hcaca;
    L6MUX21 debug_rd_3__I_0_i1 (.D0(debug_rd_3__N_1123[0]), .D1(debug_rd_3__N_1127[0]), 
            .SD(debug_rd_3__N_1131), .Z(debug_rd[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_4_lut_adj_222 (.A(\cycle[0] ), .B(n8461), .C(n25435), .D(n22770), 
         .Z(n15)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_4_lut_adj_222.init = 16'hfffd;
    LUT4 i1_2_lut (.A(counter_hi[2]), .B(cycle[1]), .Z(n22770)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(96[19:40])
    defparam i1_2_lut.init = 16'heeee;
    PFUMX i22016 (.BLUT(debug_rd_3__N_1298[1]), .ALUT(n24280), .C0(debug_rd_3__N_1306), 
          .Z(n24281));
    LUT4 mux_3105_i2_4_lut (.A(n5003[1]), .B(mepc[1]), .C(\imm[0] ), .D(n20677), 
         .Z(n5035[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3105_i2_4_lut.init = 16'hca0a;
    LUT4 tmp_data_31__I_0_542_i8_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[7]), 
         .D(tmp_data[11]), .Z(\addr_out[7] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 i21744_4_lut (.A(\imm[6] ), .B(n25369), .C(\imm[2] ), .D(n20561), 
         .Z(n1092)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i21744_4_lut.init = 16'h0080;
    LUT4 mux_73_i1_4_lut (.A(cmp), .B(tmp_data[0]), .C(n25410), .D(n25404), 
         .Z(n196[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(170[18] 174[35])
    defparam mux_73_i1_4_lut.init = 16'hca0a;
    LUT4 mux_72_i1_4_lut (.A(accum[0]), .B(alu_out[0]), .C(n25405), .D(d_3__N_1599[0]), 
         .Z(n191[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(174[17:35])
    defparam mux_72_i1_4_lut.init = 16'hc5ca;
    LUT4 i1_4_lut_adj_223 (.A(n18_c), .B(n21), .C(n16), .D(n22698), 
         .Z(n20561)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam i1_4_lut_adj_223.init = 16'hfffe;
    LUT4 i1_2_lut_adj_224 (.A(\imm[0] ), .B(\imm[1] ), .Z(n22698)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam i1_2_lut_adj_224.init = 16'heeee;
    LUT4 imm_lo_11__I_0_536_i18_2_lut (.A(\imm[7] ), .B(\imm[8] ), .Z(n18_c)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam imm_lo_11__I_0_536_i18_2_lut.init = 16'hbbbb;
    LUT4 i1_3_lut (.A(\imm[10] ), .B(\imm[9] ), .C(\imm[11] ), .Z(n21)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_3_lut.init = 16'hfbfb;
    LUT4 mux_87_i1_3_lut (.A(n24938), .B(\debug_branch_N_181[0] ), .C(n23306), 
         .Z(debug_rd_3__N_1302[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam mux_87_i1_3_lut.init = 16'hcaca;
    LUT4 tmp_data_31__I_0_542_i5_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[4]), 
         .D(tmp_data[8]), .Z(\addr_out[4] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_72_i2_3_lut (.A(\mul_out[1] ), .B(alu_out[1]), .C(n25405), 
         .Z(n191[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(174[17:35])
    defparam mux_72_i2_3_lut.init = 16'hcaca;
    PFUMX i22246 (.BLUT(n24694), .ALUT(n24693), .C0(\imm[10] ), .Z(n24695));
    LUT4 mux_149_i1_3_lut_4_lut (.A(n25421), .B(n25405), .C(alu_out[0]), 
         .D(data_rs2[0]), .Z(tmp_data_in_3__N_1313[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i1_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX tmp_data_i0_i2 (.D(tmp_data[6]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i2.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i3 (.D(tmp_data[7]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i3.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i4 (.D(tmp_data[8]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i4.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i5 (.D(tmp_data[9]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i5.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i6 (.D(tmp_data[10]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i6.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i7 (.D(tmp_data[11]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i7.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i8 (.D(tmp_data[12]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i8.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i9 (.D(tmp_data[13]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i9.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i10 (.D(tmp_data[14]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i10.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i11 (.D(tmp_data[15]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i11.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i12 (.D(tmp_data[16]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i12.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i13 (.D(tmp_data[17]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i13.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i14 (.D(tmp_data[18]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i14.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i15 (.D(tmp_data[19]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i15.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i16 (.D(tmp_data[20]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i16.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i17 (.D(tmp_data[21]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i17.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i18 (.D(tmp_data[22]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i18.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i19 (.D(tmp_data[23]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i19.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i20 (.D(tmp_data[24]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i20.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i21 (.D(tmp_data[25]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i21.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i22 (.D(tmp_data[26]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i22.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i23 (.D(tmp_data[27]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i23.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i24 (.D(tmp_data[28]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i24.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i25 (.D(tmp_data[29]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i25.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i26 (.D(tmp_data[30]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i26.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i27 (.D(tmp_data[31]), .SP(clk_c_enable_255), .CK(clk_c), 
            .Q(tmp_data[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i27.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i30 (.D(tmp_data_in[2]), .SP(clk_c_enable_255), 
            .CK(clk_c), .Q(tmp_data[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i30.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i31 (.D(tmp_data_in[3]), .SP(clk_c_enable_255), 
            .CK(clk_c), .Q(tmp_data[31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i31.GSR = "DISABLED";
    FD1P3AX mepc_i0_i1 (.D(mepc[5]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i1.GSR = "DISABLED";
    LUT4 imm_3__I_0_i1_3_lut (.A(\debug_rd_3__N_136[28] ), .B(data_rs2[0]), 
         .C(alu_b_in_3__N_1235), .Z(alu_b_in[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 mux_149_i2_3_lut_4_lut (.A(n25421), .B(n25405), .C(alu_out[1]), 
         .D(data_rs2[1]), .Z(tmp_data_in_3__N_1313[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_149_i3_3_lut_4_lut (.A(n25421), .B(n25405), .C(alu_out[2]), 
         .D(data_rs2[2]), .Z(tmp_data_in_3__N_1313[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_149_i4_3_lut_4_lut (.A(n25421), .B(n25405), .C(alu_out[3]), 
         .D(data_rs2[3]), .Z(tmp_data_in_3__N_1313[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 tmp_data_in_3__I_99_i3_4_lut (.A(data_rs1_c[2]), .B(mstatus_mte), 
         .C(n25316), .D(n25323), .Z(tmp_data_in_3__N_1245[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_99_i3_4_lut.init = 16'hca0a;
    LUT4 mux_2671_i3_3_lut_4_lut (.A(\alu_op[0] ), .B(n25410), .C(alu_b_in_c[2]), 
         .D(alu_a_in[2]), .Z(n4411[2])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam mux_2671_i3_3_lut_4_lut.init = 16'hfdd0;
    FD1P3AX mepc_i0_i2 (.D(mepc[6]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i2.GSR = "DISABLED";
    FD1P3AX mepc_i0_i3 (.D(mepc[7]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i3.GSR = "DISABLED";
    FD1P3AX mepc_i0_i4 (.D(mepc[8]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i4.GSR = "DISABLED";
    FD1P3AX mepc_i0_i5 (.D(mepc[9]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i5.GSR = "DISABLED";
    FD1P3AX mepc_i0_i6 (.D(mepc[10]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i6.GSR = "DISABLED";
    FD1P3AX mepc_i0_i7 (.D(mepc[11]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i7.GSR = "DISABLED";
    FD1P3AX mepc_i0_i8 (.D(mepc[12]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i8.GSR = "DISABLED";
    FD1P3AX mepc_i0_i9 (.D(mepc[13]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i9.GSR = "DISABLED";
    FD1P3AX mepc_i0_i10 (.D(mepc[14]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i10.GSR = "DISABLED";
    FD1P3AX mepc_i0_i11 (.D(mepc[15]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i11.GSR = "DISABLED";
    FD1P3AX mepc_i0_i12 (.D(mepc[16]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i12.GSR = "DISABLED";
    FD1P3AX mepc_i0_i13 (.D(mepc[17]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i13.GSR = "DISABLED";
    FD1P3AX mepc_i0_i14 (.D(mepc[18]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i14.GSR = "DISABLED";
    FD1P3AX mepc_i0_i15 (.D(mepc[19]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i15.GSR = "DISABLED";
    FD1P3AX mepc_i0_i16 (.D(mepc[20]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i16.GSR = "DISABLED";
    FD1P3AX mepc_i0_i17 (.D(mepc[21]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i17.GSR = "DISABLED";
    FD1P3AX mepc_i0_i18 (.D(mepc[22]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i18.GSR = "DISABLED";
    FD1P3AX mepc_i0_i19 (.D(mepc[23]), .SP(clk_c_enable_396), .CK(clk_c), 
            .Q(mepc[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i19.GSR = "DISABLED";
    FD1P3IX mcause__i1 (.D(n611[1]), .SP(clk_c_enable_279), .CD(n25424), 
            .CK(clk_c), .Q(mcause[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i1.GSR = "DISABLED";
    LUT4 n24571_bdd_3_lut_4_lut (.A(\alu_op[0] ), .B(n25410), .C(n24569), 
         .D(n24571), .Z(cmp_out)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam n24571_bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 tmp_data_31__I_0_542_i9_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[8]), 
         .D(tmp_data[12]), .Z(\addr_out[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 i11856_2_lut (.A(n24866), .B(n15), .Z(debug_rd_3__N_1290[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[18] 174[35])
    defparam i11856_2_lut.init = 16'h8888;
    LUT4 mux_72_i4_3_lut (.A(\mul_out[3] ), .B(alu_out[3]), .C(n25405), 
         .Z(n191[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(174[17:35])
    defparam mux_72_i4_3_lut.init = 16'hcaca;
    FD1P3IX mcause__i2 (.D(n611[2]), .SP(clk_c_enable_279), .CD(n25424), 
            .CK(clk_c), .Q(\mcause[2] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i2.GSR = "DISABLED";
    FD1P3IX mcause__i3 (.D(n21695), .SP(clk_c_enable_279), .CD(n25424), 
            .CK(clk_c), .Q(mcause[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i3.GSR = "DISABLED";
    FD1P3IX mcause__i4 (.D(n611[4]), .SP(clk_c_enable_279), .CD(n25424), 
            .CK(clk_c), .Q(mcause[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i4.GSR = "DISABLED";
    FD1P3IX mcause__i5 (.D(interrupt_core), .SP(clk_c_enable_279), .CD(n25424), 
            .CK(clk_c), .Q(mcause[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i5.GSR = "DISABLED";
    FD1P3AX last_interrupt_req_i0_i1 (.D(\ui_in_sync[1] ), .SP(clk_c_enable_280), 
            .CK(clk_c), .Q(last_interrupt_req[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam last_interrupt_req_i0_i1.GSR = "DISABLED";
    LUT4 mux_2671_i2_3_lut_4_lut (.A(\alu_op[0] ), .B(n25410), .C(\alu_b_in[1] ), 
         .D(\alu_a_in[1] ), .Z(n4411[1])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam mux_2671_i2_3_lut_4_lut.init = 16'hfdd0;
    LUT4 mux_2671_i4_3_lut_4_lut (.A(\alu_op[0] ), .B(n25410), .C(alu_b_in_c[3]), 
         .D(alu_a_in[3]), .Z(n4411[3])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam mux_2671_i4_3_lut_4_lut.init = 16'hfdd0;
    LUT4 i1_3_lut_adj_225 (.A(tmp_data[30]), .B(tmp_data[31]), .C(\cycle[0] ), 
         .Z(instr_complete_N_1387)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_adj_225.init = 16'hf7f7;
    LUT4 cycle_0__I_0_548_3_lut (.A(\cycle[0] ), .B(cmp_out), .C(\alu_op[0] ), 
         .Z(instr_complete_N_1385)) /* synthesis lut_function=(A+!(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(224[34:67])
    defparam cycle_0__I_0_548_3_lut.init = 16'hbebe;
    LUT4 mux_3109_i1_3_lut (.A(n5041[0]), .B(n23081), .C(n5040), .Z(n5047[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3109_i1_3_lut.init = 16'hcaca;
    LUT4 mux_2671_i1_3_lut_4_lut (.A(\alu_op[0] ), .B(n25410), .C(alu_b_in[0]), 
         .D(\alu_a_in[0] ), .Z(n4411[0])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam mux_2671_i1_3_lut_4_lut.init = 16'hfdd0;
    LUT4 i1_3_lut_adj_226 (.A(n25369), .B(n46), .C(\imm[7] ), .Z(n6657)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(190[18] 194[12])
    defparam i1_3_lut_adj_226.init = 16'h0808;
    LUT4 i1_4_lut_adj_227 (.A(n20584), .B(n8500), .C(\imm[7] ), .D(\imm[11] ), 
         .Z(n5040)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_227.init = 16'h0008;
    LUT4 debug_branch_N_172_I_0_2_lut_3_lut_4_lut (.A(n26608), .B(n25388), 
         .C(was_early_branch), .D(n21036), .Z(instr_fetch_restart_N_678)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam debug_branch_N_172_I_0_2_lut_3_lut_4_lut.init = 16'hf7ff;
    LUT4 i11864_2_lut (.A(data_rs2[1]), .B(data_out_3__N_1116), .Z(\data_out_slice[1] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i11864_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut (.A(counter_hi[4]), .B(n25388), .C(n21402), 
         .D(n21036), .Z(n22354)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i1_3_lut_4_lut_adj_228 (.A(counter_hi[4]), .B(n25388), .C(mstatus_mie), 
         .D(interrupt_pending_N_1402), .Z(n21750)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_228.init = 16'h8000;
    LUT4 cycle_count_wide_6__I_0_3_lut_4_lut (.A(counter_hi[4]), .B(n25388), 
         .C(time_hi[2]), .D(cycle_count_wide_c[6]), .Z(time_count[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam cycle_count_wide_6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_229 (.A(counter_hi[4]), .B(n25388), .C(n22028), 
         .D(n21036), .Z(n22030)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_229.init = 16'h70f0;
    LUT4 i1_3_lut_rep_444_4_lut (.A(n26608), .B(n25388), .C(instr_complete_N_1378), 
         .D(n25349), .Z(n25180)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_rep_444_4_lut.init = 16'h0080;
    LUT4 cycle_count_wide_5__I_0_3_lut_4_lut (.A(counter_hi[4]), .B(n25388), 
         .C(time_hi[1]), .D(cycle_count_wide_c[5]), .Z(time_count[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam cycle_count_wide_5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i11727_2_lut_3_lut_4_lut (.A(counter_hi[4]), .B(n25388), .C(interrupt_core), 
         .D(n25349), .Z(n13946)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;
    defparam i11727_2_lut_3_lut_4_lut.init = 16'h7f77;
    LUT4 i21735_2_lut_3_lut_4_lut (.A(counter_hi[4]), .B(n25388), .C(rst_reg_n), 
         .D(n14111), .Z(clk_c_enable_94)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i21735_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i18656_2_lut_3_lut_4_lut (.A(counter_hi[4]), .B(n25388), .C(rst_reg_n), 
         .D(n21036), .Z(n20807)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i18656_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 cycle_count_wide_4__I_0_3_lut_4_lut (.A(counter_hi[4]), .B(n25388), 
         .C(time_hi[0]), .D(cycle_count_wide_c[4]), .Z(time_count[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam cycle_count_wide_4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_230 (.A(n26608), .B(n25388), .C(\next_pc_offset[3] ), 
         .D(any_additional_mem_ops), .Z(n21864)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_230.init = 16'h0080;
    LUT4 i1_3_lut_rep_603_4_lut (.A(n26608), .B(n25388), .C(n25422), .D(n5_adj_1), 
         .Z(clk_c_enable_54)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_rep_603_4_lut.init = 16'h8000;
    LUT4 tmp_data_31__I_0_542_i11_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[10]), 
         .D(tmp_data[14]), .Z(\addr_out[10] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 i6467_4_lut (.A(mem_op[1]), .B(mem_op[0]), .C(n26608), .D(counter_hi[3]), 
         .Z(data_out_3__N_1116)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[13] 272[50])
    defparam i6467_4_lut.init = 16'h5150;
    LUT4 mux_3109_i4_3_lut (.A(n23078), .B(n5035[3]), .C(n5040), .Z(n5047[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3109_i4_3_lut.init = 16'hcaca;
    LUT4 i21547_3_lut_4_lut (.A(n25404), .B(n25428), .C(n191[1]), .D(shift_out[1]), 
         .Z(n196[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i21547_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i21886_3_lut_4_lut (.A(n25404), .B(n25428), .C(n15), .D(n25410), 
         .Z(n23385)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i21886_3_lut_4_lut.init = 16'hffdf;
    LUT4 i21540_4_lut_4_lut (.A(n25410), .B(n15), .C(n196[0]), .D(n191[0]), 
         .Z(debug_rd_3__N_1290[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;
    defparam i21540_4_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_3105_i4_4_lut (.A(n24222), .B(mepc[3]), .C(\imm[0] ), .D(n20677), 
         .Z(n5035[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3105_i4_4_lut.init = 16'hca0a;
    LUT4 i11778_4_lut_4_lut (.A(n25410), .B(n23094), .C(\debug_branch_N_173[28] ), 
         .D(n22941), .Z(\alu_a_in[0] )) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;
    defparam i11778_4_lut_4_lut.init = 16'h5410;
    LUT4 tmp_data_31__I_0_542_i1_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[0]), 
         .D(tmp_data[4]), .Z(\addr_out[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i18702_3_lut_4_lut_3_lut_4_lut_4_lut (.A(n25430), .B(\alu_op[0] ), 
         .C(\alu_op[1] ), .D(data_rs1[0]), .Z(n20855)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(75[19:52])
    defparam i18702_3_lut_4_lut_3_lut_4_lut_4_lut.init = 16'h20a0;
    LUT4 i1_4_lut_adj_231 (.A(n21778), .B(cmp_out), .C(n25411), .D(mem_op[0]), 
         .Z(n21036)) /* synthesis lut_function=(A+!(B ((D)+!C)+!B !(C (D)))) */ ;
    defparam i1_4_lut_adj_231.init = 16'hbaea;
    FD1P3AX mstatus_mie_524 (.D(mstatus_mie_N_1438), .SP(clk_c_enable_320), 
            .CK(clk_c), .Q(mstatus_mie)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam mstatus_mie_524.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_232 (.A(n25344), .B(n25333), .C(n25359), .D(interrupt_core), 
         .Z(n21778)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_232.init = 16'hfffe;
    LUT4 next_pc_for_core_23__bdd_3_lut (.A(\next_pc_for_core[15] ), .B(\next_pc_for_core[11] ), 
         .C(counter_hi[2]), .Z(n24265)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam next_pc_for_core_23__bdd_3_lut.init = 16'hacac;
    FD1P3IX load_top_bit_513 (.D(\debug_branch_N_181[3] ), .SP(clk_c_enable_359), 
            .CD(n14438), .CK(clk_c), .Q(load_top_bit)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(156[12] 157[43])
    defparam load_top_bit_513.GSR = "DISABLED";
    LUT4 cy_I_0_3_lut_rep_582_3_lut_4_lut (.A(n25435), .B(counter_hi[2]), 
         .C(cy), .D(n25352), .Z(n25318)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam cy_I_0_3_lut_rep_582_3_lut_4_lut.init = 16'hf1e0;
    LUT4 cy_I_0_3_lut_rep_572_3_lut_4_lut (.A(n25435), .B(counter_hi[2]), 
         .C(cy_adj_2), .D(instr_retired), .Z(n25308)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam cy_I_0_3_lut_rep_572_3_lut_4_lut.init = 16'hf1e0;
    LUT4 imm_10__bdd_3_lut_22245_3_lut_4_lut (.A(n25435), .B(counter_hi[2]), 
         .C(instrret_count[1]), .D(\imm[0] ), .Z(n24693)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam imm_10__bdd_3_lut_22245_3_lut_4_lut.init = 16'h11f0;
    LUT4 imm_10__bdd_3_lut_3_lut_4_lut (.A(n25435), .B(counter_hi[2]), .C(\imm[1] ), 
         .D(mcause[1]), .Z(n24694)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam imm_10__bdd_3_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 data_ready_sync_I_0_3_lut_3_lut_4_lut (.A(n25435), .B(counter_hi[2]), 
         .C(data_ready_sync), .D(n25197), .Z(data_ready_core)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam data_ready_sync_I_0_3_lut_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX cycle__i0 (.D(n24186), .CK(clk_c), .Q(\cycle[0] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam cycle__i0.GSR = "DISABLED";
    LUT4 i3918_2_lut_3_lut_3_lut_4_lut (.A(n25435), .B(counter_hi[2]), .C(cy_adj_3), 
         .D(cycle_count_wide[0]), .Z(increment_result_3__N_1642[0])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam i3918_2_lut_3_lut_3_lut_4_lut.init = 16'h0ef1;
    LUT4 counter_hi_2__bdd_4_lut_22180 (.A(mie[10]), .B(mie[2]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n24258)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam counter_hi_2__bdd_4_lut_22180.init = 16'hacaa;
    LUT4 tmp_data_31__I_0_542_i6_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[5]), 
         .D(tmp_data[9]), .Z(\addr_out[5] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 i3920_2_lut_rep_562_3_lut_3_lut_4_lut (.A(n25435), .B(counter_hi[2]), 
         .C(cy_adj_3), .D(cycle_count_wide[0]), .Z(n25298)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (D))) */ ;
    defparam i3920_2_lut_rep_562_3_lut_3_lut_4_lut.init = 16'hf100;
    LUT4 i20736_3_lut_3_lut_4_lut (.A(n25435), .B(counter_hi[2]), .C(\instrret_count[0] ), 
         .D(\imm[0] ), .Z(n23011)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam i20736_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i1_2_lut_rep_587_3_lut_4_lut (.A(n25435), .B(counter_hi[2]), .C(n20692), 
         .D(n25436), .Z(n25323)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_587_3_lut_4_lut.init = 16'h0010;
    LUT4 equal_153_i6_1_lut_rep_595_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(clk_c_enable_205)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam equal_153_i6_1_lut_rep_595_2_lut_3_lut.init = 16'h0101;
    LUT4 counter_hi_2__bdd_4_lut_22001 (.A(mie[6]), .B(mie[14]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n24257)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam counter_hi_2__bdd_4_lut_22001.init = 16'hcac0;
    LUT4 i1_3_lut_adj_233 (.A(\mie[0] ), .B(n17061), .C(n8_adj_2353), 
         .Z(n795)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_233.init = 16'hcece;
    LUT4 counter_hi_2__bdd_3_lut (.A(n25408), .B(mie[9]), .C(mie[1]), 
         .Z(n24577)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam counter_hi_2__bdd_3_lut.init = 16'he4e4;
    LUT4 counter_hi_2__bdd_4_lut (.A(n25408), .B(mie[5]), .C(mie[13]), 
         .D(counter_hi[3]), .Z(n24576)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;
    defparam counter_hi_2__bdd_4_lut.init = 16'h5044;
    PFUMX i22002 (.BLUT(n24258), .ALUT(n24257), .C0(counter_hi[2]), .Z(n24259));
    LUT4 i21902_2_lut_rep_640 (.A(\imm[1] ), .B(\imm[0] ), .Z(n25376)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i21902_2_lut_rep_640.init = 16'hbbbb;
    LUT4 i21904_2_lut_3_lut (.A(\imm[1] ), .B(\imm[0] ), .C(\imm[10] ), 
         .Z(n23368)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i21904_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i1_3_lut_4_lut_adj_234 (.A(mip_reg[17]), .B(mie[1]), .C(n25378), 
         .D(n82), .Z(interrupt_pending_N_1402)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(321[17:24])
    defparam i1_3_lut_4_lut_adj_234.init = 16'hfff8;
    LUT4 i1_3_lut_4_lut_adj_235 (.A(mip_reg[17]), .B(mie[1]), .C(n82), 
         .D(n25378), .Z(n5_adj_2354)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(321[17:24])
    defparam i1_3_lut_4_lut_adj_235.init = 16'hff08;
    LUT4 i1_2_lut_rep_642 (.A(mie[16]), .B(timer_interrupt), .Z(n25378)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam i1_2_lut_rep_642.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(mie[16]), .B(timer_interrupt), .C(interrupt_core), 
         .Z(n611[2])) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_236 (.A(mie[16]), .B(timer_interrupt), .C(interrupt_core), 
         .Z(n611[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam i1_2_lut_3_lut_adj_236.init = 16'h7070;
    LUT4 i11998_4_lut (.A(data_rs1_c[2]), .B(n25410), .C(\debug_branch_N_173[30] ), 
         .D(n25402), .Z(alu_a_in[2])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i11998_4_lut.init = 16'h3022;
    LUT4 i11974_2_lut_rep_652 (.A(n26610), .B(counter_hi[2]), .Z(n25388)) /* synthesis lut_function=(A (B)) */ ;
    defparam i11974_2_lut_rep_652.init = 16'h8888;
    LUT4 i12200_2_lut_rep_626_3_lut (.A(n26610), .B(counter_hi[2]), .C(n26608), 
         .Z(clk_c_enable_206)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i12200_2_lut_rep_626_3_lut.init = 16'h8080;
    LUT4 i18774_2_lut_rep_446_3_lut_4_lut (.A(n26610), .B(counter_hi[2]), 
         .C(n21036), .D(n26608), .Z(n25182)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18774_2_lut_rep_446_3_lut_4_lut.init = 16'h8000;
    LUT4 i21872_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(n25350), .D(counter_hi[4]), .Z(clk_c_enable_336)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i21872_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_3_lut_4_lut_adj_237 (.A(n26610), .B(counter_hi[2]), .C(debug_instr_valid), 
         .D(n26608), .Z(n21402)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_237.init = 16'hf7ff;
    LUT4 i16401_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(counter_hi[4]), 
         .Z(n18)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;
    defparam i16401_2_lut_3_lut.init = 16'h7878;
    LUT4 i1_2_lut_rep_591_3_lut_4_lut (.A(n26610), .B(counter_hi[2]), .C(any_additional_mem_ops), 
         .D(n26608), .Z(n25327)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_591_3_lut_4_lut.init = 16'h0800;
    LUT4 i21717_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(rst_reg_n), .D(counter_hi[4]), .Z(clk_c_enable_197)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;
    defparam i21717_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i18774_rep_126_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(n21036), .D(counter_hi[4]), .Z(n23898)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18774_rep_126_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3IX mepc_i0_i22 (.D(n658[2]), .SP(clk_c_enable_396), .CD(n9321), 
            .CK(clk_c), .Q(mepc[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i22.GSR = "DISABLED";
    FD1P3IX mepc_i0_i21 (.D(n658[1]), .SP(clk_c_enable_396), .CD(n9321), 
            .CK(clk_c), .Q(mepc[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i21.GSR = "DISABLED";
    FD1P3IX mepc_i0_i20 (.D(n658[0]), .SP(clk_c_enable_396), .CD(n9321), 
            .CK(clk_c), .Q(mepc[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i20.GSR = "DISABLED";
    LUT4 i18774_rep_125_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(n21036), .D(counter_hi[4]), .Z(n23897)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18774_rep_125_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i18774_rep_124_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(n21036), .D(counter_hi[4]), .Z(n23896)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18774_rep_124_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i18774_rep_123_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(n21036), .D(counter_hi[4]), .Z(n23895)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18774_rep_123_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 tmp_data_in_3__I_99_i2_3_lut (.A(tmp_data_in_3__N_1313[1]), .B(data_rs1_c[1]), 
         .C(n5094), .Z(tmp_data_in_3__N_1245[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_99_i2_3_lut.init = 16'hcaca;
    LUT4 i18774_rep_122_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(n21036), .D(counter_hi[4]), .Z(n23894)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18774_rep_122_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_238 (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(mcause[5]), .D(counter_hi[4]), .Z(n22604)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_238.init = 16'h8000;
    LUT4 i13_rep_653 (.A(counter_hi[3]), .B(counter_hi[2]), .C(counter_hi[4]), 
         .Z(n25389)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;
    defparam i13_rep_653.init = 16'h8181;
    LUT4 equal_3119_i8_2_lut_rep_629_3_lut (.A(n26610), .B(n26608), .C(counter_hi[2]), 
         .Z(n25365)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam equal_3119_i8_2_lut_rep_629_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_654 (.A(\imm[9] ), .B(\imm[8] ), .Z(n25390)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_654.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_239 (.A(\imm[9] ), .B(\imm[8] ), .C(\imm[4] ), 
         .D(\imm[10] ), .Z(n20584)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_239.init = 16'h0008;
    LUT4 i11862_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[30]), 
         .D(n20692), .Z(\addr_out[26] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i11862_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i11863_2_lut_rep_571_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[31]), 
         .D(n20692), .Z(n25307)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i11863_2_lut_rep_571_3_lut_4_lut.init = 16'h70f0;
    LUT4 i11861_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[29]), 
         .D(n20692), .Z(\addr_out[25] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i11861_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i1_2_lut_rep_597_3_lut (.A(\imm[9] ), .B(\imm[8] ), .C(n20692), 
         .Z(n25333)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_597_3_lut.init = 16'h8080;
    LUT4 i11860_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[28]), 
         .D(n20692), .Z(\addr_out[24] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i11860_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i11_4_lut (.A(\alu_op[0] ), .B(\alu_op[3] ), .C(\alu_op[1] ), 
         .D(\alu_op_in[2] ), .Z(n5094)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i11_4_lut.init = 16'hca0a;
    LUT4 i5653_3_lut_4_lut (.A(is_alu_imm), .B(is_alu_reg), .C(is_auipc), 
         .D(debug_instr_valid), .Z(debug_rd_3__N_1131)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(225[22:46])
    defparam i5653_3_lut_4_lut.init = 16'hfe00;
    LUT4 i4469_2_lut_3_lut (.A(is_alu_imm), .B(is_alu_reg), .C(debug_instr_valid), 
         .Z(debug_rd_3__N_1132)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(225[22:46])
    defparam i4469_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_3_lut_3_lut (.A(\imm[6] ), .B(n24259), .C(n4404), .Z(n21446)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i1_3_lut_3_lut.init = 16'h4040;
    LUT4 i1_4_lut_4_lut_adj_240 (.A(\imm[6] ), .B(n25425), .C(n40), .D(n22590), 
         .Z(n21576)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i1_4_lut_4_lut_adj_240.init = 16'h4000;
    LUT4 i21891_2_lut_rep_665 (.A(counter_hi[3]), .B(counter_hi[4]), .Z(clk_c_enable_396)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i21891_2_lut_rep_665.init = 16'h7777;
    LUT4 i1_2_lut_3_lut_adj_241 (.A(n26610), .B(counter_hi[4]), .C(\imm[6] ), 
         .Z(n20677)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut_adj_241.init = 16'h7070;
    LUT4 i21817_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), .C(rst_reg_n), 
         .Z(n9321)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam i21817_2_lut_3_lut.init = 16'h0707;
    LUT4 tmp_data_in_3__I_99_i1_3_lut (.A(tmp_data_in_3__N_1313[0]), .B(data_rs1[0]), 
         .C(n5094), .Z(tmp_data_in_3__N_1245[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_99_i1_3_lut.init = 16'hcaca;
    LUT4 i11997_4_lut (.A(data_rs1_c[1]), .B(n25410), .C(\debug_branch_N_173[29] ), 
         .D(n25402), .Z(\alu_a_in[1] )) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i11997_4_lut.init = 16'h3022;
    LUT4 i11589_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), .C(mepc[0]), 
         .Z(csr_read_3__N_1182[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i11589_2_lut_3_lut.init = 16'h7070;
    LUT4 i4452_3_lut_rep_666 (.A(debug_instr_valid), .B(is_auipc), .C(is_jal), 
         .Z(n25402)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(108[27:47])
    defparam i4452_3_lut_rep_666.init = 16'ha8a8;
    LUT4 i20819_2_lut_4_lut (.A(debug_instr_valid), .B(is_auipc), .C(is_jal), 
         .D(n25426), .Z(n23094)) /* synthesis lut_function=(A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(108[27:47])
    defparam i20819_2_lut_4_lut.init = 16'ha800;
    LUT4 i21769_2_lut_rep_668 (.A(\cycle[0] ), .B(cycle[1]), .Z(n25404)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam i21769_2_lut_rep_668.init = 16'h2222;
    LUT4 i11563_3_lut_4_lut (.A(\cycle[0] ), .B(cycle[1]), .C(n25405), 
         .D(n25428), .Z(clk_c_enable_255)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam i11563_3_lut_4_lut.init = 16'hfddd;
    LUT4 i11852_2_lut_3_lut (.A(\cycle[0] ), .B(cycle[1]), .C(tmp_data[1]), 
         .Z(debug_rd_3__N_1294[1])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam i11852_2_lut_3_lut.init = 16'h2020;
    LUT4 i11853_2_lut_3_lut (.A(\cycle[0] ), .B(cycle[1]), .C(tmp_data[2]), 
         .Z(debug_rd_3__N_1294[2])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam i11853_2_lut_3_lut.init = 16'h2020;
    LUT4 i4301_2_lut (.A(time_hi[0]), .B(clk_c_enable_170), .Z(n1[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam i4301_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_242 (.A(n25292), .B(instr_complete_N_1379), .C(n13853), 
         .D(n8720), .Z(n14111)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(220[18] 228[36])
    defparam i1_4_lut_adj_242.init = 16'hffef;
    LUT4 i1_3_lut_rep_669 (.A(\alu_op[3] ), .B(\alu_op[1] ), .C(\alu_op_in[2] ), 
         .Z(n25405)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_rep_669.init = 16'hf7f7;
    LUT4 i11634_2_lut (.A(\cycle[0] ), .B(cycle[1]), .Z(n13853)) /* synthesis lut_function=(A (B)) */ ;
    defparam i11634_2_lut.init = 16'h8888;
    LUT4 mux_3084_i4_4_lut_4_lut (.A(\imm[0] ), .B(\imm[1] ), .C(instrret_count[3]), 
         .D(cycle_count_wide[3]), .Z(n4994[3])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam mux_3084_i4_4_lut_4_lut.init = 16'h7340;
    LUT4 imm_3__I_0_i2_3_lut (.A(\debug_rd_3__N_136[29] ), .B(data_rs2[1]), 
         .C(alu_b_in_3__N_1235), .Z(\alu_b_in[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 mux_3084_i3_4_lut_4_lut (.A(\imm[0] ), .B(\imm[1] ), .C(instrret_count[2]), 
         .D(cycle_count_wide_c[2]), .Z(n4996)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam mux_3084_i3_4_lut_4_lut.init = 16'h7340;
    LUT4 i1_3_lut_rep_672 (.A(n26610), .B(counter_hi[2]), .C(counter_hi[4]), 
         .Z(n25408)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;
    defparam i1_3_lut_rep_672.init = 16'h1414;
    LUT4 i21915_2_lut_rep_615_3_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(counter_hi[4]), .Z(n25351)) /* synthesis lut_function=(!(A (B)+!A (B (C)))) */ ;
    defparam i21915_2_lut_rep_615_3_lut.init = 16'h3737;
    LUT4 i1_4_lut_adj_243 (.A(\imm[1] ), .B(n25425), .C(\imm[0] ), .D(\imm[2] ), 
         .Z(n8500)) /* synthesis lut_function=(!(A+((C (D)+!C !(D))+!B))) */ ;
    defparam i1_4_lut_adj_243.init = 16'h0440;
    LUT4 i4264_2_lut (.A(\imm[6] ), .B(\imm[1] ), .Z(n6452)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i4264_2_lut.init = 16'h6666;
    LUT4 i1_2_lut_adj_244 (.A(\imm[2] ), .B(\imm[10] ), .Z(n22590)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_244.init = 16'h4444;
    LUT4 i67_4_lut (.A(n13929), .B(n25390), .C(\imm[4] ), .D(n25436), 
         .Z(n40)) /* synthesis lut_function=(A (B (C))+!A !(C+(D))) */ ;
    defparam i67_4_lut.init = 16'h8085;
    LUT4 i11710_2_lut (.A(\imm[1] ), .B(\imm[0] ), .Z(n13929)) /* synthesis lut_function=(A (B)) */ ;
    defparam i11710_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_rep_674 (.A(\alu_op[1] ), .B(\alu_op_in[2] ), .C(\alu_op[3] ), 
         .Z(n25410)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_674.init = 16'h8080;
    LUT4 i1_3_lut_adj_245 (.A(\alu_op_in[2] ), .B(\alu_op[1] ), .C(\alu_op[3] ), 
         .Z(n8461)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(64[33:56])
    defparam i1_3_lut_adj_245.init = 16'hfbfb;
    LUT4 i4295_2_lut_rep_518_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in[0]), .Z(n25254)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i4295_2_lut_rep_518_4_lut_4_lut.init = 16'h857a;
    LUT4 i11731_3_lut_rep_616_3_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .Z(n25352)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;
    defparam i11731_3_lut_rep_616_3_lut.init = 16'h7a7a;
    LUT4 i4297_2_lut_rep_514_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in_c[2]), .Z(n25250)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i4297_2_lut_rep_514_4_lut_4_lut.init = 16'h857a;
    LUT4 i4296_2_lut_rep_515_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in_c[3]), .Z(n25251)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i4296_2_lut_rep_515_4_lut_4_lut.init = 16'h857a;
    LUT4 i12199_1_lut_rep_631_3_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .Z(n25367)) /* synthesis lut_function=(!(A (B (C)))) */ ;
    defparam i12199_1_lut_rep_631_3_lut.init = 16'h7f7f;
    LUT4 i4298_2_lut_rep_538_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(\alu_b_in[1] ), .Z(n25274)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i4298_2_lut_rep_538_4_lut_4_lut.init = 16'h857a;
    LUT4 i11849_2_lut_rep_621_3_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .Z(n25357)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i11849_2_lut_rep_621_3_lut.init = 16'h2a2a;
    LUT4 i11539_2_lut_rep_622_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(\alu_op[0] ), .Z(n25358)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;
    defparam i11539_2_lut_rep_622_4_lut.init = 16'h7f00;
    PFUMX i22006 (.BLUT(n24265), .ALUT(n24264), .C0(counter_hi[4]), .Z(n24266));
    LUT4 is_jal_I_0_2_lut_rep_676 (.A(is_jal), .B(is_jalr), .Z(n25412)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam is_jal_I_0_2_lut_rep_676.init = 16'heeee;
    LUT4 i21120_2_lut_3_lut_4_lut (.A(is_jal), .B(is_jalr), .C(n25426), 
         .D(debug_instr_valid), .Z(n23395)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam i21120_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i4462_2_lut_rep_623_3_lut (.A(is_jal), .B(is_jalr), .C(debug_instr_valid), 
         .Z(n25359)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam i4462_2_lut_rep_623_3_lut.init = 16'he0e0;
    LUT4 i21921_2_lut_3_lut_3_lut_4_lut (.A(is_jal), .B(is_jalr), .C(debug_instr_valid), 
         .D(is_lui), .Z(n23325)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam i21921_2_lut_3_lut_3_lut_4_lut.init = 16'hff1f;
    LUT4 i21906_2_lut_rep_677 (.A(\imm[10] ), .B(\imm[1] ), .Z(n25413)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i21906_2_lut_rep_677.init = 16'hdddd;
    LUT4 i21447_3_lut_4_lut (.A(\imm[10] ), .B(\imm[1] ), .C(n24695), 
         .D(n23001), .Z(n5041[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i21447_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i1_2_lut_rep_636_3_lut (.A(n26610), .B(n26608), .C(counter_hi[2]), 
         .Z(n25372)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_636_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_adj_246 (.A(n26608), .B(counter_hi[2]), .C(counter_hi[3]), 
         .Z(n4404)) /* synthesis lut_function=(A+!((C)+!B)) */ ;
    defparam i1_3_lut_adj_246.init = 16'haeae;
    LUT4 equal_3123_i6_2_lut_rep_685 (.A(\cycle[0] ), .B(cycle[1]), .Z(n25421)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(57[23:37])
    defparam equal_3123_i6_2_lut_rep_685.init = 16'heeee;
    LUT4 i21786_2_lut_3_lut_4_lut (.A(\cycle[0] ), .B(cycle[1]), .C(counter_hi[2]), 
         .D(n25435), .Z(clk_c_enable_161)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(57[23:37])
    defparam i21786_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_3_lut_4_lut_adj_247 (.A(\cycle[0] ), .B(cycle[1]), .C(is_load), 
         .D(is_store), .Z(n5_adj_1)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(57[23:37])
    defparam i1_2_lut_3_lut_4_lut_adj_247.init = 16'h1110;
    LUT4 i21863_2_lut_3_lut_4_lut (.A(\cycle[0] ), .B(cycle[1]), .C(n25435), 
         .D(counter_hi[2]), .Z(clk_c_enable_158)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(57[23:37])
    defparam i21863_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 n24279_bdd_3_lut (.A(n24279), .B(load_top_bit), .C(data_out_3__N_1116), 
         .Z(n24280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24279_bdd_3_lut.init = 16'hcaca;
    LUT4 i11566_2_lut (.A(data_rs2[0]), .B(data_out_3__N_1116), .Z(\data_out_slice[0] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i11566_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_248 (.A(n25273), .B(n22937), .C(n25296), .D(n14477), 
         .Z(clk_c_enable_162)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i1_4_lut_adj_248.init = 16'hfbfa;
    LUT4 i20721_4_lut (.A(n25333), .B(n25309), .C(n25365), .D(\imm[2] ), 
         .Z(n22937)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20721_4_lut.init = 16'hfffe;
    LUT4 i11477_4_lut (.A(n25270), .B(n25273), .C(mstatus_mie), .D(n25296), 
         .Z(n5400)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam i11477_4_lut.init = 16'h3022;
    LUT4 debug_branch_N_571_29__bdd_3_lut_22279 (.A(\debug_branch_N_571[29] ), 
         .B(\timer_data[1] ), .C(is_timer_addr), .Z(n24279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam debug_branch_N_571_29__bdd_3_lut_22279.init = 16'hcaca;
    LUT4 i21858_2_lut_rep_689 (.A(\imm[5] ), .B(\imm[3] ), .Z(n25425)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21858_2_lut_rep_689.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_adj_249 (.A(\imm[5] ), .B(\imm[3] ), .C(\imm[4] ), 
         .Z(n16)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut_adj_249.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut_adj_250 (.A(\imm[5] ), .B(\imm[3] ), .C(\imm[2] ), 
         .D(\imm[0] ), .Z(n22602)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_250.init = 16'hfffe;
    LUT4 i4453_3_lut (.A(debug_instr_valid), .B(is_alu_reg), .C(is_branch), 
         .Z(alu_b_in_3__N_1235)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:52])
    defparam i4453_3_lut.init = 16'ha8a8;
    LUT4 i11866_2_lut_rep_541 (.A(data_rs2[3]), .B(data_out_3__N_1116), 
         .Z(n25277)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i11866_2_lut_rep_541.init = 16'h2222;
    LUT4 i3731_3_lut (.A(time_hi[2]), .B(time_hi[1]), .C(time_hi[0]), 
         .Z(n498[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(295[55:71])
    defparam i3731_3_lut.init = 16'h6a6a;
    LUT4 i3724_2_lut (.A(time_hi[1]), .B(time_hi[0]), .Z(n498[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(295[55:71])
    defparam i3724_2_lut.init = 16'h6666;
    LUT4 debug_rd_3__N_1298_1__bdd_4_lut (.A(n196[1]), .B(debug_rd_3__N_1294[1]), 
         .C(n25410), .D(n15), .Z(n24278)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam debug_rd_3__N_1298_1__bdd_4_lut.init = 16'hcac0;
    LUT4 equal_3122_i6_2_lut_rep_692 (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .Z(n25428)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam equal_3122_i6_2_lut_rep_692.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_251 (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .C(mip_reg[16]), .D(n25369), .Z(n22674)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i1_2_lut_3_lut_4_lut_adj_251.init = 16'hd0f0;
    LUT4 equal_3122_i7_2_lut_rep_630_3_lut_4_lut (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .C(cycle[1]), .D(\cycle[0] ), .Z(n25366)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam equal_3122_i7_2_lut_rep_630_3_lut_4_lut.init = 16'hfdff;
    LUT4 i1_3_lut_adj_252 (.A(mie[14]), .B(n12484), .C(n8_adj_2356), .Z(n926)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_252.init = 16'hcece;
    LUT4 i12247_3_lut_4_lut_4_lut_4_lut (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .C(\data_rs1[3] ), .D(n25369), .Z(n14477)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i12247_3_lut_4_lut_4_lut_4_lut.init = 16'he200;
    L6MUX21 instr_complete_I_106 (.D0(instr_complete_N_1381), .D1(instr_complete_N_1380), 
            .SD(n23111), .Z(instr_complete_N_1379)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_adj_253 (.A(mie[12]), .B(n17061), .C(n8_adj_2353), .Z(n928)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_253.init = 16'hcece;
    LUT4 i1_4_lut_adj_254 (.A(n25375), .B(n25295), .C(n25365), .D(n22798), 
         .Z(clk_c_enable_184)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(429[18] 459[12])
    defparam i1_4_lut_adj_254.init = 16'h2000;
    LUT4 i1_3_lut_adj_255 (.A(mie[10]), .B(n12484), .C(n8_adj_2356), .Z(n893)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_255.init = 16'hcece;
    PFUMX instr_complete_I_107 (.BLUT(instr_complete_N_1385), .ALUT(instr_complete_N_1387), 
          .C0(n25387), .Z(instr_complete_N_1380)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_adj_256 (.A(\mie[8] ), .B(n17061), .C(n8_adj_2353), 
         .Z(n895)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_256.init = 16'hcece;
    LUT4 imm_3__I_0_i4_3_lut (.A(\debug_rd_3__N_136[31] ), .B(data_rs2[3]), 
         .C(alu_b_in_3__N_1235), .Z(alu_b_in_c[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i4_3_lut.init = 16'hcaca;
    PFUMX tmp_data_in_3__I_0_i4 (.BLUT(tmp_data_in_3__N_1313[3]), .ALUT(\tmp_data_in_3__N_1245[3] ), 
          .C0(n23334), .Z(tmp_data_in[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i353_4_lut (.A(n39), .B(data_rs1_c[2]), .C(n25343), .D(n25319), 
         .Z(n860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(444[22] 445[73])
    defparam i353_4_lut.init = 16'hceca;
    PFUMX debug_rd_3__I_96_i3 (.BLUT(debug_rd_3__N_1294[2]), .ALUT(debug_rd_3__N_1290[2]), 
          .C0(n25367), .Z(debug_rd_3__N_1127[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 imm_3__I_0_i3_3_lut (.A(\debug_rd_3__N_136[30] ), .B(data_rs2[2]), 
         .C(alu_b_in_3__N_1235), .Z(alu_b_in_c[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_257 (.A(mie[4]), .B(n17061), .C(n8_adj_2353), .Z(n862)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_257.init = 16'hcece;
    LUT4 n24281_bdd_3_lut (.A(n24281), .B(n24278), .C(debug_rd_3__N_1131), 
         .Z(debug_rd[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24281_bdd_3_lut.init = 16'hcaca;
    LUT4 tmp_data_31__I_0_542_i10_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[9]), 
         .D(tmp_data[13]), .Z(\addr_out[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i11999_4_lut (.A(\data_rs1[3] ), .B(n25410), .C(\debug_branch_N_173[31] ), 
         .D(n25402), .Z(alu_a_in[3])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i11999_4_lut.init = 16'h3022;
    PFUMX tmp_data_in_3__I_0_i3 (.BLUT(tmp_data_in_3__N_1313[2]), .ALUT(tmp_data_in_3__N_1245[2]), 
          .C0(n23334), .Z(tmp_data_in[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_4_lut_adj_258 (.A(n25301), .B(\data_rs1[3] ), .C(n20), 
         .D(mie[16]), .Z(n20019)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_258.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_259 (.A(n25301), .B(\data_rs1[3] ), .C(n22935), 
         .D(mie[15]), .Z(n925)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_259.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_260 (.A(n25301), .B(\data_rs1[3] ), .C(n22935), 
         .D(mie[11]), .Z(n892)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_260.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_261 (.A(n25301), .B(\data_rs1[3] ), .C(n22935), 
         .D(mie[7]), .Z(n859)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_261.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_262 (.A(n25301), .B(\data_rs1[3] ), .C(n20), 
         .D(mie[3]), .Z(n20021)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_262.init = 16'h8f88;
    LUT4 i40_3_lut_4_lut (.A(n25301), .B(\data_rs1[3] ), .C(n25333), .D(mstatus_mpie), 
         .Z(n33)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i40_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_3_lut_adj_263 (.A(mie[2]), .B(n12484), .C(n8_adj_2356), .Z(n793)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_263.init = 16'hcece;
    LUT4 i1_4_lut_adj_264 (.A(n8448), .B(n25344), .C(\debug_rd_3__N_136[28] ), 
         .D(interrupt_core), .Z(n21695)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_264.init = 16'h0004;
    LUT4 i1_3_lut_adj_265 (.A(\debug_rd_3__N_136[30] ), .B(\debug_rd_3__N_136[29] ), 
         .C(\debug_rd_3__N_136[31] ), .Z(n8448)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(353[26:40])
    defparam i1_3_lut_adj_265.init = 16'hfefe;
    PFUMX debug_rd_3__I_97_i1 (.BLUT(\debug_rd_3__N_1298[0] ), .ALUT(debug_rd_3__N_1302[0]), 
          .C0(debug_rd_3__N_1306), .Z(debug_rd_3__N_1123[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX debug_rd_3__I_96_i1 (.BLUT(shift_out[0]), .ALUT(debug_rd_3__N_1290[0]), 
          .C0(n23385), .Z(debug_rd_3__N_1127[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_4_lut_adj_266 (.A(rst_reg_n), .B(n25293), .C(n33), .D(n25296), 
         .Z(mstatus_mie_N_1438)) /* synthesis lut_function=((B+!((D)+!C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(395[13:37])
    defparam i1_3_lut_4_lut_adj_266.init = 16'hddfd;
    LUT4 i1_3_lut_4_lut_adj_267 (.A(rst_reg_n), .B(n25293), .C(n25365), 
         .D(n11558), .Z(clk_c_enable_280)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(395[13:37])
    defparam i1_3_lut_4_lut_adj_267.init = 16'h2000;
    LUT4 i11957_2_lut_3_lut_4_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(csr_read_3__N_1174[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i11957_2_lut_3_lut_4_lut_3_lut.init = 16'h1010;
    LUT4 i21838_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_top_bit_next_N_1462), .D(counter_hi[2]), .Z(n14438)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i21838_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i7_3_lut (.A(mie[4]), .B(mie[12]), .C(counter_hi[3]), .Z(n3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(139[15:25])
    defparam i7_3_lut.init = 16'hcaca;
    LUT4 i3296_2_lut_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(mstatus_mte), .D(counter_hi[2]), .Z(n5287)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3296_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_top_bit_next_N_1462), .D(counter_hi[2]), .Z(clk_c_enable_359)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i11737_2_lut_rep_579_2_lut_3_lut_4_lut (.A(n26610), .B(n26608), 
         .C(cy_adj_3), .D(counter_hi[2]), .Z(n25315)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;
    defparam i11737_2_lut_rep_579_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i12051_2_lut_rep_700 (.A(\imm[8] ), .B(\imm[9] ), .Z(n25436)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12051_2_lut_rep_700.init = 16'heeee;
    LUT4 i1_2_lut_rep_608_3_lut (.A(\imm[8] ), .B(\imm[9] ), .C(n20692), 
         .Z(n25344)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_608_3_lut.init = 16'h1010;
    LUT4 is_trap_I_0_586_2_lut_rep_580_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), 
         .C(interrupt_core), .D(n20692), .Z(n25316)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam is_trap_I_0_586_2_lut_rep_580_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i1_2_lut_rep_570_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), .C(interrupt_core), 
         .D(n20692), .Z(n25306)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i1_2_lut_rep_570_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i11574_2_lut_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), .C(n8448), 
         .D(n20692), .Z(n4495[0])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i11574_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 mtimecmp_7__I_0_3_lut_4_lut (.A(data_rs2[3]), .B(data_out_3__N_1116), 
         .C(n25282), .D(\mtimecmp[7] ), .Z(mtimecmp_3__N_1666)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam mtimecmp_7__I_0_3_lut_4_lut.init = 16'h2f20;
    LUT4 i11865_2_lut (.A(data_rs2[2]), .B(data_out_3__N_1116), .Z(\data_out_slice[2] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i11865_2_lut.init = 16'h2222;
    LUT4 debug_rd_3__I_0_i3_4_lut (.A(debug_rd_3__N_1302[2]), .B(debug_rd_3__N_1123[2]), 
         .C(debug_rd_3__N_1131), .D(debug_rd_3__N_1306), .Z(debug_rd[2])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(176[18] 194[12])
    defparam debug_rd_3__I_0_i3_4_lut.init = 16'hcacc;
    LUT4 i6466_4_lut (.A(debug_instr_valid), .B(n22450), .C(is_lui), .D(is_jal), 
         .Z(n8720)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(218[17:110])
    defparam i6466_4_lut.init = 16'haaa8;
    LUT4 mux_87_i3_3_lut (.A(n24932), .B(\debug_branch_N_181[2] ), .C(n23306), 
         .Z(debug_rd_3__N_1302[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam mux_87_i3_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_268 (.A(is_branch), .B(is_jalr), .C(is_auipc), .D(is_system), 
         .Z(n22450)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(218[17:110])
    defparam i1_4_lut_adj_268.init = 16'hfffe;
    LUT4 i21925_3_lut (.A(data_out_3__N_1116), .B(is_timer_addr), .C(n26608), 
         .Z(n23306)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam i21925_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_adj_269 (.A(interrupt_pending_N_1402), .B(no_write_in_progress), 
         .C(mstatus_mie), .Z(n21786)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_adj_269.init = 16'h8080;
    LUT4 i1_3_lut_4_lut_adj_270 (.A(data_rs1_c[1]), .B(n25301), .C(n20_adj_2357), 
         .D(mie[1]), .Z(n20023)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(450[22] 451[75])
    defparam i1_3_lut_4_lut_adj_270.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_271 (.A(data_rs1_c[1]), .B(n25301), .C(n20_adj_2357), 
         .D(mie[13]), .Z(n20033)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(450[22] 451[75])
    defparam i1_3_lut_4_lut_adj_271.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_272 (.A(data_rs1_c[1]), .B(n25301), .C(n20_adj_2357), 
         .D(mie[9]), .Z(n20031)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(450[22] 451[75])
    defparam i1_3_lut_4_lut_adj_272.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_273 (.A(data_rs1_c[1]), .B(n25301), .C(n20_adj_2357), 
         .D(mie[5]), .Z(n20029)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(450[22] 451[75])
    defparam i1_3_lut_4_lut_adj_273.init = 16'h8f88;
    PFUMX mux_443_i1 (.BLUT(n822[0]), .ALUT(n948[0]), .C0(n25348), .Z(n979[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_4_lut_adj_274 (.A(n25306), .B(n25326), .C(n8720), .D(instr_complete_N_1379), 
         .Z(instr_complete_N_1378)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i1_3_lut_4_lut_adj_274.init = 16'hfffe;
    LUT4 rstn_N_1310_I_0_2_lut_rep_537_4_lut (.A(mstatus_mte), .B(is_double_fault_r), 
         .C(n25323), .D(rst_reg_n), .Z(n25273)) /* synthesis lut_function=(A (B+!(D))+!A (B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(365[28:90])
    defparam rstn_N_1310_I_0_2_lut_rep_537_4_lut.init = 16'hdcff;
    LUT4 i1_2_lut_4_lut_adj_275 (.A(mstatus_mte), .B(is_double_fault_r), 
         .C(n25323), .D(n25296), .Z(mstatus_mte_N_1434)) /* synthesis lut_function=(A (B+!(D))+!A (B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(365[28:90])
    defparam i1_2_lut_4_lut_adj_275.init = 16'hdcff;
    LUT4 mux_93_i2_3_lut (.A(n23069), .B(n234[1]), .C(n23322), .Z(debug_rd_3__N_1298[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(187[18] 194[12])
    defparam mux_93_i2_3_lut.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_4_lut_adj_276 (.A(\imm[2] ), .B(n25309), .C(clk_c_enable_206), 
         .D(n25365), .Z(clk_c_enable_180)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i1_2_lut_3_lut_4_lut_adj_276.init = 16'h2000;
    PFUMX i20802 (.BLUT(time_count[3]), .ALUT(n4994[3]), .C0(n25376), 
          .Z(n23077));
    LUT4 i2_2_lut_3_lut_4_lut (.A(\imm[2] ), .B(n25309), .C(n11558), .D(n25365), 
         .Z(clk_c_enable_189)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_277 (.A(\imm[2] ), .B(n25309), .C(n25348), 
         .D(n25365), .Z(clk_c_enable_190)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i1_2_lut_3_lut_4_lut_adj_277.init = 16'h0200;
    LUT4 i101_2_lut (.A(mip_reg[16]), .B(\mie[0] ), .Z(n82)) /* synthesis lut_function=(A (B)) */ ;
    defparam i101_2_lut.init = 16'h8888;
    LUT4 tmp_data_31__I_0_542_i2_3_lut_4_lut (.A(n25390), .B(n20692), .C(mepc[1]), 
         .D(tmp_data[5]), .Z(\addr_out[1] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_278 (.A(n14329), .B(debug_rd_3__N_1306), .C(mem_op[1]), 
         .D(mem_op[2]), .Z(load_top_bit_next_N_1462)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_278.init = 16'h0004;
    LUT4 mux_87_i4_3_lut_4_lut (.A(data_out_3__N_1116), .B(is_timer_addr), 
         .C(n22944), .D(\debug_branch_N_571[31] ), .Z(debug_rd_3__N_1302[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam mux_87_i4_3_lut_4_lut.init = 16'hf1e0;
    PFUMX mux_91_i4 (.BLUT(n23073), .ALUT(\debug_branch_N_177[31] ), .C0(n23325), 
          .Z(n234[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 dr_3__N_1595_32__bdd_3_lut_22351 (.A(alu_out[2]), .B(\mul_out[2] ), 
         .C(n25405), .Z(n24863)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam dr_3__N_1595_32__bdd_3_lut_22351.init = 16'hacac;
    PFUMX mux_91_i2 (.BLUT(n23067), .ALUT(\debug_branch_N_177[29] ), .C0(n23325), 
          .Z(n234[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 next_pc_for_core_22__bdd_3_lut_23107 (.A(\next_pc_for_core[14] ), 
         .B(\next_pc_for_core[10] ), .C(counter_hi[2]), .Z(n25653)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam next_pc_for_core_22__bdd_3_lut_23107.init = 16'hacac;
    LUT4 i21741_3_lut_4_lut (.A(n25344), .B(interrupt_core), .C(n25372), 
         .D(rst_reg_n), .Z(clk_c_enable_279)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i21741_3_lut_4_lut.init = 16'h0eff;
    LUT4 i10016_3_lut_4_lut (.A(tmp_data[31]), .B(n25333), .C(n5_adj_1), 
         .D(n66), .Z(n12257)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(267[23:65])
    defparam i10016_3_lut_4_lut.init = 16'h2f20;
    LUT4 debug_rd_3__N_1306_bdd_4_lut_22600 (.A(n25369), .B(n25412), .C(debug_instr_valid), 
         .D(is_lui), .Z(n24883)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam debug_rd_3__N_1306_bdd_4_lut_22600.init = 16'hfaea;
    LUT4 dr_3__N_1595_32__bdd_3_lut_22610 (.A(dr_3__N_1595[32]), .B(dr_3__N_1595[33]), 
         .C(\alu_op_in[2] ), .Z(n24864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam dr_3__N_1595_32__bdd_3_lut_22610.init = 16'hcaca;
    LUT4 i1_2_lut_rep_573 (.A(\imm[6] ), .B(n20561), .Z(n25309)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam i1_2_lut_rep_573.init = 16'heeee;
    LUT4 i21738_2_lut_3_lut_4_lut (.A(\imm[6] ), .B(n20561), .C(n25365), 
         .D(\imm[2] ), .Z(clk_c_enable_176)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam i21738_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_559_3_lut (.A(\imm[6] ), .B(n20561), .C(\imm[2] ), 
         .Z(n25295)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam i1_2_lut_rep_559_3_lut.init = 16'hefef;
    LUT4 i20712_3_lut_4_lut (.A(\imm[6] ), .B(n20561), .C(\imm[2] ), .D(n25372), 
         .Z(n22927)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam i20712_3_lut_4_lut.init = 16'hfffe;
    LUT4 i3582_2_lut_4_lut (.A(tmp_data[6]), .B(mepc[2]), .C(n25333), 
         .D(\addr_offset[2] ), .Z(n701)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(267[23:65])
    defparam i3582_2_lut_4_lut.init = 16'h35ca;
    LUT4 n24883_bdd_2_lut (.A(n24883), .B(debug_rd_3__N_1306), .Z(n24884)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n24883_bdd_2_lut.init = 16'heeee;
    PFUMX mux_443_i2 (.BLUT(n822[1]), .ALUT(n948[1]), .C0(n25348), .Z(n979[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX mux_91_i3 (.BLUT(n23070), .ALUT(\debug_branch_N_177[30] ), .C0(n23325), 
          .Z(n234[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 mux_252_i3_3_lut_4_lut (.A(n25344), .B(interrupt_core), .C(\debug_branch_N_173[30] ), 
         .D(n653[2]), .Z(n658[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i2_3_lut_4_lut (.A(n25344), .B(interrupt_core), .C(\debug_branch_N_173[29] ), 
         .D(n653[1]), .Z(n658[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i4_3_lut_4_lut (.A(n25344), .B(interrupt_core), .C(\debug_branch_N_173[31] ), 
         .D(n653[3]), .Z(n658[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i4_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i22739 (.D0(n25850), .D1(n25848), .SD(debug_rd_3__N_1131), 
            .Z(debug_rd[3]));
    PFUMX i22737 (.BLUT(n25849), .ALUT(debug_rd_3__N_1302[3]), .C0(debug_rd_3__N_1306), 
          .Z(n25850));
    PFUMX i22735 (.BLUT(n25847), .ALUT(n25846), .C0(n25410), .Z(n25848));
    LUT4 debug_rd_3__N_1306_bdd_4_lut_22363 (.A(\alu_op[3] ), .B(\alu_op[1] ), 
         .C(\alu_op_in[2] ), .D(\cycle[0] ), .Z(n24882)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam debug_rd_3__N_1306_bdd_4_lut_22363.init = 16'hfff7;
    LUT4 data_rs1_3__I_0_i1_2_lut (.A(data_rs1[0]), .B(\cycle[0] ), .Z(mul_out_3__N_1241[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i1_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i2_2_lut (.A(data_rs1_c[1]), .B(\cycle[0] ), .Z(mul_out_3__N_1241[1])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i2_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i3_2_lut (.A(data_rs1_c[2]), .B(\cycle[0] ), .Z(mul_out_3__N_1241[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i3_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i4_2_lut (.A(\data_rs1[3] ), .B(\cycle[0] ), .Z(mul_out_3__N_1241[3])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i4_2_lut.init = 16'h8888;
    LUT4 i7000_2_lut_rep_534_3_lut_4_lut (.A(\alu_op[0] ), .B(n25341), .C(\data_rs1[3] ), 
         .D(n25343), .Z(n25270)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i7000_2_lut_rep_534_3_lut_4_lut.init = 16'hf040;
    PFUMX i20805 (.BLUT(csr_read_3__N_1174[0]), .ALUT(csr_read_3__N_1182[0]), 
          .C0(\imm[6] ), .Z(n23080));
    LUT4 i1_2_lut_3_lut_4_lut_adj_279 (.A(\alu_op[0] ), .B(n25341), .C(data_rs1_c[2]), 
         .D(n25343), .Z(n12484)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_279.init = 16'hf040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_280 (.A(\alu_op[0] ), .B(n25341), .C(data_rs1[0]), 
         .D(n25343), .Z(n17061)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_280.init = 16'hf040;
    LUT4 mux_251_i4_3_lut (.A(mepc[3]), .B(\data_rs1[3] ), .C(n652), .Z(n653[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i4_3_lut.init = 16'hcaca;
    LUT4 i25_3_lut_4_lut (.A(\alu_op[0] ), .B(n25341), .C(data_rs1_c[1]), 
         .D(n25343), .Z(n20_adj_2357)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i25_3_lut_4_lut.init = 16'h8f80;
    LUT4 i20719_3_lut_4_lut (.A(\alu_op[0] ), .B(n25341), .C(\data_rs1[3] ), 
         .D(n25343), .Z(n22935)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i20719_3_lut_4_lut.init = 16'hff80;
    LUT4 i1_4_lut_adj_281 (.A(n18_c), .B(n25343), .C(n21), .D(n22782), 
         .Z(n652)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_281.init = 16'h0400;
    LUT4 i1_4_lut_adj_282 (.A(\imm[2] ), .B(n16), .C(\imm[1] ), .D(n22776), 
         .Z(n22782)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_282.init = 16'h0100;
    LUT4 i1_2_lut_adj_283 (.A(\imm[0] ), .B(\imm[6] ), .Z(n22776)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_283.init = 16'h8888;
    LUT4 i13_3_lut_4_lut (.A(\alu_op[0] ), .B(n25341), .C(data_rs1[0]), 
         .D(n25343), .Z(n8_adj_2353)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i25_3_lut_4_lut_adj_284 (.A(\alu_op[0] ), .B(n25341), .C(\data_rs1[3] ), 
         .D(n25343), .Z(n20)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i25_3_lut_4_lut_adj_284.init = 16'h8f80;
    LUT4 i13_3_lut_4_lut_adj_285 (.A(\alu_op[0] ), .B(n25341), .C(data_rs1_c[2]), 
         .D(n25343), .Z(n8_adj_2356)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i13_3_lut_4_lut_adj_285.init = 16'h8f80;
    LUT4 i1_3_lut_4_lut_adj_286 (.A(\alu_op[0] ), .B(n25341), .C(mie[6]), 
         .D(data_rs1_c[2]), .Z(n39)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i1_3_lut_4_lut_adj_286.init = 16'h70f0;
    LUT4 i1_4_lut_adj_287 (.A(\cycle[0] ), .B(n8461), .C(n25405), .D(n25428), 
         .Z(instr_complete_N_1383)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam i1_4_lut_adj_287.init = 16'h6aaa;
    LUT4 i1_4_lut_adj_288 (.A(n25273), .B(n22927), .C(n25271), .D(n14477), 
         .Z(clk_c_enable_320)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i1_4_lut_adj_288.init = 16'hfbfa;
    LUT4 is_double_fault_I_0_3_lut_rep_557_4_lut (.A(n25372), .B(n25344), 
         .C(is_double_fault_r), .D(mstatus_mte), .Z(n25293)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;
    defparam is_double_fault_I_0_3_lut_rep_557_4_lut.init = 16'hf0f4;
    PFUMX mux_252_i1 (.BLUT(n653[0]), .ALUT(n22939), .C0(n25316), .Z(n658[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX mux_3109_i2 (.BLUT(n5041[1]), .ALUT(n5035[1]), .C0(n5040), .Z(n5047[1]));
    LUT4 i1_4_lut_adj_289 (.A(n8500), .B(n20584), .C(n22602), .D(n6452), 
         .Z(n20586)) /* synthesis lut_function=(A (B)+!A !((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_289.init = 16'h888c;
    LUT4 i1_3_lut_rep_445_4_lut (.A(clk_c_enable_206), .B(any_additional_mem_ops), 
         .C(instr_complete_N_1378), .D(n25349), .Z(n25181)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_rep_445_4_lut.init = 16'h0020;
    L6MUX21 i20803 (.D0(n23076), .D1(n23077), .SD(\imm[10] ), .Z(n23078));
    L6MUX21 i20806 (.D0(n23079), .D1(n23080), .SD(\imm[0] ), .Z(n23081));
    L6MUX21 i22628 (.D0(n234[2]), .D1(n25654), .SD(n23322), .Z(n25655));
    PFUMX i22626 (.BLUT(n25653), .ALUT(n25652), .C0(counter_hi[4]), .Z(n25654));
    L6MUX21 mux_3109_i3 (.D0(n5041[2]), .D1(n5035[2]), .SD(n5040), .Z(n5047[2]));
    PFUMX mux_3107_i1 (.BLUT(n23010), .ALUT(n23012), .C0(n25413), .Z(n5041[0]));
    PFUMX i22545 (.BLUT(n25473), .ALUT(n25474), .C0(counter_hi[2]), .Z(n25475));
    PFUMX mux_233_i1 (.BLUT(n4495[0]), .ALUT(n5_adj_2354), .C0(interrupt_core), 
          .Z(n611[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX mux_3089_i2 (.BLUT(csr_read_3__N_1178[1]), .ALUT(csr_read_3__N_1190[1]), 
          .C0(\imm[6] ), .Z(n5003[1]));
    PFUMX i22537 (.BLUT(n25459), .ALUT(n25460), .C0(data_rs1_c[1]), .Z(n25461));
    PFUMX mux_3105_i3 (.BLUT(n21446), .ALUT(n5013[2]), .C0(\imm[0] ), 
          .Z(n5035[2]));
    PFUMX i20804 (.BLUT(csr_read_3__N_1178[0]), .ALUT(csr_read_3__N_1190[0]), 
          .C0(\imm[6] ), .Z(n23079));
    PFUMX i20801 (.BLUT(\csr_read_3__N_1170[3] ), .ALUT(csr_read_3__N_1186[3]), 
          .C0(\imm[1] ), .Z(n23076));
    tinyqv_mul multiplier (.accum({accum}), .\next_accum[6] (\next_accum[6] ), 
            .\next_accum[7] (\next_accum[7] ), .\next_accum[8] (\next_accum[8] ), 
            .\next_accum[9] (\next_accum[9] ), .\next_accum[10] (\next_accum[10] ), 
            .\next_accum[11] (\next_accum[11] ), .\next_accum[12] (\next_accum[12] ), 
            .\next_accum[13] (\next_accum[13] ), .\next_accum[14] (\next_accum[14] ), 
            .\next_accum[15] (\next_accum[15] ), .clk_c(clk_c), .mul_out_3__N_1241({mul_out_3__N_1241}), 
            .\tmp_data[0] (tmp_data[0]), .\tmp_data[1] (tmp_data[1]), .\tmp_data[2] (tmp_data[2]), 
            .\tmp_data[3] (tmp_data[3]), .\tmp_data[4] (tmp_data[4]), .\tmp_data[5] (tmp_data[5]), 
            .\tmp_data[6] (tmp_data[6]), .\tmp_data[7] (tmp_data[7]), .\tmp_data[8] (tmp_data[8]), 
            .\tmp_data[9] (tmp_data[9]), .\tmp_data[10] (tmp_data[10]), 
            .\tmp_data[11] (tmp_data[11]), .\tmp_data[12] (tmp_data[12]), 
            .\tmp_data[13] (tmp_data[13]), .\tmp_data[14] (tmp_data[14]), 
            .\tmp_data[15] (tmp_data[15]), .d_3__N_1599({d_3__N_1599}), 
            .GND_net(GND_net), .VCC_net(VCC_net), .\next_accum[16] (\next_accum[16] ), 
            .\next_accum[17] (\next_accum[17] ), .\next_accum[18] (\next_accum[18] ), 
            .\next_accum[19] (\next_accum[19] ), .\next_accum[5] (\next_accum[5] ), 
            .\next_accum[4] (\next_accum[4] ), .\cycle[0] (\cycle[0] ), 
            .data_rs1({\data_rs1[3] , data_rs1_c[2:1], data_rs1[0]})) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[31:97])
    tinyqv_shifter i_shift (.tmp_data({tmp_data}), .\alu_op[3] (\alu_op[3] ), 
            .n24268(n24268), .n24864(n24864), .n24865(n24865), .\shift_amt[0] (shift_amt[0]), 
            .n26610(n26610), .\alu_op_in[2] (\alu_op_in[2] ), .\dr_3__N_1595[33] (dr_3__N_1595[33]), 
            .\dr_3__N_1595[32] (dr_3__N_1595[32]), .\shift_amt[1] (shift_amt[1]), 
            .\shift_amt[2] (shift_amt_adj_2358[2]), .\shift_amt[3] (shift_amt_adj_2358[3]), 
            .\counter_hi[2] (counter_hi[2]), .n26608(n26608), .\shift_amt[4] (shift_amt_adj_2358[4]), 
            .\counter_hi[4] (counter_hi[4]), .\shift_out[0] (shift_out[0]), 
            .\shift_out[1] (shift_out[1])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(133[20:81])
    tinyqv_registers i_registers (.rs2({rs2}), .data_rs2({data_rs2}), .rs1({rs1}), 
            .data_rs1({\data_rs1[3] , data_rs1_c[2:1], data_rs1[0]}), 
            .rd({rd}), .debug_reg_wen(debug_reg_wen), .clk_c(clk_c), .return_addr({return_addr}), 
            .debug_rd({debug_rd}), .\reg_access[4][3] (\reg_access[4][3] ), 
            .\reg_access[3][2] (\reg_access[3][2] ), .n26608(n26608), .n26610(n26610), 
            .\counter_hi[2] (counter_hi[2]), .\instr[12] (\instr[12] ), 
            .n25180(n25180), .any_additional_mem_ops(any_additional_mem_ops), 
            .n3645(n3645)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(91[9:103])
    tinyqv_counter_U0 i_instrret (.cy(cy_adj_2), .clk_c(clk_c), .n25424(n25424), 
            .\increment_result_3__N_1656[0] (\increment_result_3__N_1656[0] ), 
            .instrret_count({instrret_count[3:1], \instrret_count[0] }), 
            .n25294(n25294), .n25308(n25308)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(307[20] 315[6])
    \tinyqv_counter(OUTPUT_WIDTH=7)  i_cycles (.cy(cy_adj_3), .clk_c(clk_c), 
            .n25424(n25424), .\increment_result_3__N_1642[1] (\increment_result_3__N_1642[1] ), 
            .\increment_result_3__N_1642[0] (increment_result_3__N_1642[0]), 
            .cycle_count_wide({cycle_count_wide_c[6:4], cycle_count_wide[3], 
            cycle_count_wide_c[2], cycle_count_wide[1:0]}), .n25298(n25298), 
            .n25315(n25315), .n25246(n25246)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(281[40] 290[6])
    tinyqv_alu i_alu (.n22558(n22558), .\alu_op_in[2] (\alu_op_in[2] ), 
            .n25254(n25254), .alu_a_in({alu_a_in[3:2], \alu_a_in[1] , 
            \alu_a_in[0] }), .n25218(n25218), .n25274(n25274), .alu_b_in({alu_b_in_c[3:2], 
            \alu_b_in[1] , alu_b_in[0]}), .n21812(n21812), .n25251(n25251), 
            .cy_out(cy_out), .n24569(n24569), .n25250(n25250), .n25352(n25352), 
            .n25318(n25318), .n25357(n25357), .n24571(n24571), .n4411({n4411}), 
            .n25358(n25358), .alu_out({alu_out})) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(115[16:93])
    
endmodule
//
// Verilog Description of module tinyqv_mul
//

module tinyqv_mul (accum, \next_accum[6] , \next_accum[7] , \next_accum[8] , 
            \next_accum[9] , \next_accum[10] , \next_accum[11] , \next_accum[12] , 
            \next_accum[13] , \next_accum[14] , \next_accum[15] , clk_c, 
            mul_out_3__N_1241, \tmp_data[0] , \tmp_data[1] , \tmp_data[2] , 
            \tmp_data[3] , \tmp_data[4] , \tmp_data[5] , \tmp_data[6] , 
            \tmp_data[7] , \tmp_data[8] , \tmp_data[9] , \tmp_data[10] , 
            \tmp_data[11] , \tmp_data[12] , \tmp_data[13] , \tmp_data[14] , 
            \tmp_data[15] , d_3__N_1599, GND_net, VCC_net, \next_accum[16] , 
            \next_accum[17] , \next_accum[18] , \next_accum[19] , \next_accum[5] , 
            \next_accum[4] , \cycle[0] , data_rs1) /* synthesis syn_module_defined=1 */ ;
    output [15:0]accum;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input clk_c;
    input [3:0]mul_out_3__N_1241;
    input \tmp_data[0] ;
    input \tmp_data[1] ;
    input \tmp_data[2] ;
    input \tmp_data[3] ;
    input \tmp_data[4] ;
    input \tmp_data[5] ;
    input \tmp_data[6] ;
    input \tmp_data[7] ;
    input \tmp_data[8] ;
    input \tmp_data[9] ;
    input \tmp_data[10] ;
    input \tmp_data[11] ;
    input \tmp_data[12] ;
    input \tmp_data[13] ;
    input \tmp_data[14] ;
    input \tmp_data[15] ;
    output [19:0]d_3__N_1599;
    input GND_net;
    input VCC_net;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[5] ;
    input \next_accum[4] ;
    input \cycle[0] ;
    input [3:0]data_rs1;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n7;
    wire [15:0]accum_15__N_1619;
    
    wire n22740;
    
    LUT4 accum_15__I_0_i3_3_lut (.A(accum[6]), .B(\next_accum[6] ), .C(n7), 
         .Z(accum_15__N_1619[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i3_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i4_3_lut (.A(accum[7]), .B(\next_accum[7] ), .C(n7), 
         .Z(accum_15__N_1619[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i4_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i5_3_lut (.A(accum[8]), .B(\next_accum[8] ), .C(n7), 
         .Z(accum_15__N_1619[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i5_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i6_3_lut (.A(accum[9]), .B(\next_accum[9] ), .C(n7), 
         .Z(accum_15__N_1619[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i6_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i7_3_lut (.A(accum[10]), .B(\next_accum[10] ), .C(n7), 
         .Z(accum_15__N_1619[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i7_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i8_3_lut (.A(accum[11]), .B(\next_accum[11] ), .C(n7), 
         .Z(accum_15__N_1619[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i8_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i9_3_lut (.A(accum[12]), .B(\next_accum[12] ), .C(n7), 
         .Z(accum_15__N_1619[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i9_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i10_3_lut (.A(accum[13]), .B(\next_accum[13] ), .C(n7), 
         .Z(accum_15__N_1619[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i10_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i11_3_lut (.A(accum[14]), .B(\next_accum[14] ), .C(n7), 
         .Z(accum_15__N_1619[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i11_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i12_3_lut (.A(accum[15]), .B(\next_accum[15] ), .C(n7), 
         .Z(accum_15__N_1619[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i12_3_lut.init = 16'hacac;
    FD1S3AX accum_i0 (.D(accum_15__N_1619[0]), .CK(clk_c), .Q(accum[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i0.GSR = "DISABLED";
    MULT18X18D a_3__I_0_11_mult_2 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(mul_out_3__N_1241[3]), 
            .A2(mul_out_3__N_1241[2]), .A1(mul_out_3__N_1241[1]), .A0(mul_out_3__N_1241[0]), 
            .B17(GND_net), .B16(GND_net), .B15(\tmp_data[15] ), .B14(\tmp_data[14] ), 
            .B13(\tmp_data[13] ), .B12(\tmp_data[12] ), .B11(\tmp_data[11] ), 
            .B10(\tmp_data[10] ), .B9(\tmp_data[9] ), .B8(\tmp_data[8] ), 
            .B7(\tmp_data[7] ), .B6(\tmp_data[6] ), .B5(\tmp_data[5] ), 
            .B4(\tmp_data[4] ), .B3(\tmp_data[3] ), .B2(\tmp_data[2] ), 
            .B1(\tmp_data[1] ), .B0(\tmp_data[0] ), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .P19(d_3__N_1599[19]), .P18(d_3__N_1599[18]), .P17(d_3__N_1599[17]), 
            .P16(d_3__N_1599[16]), .P15(d_3__N_1599[15]), .P14(d_3__N_1599[14]), 
            .P13(d_3__N_1599[13]), .P12(d_3__N_1599[12]), .P11(d_3__N_1599[11]), 
            .P10(d_3__N_1599[10]), .P9(d_3__N_1599[9]), .P8(d_3__N_1599[8]), 
            .P7(d_3__N_1599[7]), .P6(d_3__N_1599[6]), .P5(d_3__N_1599[5]), 
            .P4(d_3__N_1599[4]), .P3(d_3__N_1599[3]), .P2(d_3__N_1599[2]), 
            .P1(d_3__N_1599[1]), .P0(d_3__N_1599[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[52:83])
    defparam a_3__I_0_11_mult_2.REG_INPUTA_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTA_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTA_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_RST = "RST0";
    defparam a_3__I_0_11_mult_2.CLK0_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK1_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK2_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK3_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.HIGHSPEED_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.GSR = "DISABLED";
    defparam a_3__I_0_11_mult_2.CAS_MATCH_REG = "FALSE";
    defparam a_3__I_0_11_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam a_3__I_0_11_mult_2.MULT_BYPASS = "DISABLED";
    defparam a_3__I_0_11_mult_2.RESETMODE = "SYNC";
    FD1S3IX accum_i12 (.D(\next_accum[16] ), .CK(clk_c), .CD(n7), .Q(accum[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i12.GSR = "DISABLED";
    FD1S3AX accum_i1 (.D(accum_15__N_1619[1]), .CK(clk_c), .Q(accum[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i1.GSR = "DISABLED";
    FD1S3AX accum_i2 (.D(accum_15__N_1619[2]), .CK(clk_c), .Q(accum[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i2.GSR = "DISABLED";
    FD1S3AX accum_i3 (.D(accum_15__N_1619[3]), .CK(clk_c), .Q(accum[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i3.GSR = "DISABLED";
    FD1S3AX accum_i4 (.D(accum_15__N_1619[4]), .CK(clk_c), .Q(accum[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i4.GSR = "DISABLED";
    FD1S3AX accum_i5 (.D(accum_15__N_1619[5]), .CK(clk_c), .Q(accum[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i5.GSR = "DISABLED";
    FD1S3AX accum_i6 (.D(accum_15__N_1619[6]), .CK(clk_c), .Q(accum[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i6.GSR = "DISABLED";
    FD1S3AX accum_i7 (.D(accum_15__N_1619[7]), .CK(clk_c), .Q(accum[7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i7.GSR = "DISABLED";
    FD1S3AX accum_i8 (.D(accum_15__N_1619[8]), .CK(clk_c), .Q(accum[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i8.GSR = "DISABLED";
    FD1S3AX accum_i9 (.D(accum_15__N_1619[9]), .CK(clk_c), .Q(accum[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i9.GSR = "DISABLED";
    FD1S3AX accum_i10 (.D(accum_15__N_1619[10]), .CK(clk_c), .Q(accum[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i10.GSR = "DISABLED";
    FD1S3AX accum_i11 (.D(accum_15__N_1619[11]), .CK(clk_c), .Q(accum[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i11.GSR = "DISABLED";
    FD1S3IX accum_i13 (.D(\next_accum[17] ), .CK(clk_c), .CD(n7), .Q(accum[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i13.GSR = "DISABLED";
    FD1S3IX accum_i14 (.D(\next_accum[18] ), .CK(clk_c), .CD(n7), .Q(accum[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i14.GSR = "DISABLED";
    FD1S3IX accum_i15 (.D(\next_accum[19] ), .CK(clk_c), .CD(n7), .Q(accum[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i15.GSR = "DISABLED";
    LUT4 accum_15__I_0_i2_3_lut (.A(accum[5]), .B(\next_accum[5] ), .C(n7), 
         .Z(accum_15__N_1619[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i2_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i1_3_lut (.A(accum[4]), .B(\next_accum[4] ), .C(n7), 
         .Z(accum_15__N_1619[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i1_3_lut.init = 16'hacac;
    LUT4 i21853_4_lut (.A(\cycle[0] ), .B(n22740), .C(data_rs1[3]), .D(data_rs1[0]), 
         .Z(n7)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:32])
    defparam i21853_4_lut.init = 16'h5557;
    LUT4 i1_2_lut (.A(data_rs1[2]), .B(data_rs1[1]), .Z(n22740)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:32])
    defparam i1_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module tinyqv_shifter
//

module tinyqv_shifter (tmp_data, \alu_op[3] , n24268, n24864, n24865, 
            \shift_amt[0] , n26610, \alu_op_in[2] , \dr_3__N_1595[33] , 
            \dr_3__N_1595[32] , \shift_amt[1] , \shift_amt[2] , \shift_amt[3] , 
            \counter_hi[2] , n26608, \shift_amt[4] , \counter_hi[4] , 
            \shift_out[0] , \shift_out[1] ) /* synthesis syn_module_defined=1 */ ;
    input [31:0]tmp_data;
    input \alu_op[3] ;
    output n24268;
    input n24864;
    output n24865;
    input \shift_amt[0] ;
    input n26610;
    input \alu_op_in[2] ;
    output \dr_3__N_1595[33] ;
    output \dr_3__N_1595[32] ;
    input \shift_amt[1] ;
    input \shift_amt[2] ;
    input \shift_amt[3] ;
    input \counter_hi[2] ;
    input n26608;
    input \shift_amt[4] ;
    input \counter_hi[4] ;
    output \shift_out[0] ;
    output \shift_out[1] ;
    
    wire [5:0]shift_amt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[16:25])
    
    wire n7762, n101, n105, n23892, n23553;
    wire [31:0]a_for_shift_right;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[17:34])
    
    wire n63, n49, n51, n53, n55, n57, n59, n61, n23508, n23509, 
        n23516, n23630;
    wire [65:0]dr_3__N_1595;
    
    wire n23510, n23511, n23517, n7758, n7202, n23512, n23513, 
        n23518, n25433, n129, n125, n121, n117, n47, n113, n43, 
        n45, n109, n58, n60, n23544, n54, n56, n23543, n50, 
        n52, n23542, n46, n48, n23541, n42, n44, n23540, n38, 
        n40, n23539, n34, n36, n23538, n23514, n23515, n23519, 
        n23530, n25395, n4, n23529, n23528, n23523, n23524, n23531, 
        n23527, n23525, n23526, n23532, n23891, n23533, n23890, 
        n41, n37, n39, n33, n35, n23534, n62, n23546, n23547, 
        n23548, n23545, n23549, n23554, n23555, n23556, n23520, 
        n23521, n23535, n23536, n23550, n23551, n23557, n23558, 
        n32;
    
    LUT4 n192_bdd_3_lut_22253_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), 
         .C(shift_amt[5]), .D(n7762), .Z(n24268)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam n192_bdd_3_lut_22253_4_lut.init = 16'h8f80;
    LUT4 n24864_bdd_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n24864), .Z(n24865)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam n24864_bdd_3_lut_4_lut.init = 16'h8f80;
    PFUMX i21278 (.BLUT(n101), .ALUT(n105), .C0(n23892), .Z(n23553));
    LUT4 top_bit_I_0_i63_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), 
         .C(\shift_amt[0] ), .D(a_for_shift_right[31]), .Z(n63)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam top_bit_I_0_i63_3_lut_4_lut.init = 16'h8f80;
    LUT4 top_bit_I_0_i49_3_lut (.A(a_for_shift_right[17]), .B(a_for_shift_right[18]), 
         .C(\shift_amt[0] ), .Z(n49)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i49_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i51_3_lut (.A(a_for_shift_right[19]), .B(a_for_shift_right[20]), 
         .C(\shift_amt[0] ), .Z(n51)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i51_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i53_3_lut (.A(a_for_shift_right[21]), .B(a_for_shift_right[22]), 
         .C(\shift_amt[0] ), .Z(n53)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i53_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i55_3_lut (.A(a_for_shift_right[23]), .B(a_for_shift_right[24]), 
         .C(\shift_amt[0] ), .Z(n55)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i55_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i57_3_lut (.A(a_for_shift_right[25]), .B(a_for_shift_right[26]), 
         .C(\shift_amt[0] ), .Z(n57)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i57_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i59_3_lut (.A(a_for_shift_right[27]), .B(a_for_shift_right[28]), 
         .C(\shift_amt[0] ), .Z(n59)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i59_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i61_3_lut (.A(a_for_shift_right[29]), .B(a_for_shift_right[30]), 
         .C(\shift_amt[0] ), .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i61_3_lut.init = 16'hcaca;
    PFUMX i21241 (.BLUT(n23508), .ALUT(n23509), .C0(shift_amt[2]), .Z(n23516));
    LUT4 i21701_2_lut (.A(n26610), .B(\alu_op_in[2] ), .Z(n23630)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i21701_2_lut.init = 16'h6666;
    LUT4 i5531_3_lut (.A(dr_3__N_1595[31]), .B(dr_3__N_1595[34]), .C(\alu_op_in[2] ), 
         .Z(n7762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i5531_3_lut.init = 16'hcaca;
    PFUMX i21242 (.BLUT(n23510), .ALUT(n23511), .C0(shift_amt[2]), .Z(n23517));
    LUT4 i5527_3_lut (.A(\dr_3__N_1595[33] ), .B(\dr_3__N_1595[32] ), .C(\alu_op_in[2] ), 
         .Z(n7758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i5527_3_lut.init = 16'hcaca;
    LUT4 i4977_3_lut (.A(dr_3__N_1595[34]), .B(dr_3__N_1595[31]), .C(\alu_op_in[2] ), 
         .Z(n7202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i4977_3_lut.init = 16'hcaca;
    PFUMX i21243 (.BLUT(n23512), .ALUT(n23513), .C0(shift_amt[2]), .Z(n23518));
    LUT4 i5017_4_lut (.A(a_for_shift_right[31]), .B(n25433), .C(\shift_amt[0] ), 
         .D(\shift_amt[1] ), .Z(n129)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam i5017_4_lut.init = 16'hccca;
    LUT4 top_bit_I_0_i125_3_lut (.A(n59), .B(n61), .C(\shift_amt[1] ), 
         .Z(n125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i125_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i121_3_lut (.A(n55), .B(n57), .C(\shift_amt[1] ), 
         .Z(n121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i121_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i117_3_lut (.A(n51), .B(n53), .C(\shift_amt[1] ), 
         .Z(n117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i117_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i113_3_lut (.A(n47), .B(n49), .C(\shift_amt[1] ), 
         .Z(n113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i113_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i109_3_lut (.A(n43), .B(n45), .C(\shift_amt[1] ), 
         .Z(n109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i109_3_lut.init = 16'hcaca;
    LUT4 i21269_3_lut (.A(n58), .B(n60), .C(\shift_amt[1] ), .Z(n23544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21269_3_lut.init = 16'hcaca;
    LUT4 i21268_3_lut (.A(n54), .B(n56), .C(\shift_amt[1] ), .Z(n23543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21268_3_lut.init = 16'hcaca;
    LUT4 i21267_3_lut (.A(n50), .B(n52), .C(\shift_amt[1] ), .Z(n23542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21267_3_lut.init = 16'hcaca;
    LUT4 i21266_3_lut (.A(n46), .B(n48), .C(\shift_amt[1] ), .Z(n23541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21266_3_lut.init = 16'hcaca;
    LUT4 i21265_3_lut (.A(n42), .B(n44), .C(\shift_amt[1] ), .Z(n23540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21265_3_lut.init = 16'hcaca;
    LUT4 i21264_3_lut (.A(n38), .B(n40), .C(\shift_amt[1] ), .Z(n23539)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21264_3_lut.init = 16'hcaca;
    LUT4 i21263_3_lut (.A(n34), .B(n36), .C(\shift_amt[1] ), .Z(n23538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21263_3_lut.init = 16'hcaca;
    PFUMX i21244 (.BLUT(n23514), .ALUT(n23515), .C0(shift_amt[2]), .Z(n23519));
    LUT4 i21255_3_lut (.A(n61), .B(n63), .C(\shift_amt[1] ), .Z(n23530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21255_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(\shift_amt[2] ), .B(n25395), .C(n23630), .D(\shift_amt[3] ), 
         .Z(shift_amt[3])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[28:55])
    defparam i2_3_lut_4_lut.init = 16'hd22d;
    LUT4 i3910_3_lut_4_lut (.A(\shift_amt[2] ), .B(n25395), .C(n23630), 
         .D(\shift_amt[3] ), .Z(n4)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[28:55])
    defparam i3910_3_lut_4_lut.init = 16'h2f02;
    LUT4 i21254_3_lut (.A(n57), .B(n59), .C(\shift_amt[1] ), .Z(n23529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21254_3_lut.init = 16'hcaca;
    LUT4 i21253_3_lut (.A(n53), .B(n55), .C(\shift_amt[1] ), .Z(n23528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21253_3_lut.init = 16'hcaca;
    PFUMX i21256 (.BLUT(n23523), .ALUT(n23524), .C0(n23892), .Z(n23531));
    LUT4 i21252_3_lut (.A(n49), .B(n51), .C(\shift_amt[1] ), .Z(n23527)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21252_3_lut.init = 16'hcaca;
    PFUMX i21257 (.BLUT(n23525), .ALUT(n23526), .C0(n23892), .Z(n23532));
    PFUMX i21258 (.BLUT(n23527), .ALUT(n23528), .C0(n23891), .Z(n23533));
    LUT4 i21699_2_lut_rep_659 (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .Z(n25395)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i21699_2_lut_rep_659.init = 16'h6666;
    LUT4 i3897_rep_121_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .C(\shift_amt[2] ), .Z(n23892)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i3897_rep_121_2_lut_3_lut.init = 16'h6969;
    LUT4 i3897_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), .C(\shift_amt[2] ), 
         .Z(shift_amt[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i3897_2_lut_3_lut.init = 16'h6969;
    LUT4 i3897_rep_120_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .C(\shift_amt[2] ), .Z(n23891)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i3897_rep_120_2_lut_3_lut.init = 16'h6969;
    LUT4 i3897_rep_119_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .C(\shift_amt[2] ), .Z(n23890)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i3897_rep_119_2_lut_3_lut.init = 16'h6969;
    LUT4 i21251_3_lut (.A(n45), .B(n47), .C(\shift_amt[1] ), .Z(n23526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21251_3_lut.init = 16'hcaca;
    LUT4 i21250_3_lut (.A(n41), .B(n43), .C(\shift_amt[1] ), .Z(n23525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21250_3_lut.init = 16'hcaca;
    LUT4 i21249_3_lut (.A(n37), .B(n39), .C(\shift_amt[1] ), .Z(n23524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21249_3_lut.init = 16'hcaca;
    LUT4 i21248_3_lut (.A(n33), .B(n35), .C(\shift_amt[1] ), .Z(n23523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21248_3_lut.init = 16'hcaca;
    PFUMX i21259 (.BLUT(n23529), .ALUT(n23530), .C0(n23891), .Z(n23534));
    LUT4 i21240_3_lut (.A(n60), .B(n62), .C(\shift_amt[1] ), .Z(n23515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21240_3_lut.init = 16'hcaca;
    LUT4 i21239_3_lut (.A(n56), .B(n58), .C(\shift_amt[1] ), .Z(n23514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21239_3_lut.init = 16'hcaca;
    LUT4 i21238_3_lut (.A(n52), .B(n54), .C(\shift_amt[1] ), .Z(n23513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21238_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i35_3_lut (.A(a_for_shift_right[3]), .B(a_for_shift_right[4]), 
         .C(\shift_amt[0] ), .Z(n35)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i35_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i37_3_lut (.A(a_for_shift_right[5]), .B(a_for_shift_right[6]), 
         .C(\shift_amt[0] ), .Z(n37)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i37_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i6_3_lut (.A(tmp_data[26]), .B(tmp_data[5]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i7_3_lut (.A(tmp_data[25]), .B(tmp_data[6]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i4_3_lut (.A(tmp_data[28]), .B(tmp_data[3]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i5_3_lut (.A(tmp_data[27]), .B(tmp_data[4]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i39_3_lut (.A(a_for_shift_right[7]), .B(a_for_shift_right[8]), 
         .C(\shift_amt[0] ), .Z(n39)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i39_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i41_3_lut (.A(a_for_shift_right[9]), .B(a_for_shift_right[10]), 
         .C(\shift_amt[0] ), .Z(n41)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i41_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i10_3_lut (.A(tmp_data[22]), .B(tmp_data[9]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i11_3_lut (.A(tmp_data[21]), .B(tmp_data[10]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i8_3_lut (.A(tmp_data[24]), .B(tmp_data[7]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i9_3_lut (.A(tmp_data[23]), .B(tmp_data[8]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 i21237_3_lut (.A(n48), .B(n50), .C(\shift_amt[1] ), .Z(n23512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21237_3_lut.init = 16'hcaca;
    LUT4 i21236_3_lut (.A(n44), .B(n46), .C(\shift_amt[1] ), .Z(n23511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21236_3_lut.init = 16'hcaca;
    LUT4 i21235_3_lut (.A(n40), .B(n42), .C(\shift_amt[1] ), .Z(n23510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21235_3_lut.init = 16'hcaca;
    PFUMX i21271 (.BLUT(n23538), .ALUT(n23539), .C0(n23892), .Z(n23546));
    PFUMX i21272 (.BLUT(n23540), .ALUT(n23541), .C0(n23891), .Z(n23547));
    PFUMX i21273 (.BLUT(n23542), .ALUT(n23543), .C0(n23891), .Z(n23548));
    PFUMX i21274 (.BLUT(n23544), .ALUT(n23545), .C0(n23890), .Z(n23549));
    PFUMX i21279 (.BLUT(n109), .ALUT(n113), .C0(n23890), .Z(n23554));
    PFUMX i21280 (.BLUT(n117), .ALUT(n121), .C0(n23890), .Z(n23555));
    PFUMX i21281 (.BLUT(n125), .ALUT(n129), .C0(n23890), .Z(n23556));
    L6MUX21 i21245 (.D0(n23516), .D1(n23517), .SD(shift_amt[3]), .Z(n23520));
    LUT4 i3917_3_lut_4_lut (.A(n26608), .B(\alu_op_in[2] ), .C(n4), .D(\shift_amt[4] ), 
         .Z(shift_amt[5])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i3917_3_lut_4_lut.init = 16'hf990;
    LUT4 i2_3_lut_4_lut_adj_205 (.A(\counter_hi[4] ), .B(\alu_op_in[2] ), 
         .C(n4), .D(\shift_amt[4] ), .Z(shift_amt[4])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i2_3_lut_4_lut_adj_205.init = 16'h9669;
    L6MUX21 i21246 (.D0(n23518), .D1(n23519), .SD(shift_amt[3]), .Z(n23521));
    L6MUX21 i21260 (.D0(n23531), .D1(n23532), .SD(shift_amt[3]), .Z(n23535));
    L6MUX21 i21261 (.D0(n23533), .D1(n23534), .SD(shift_amt[3]), .Z(n23536));
    L6MUX21 i21275 (.D0(n23546), .D1(n23547), .SD(shift_amt[3]), .Z(n23550));
    L6MUX21 i21276 (.D0(n23548), .D1(n23549), .SD(shift_amt[3]), .Z(n23551));
    LUT4 i21234_3_lut (.A(n36), .B(n38), .C(\shift_amt[1] ), .Z(n23509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21234_3_lut.init = 16'hcaca;
    L6MUX21 i21282 (.D0(n23553), .D1(n23554), .SD(shift_amt[3]), .Z(n23557));
    L6MUX21 i21283 (.D0(n23555), .D1(n23556), .SD(shift_amt[3]), .Z(n23558));
    LUT4 i21233_3_lut (.A(n32), .B(n34), .C(\shift_amt[1] ), .Z(n23508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21233_3_lut.init = 16'hcaca;
    LUT4 i11736_2_lut_rep_697 (.A(tmp_data[31]), .B(\alu_op[3] ), .Z(n25433)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i11736_2_lut_rep_697.init = 16'h8888;
    LUT4 i21270_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(\shift_amt[1] ), 
         .D(n62), .Z(n23545)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i21270_3_lut_4_lut.init = 16'h8f80;
    LUT4 i4978_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n7202), .Z(\shift_out[0] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i4978_3_lut_4_lut.init = 16'h8f80;
    LUT4 i5528_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n7758), .Z(\shift_out[1] )) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i5528_3_lut_4_lut.init = 16'h8f80;
    LUT4 top_bit_I_0_i48_3_lut (.A(a_for_shift_right[16]), .B(a_for_shift_right[17]), 
         .C(\shift_amt[0] ), .Z(n48)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i48_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i17_3_lut (.A(tmp_data[15]), .B(tmp_data[16]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i50_3_lut (.A(a_for_shift_right[18]), .B(a_for_shift_right[19]), 
         .C(\shift_amt[0] ), .Z(n50)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i50_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i19_3_lut (.A(tmp_data[13]), .B(tmp_data[18]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i20_3_lut (.A(tmp_data[12]), .B(tmp_data[19]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i18_3_lut (.A(tmp_data[14]), .B(tmp_data[17]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i52_3_lut (.A(a_for_shift_right[20]), .B(a_for_shift_right[21]), 
         .C(\shift_amt[0] ), .Z(n52)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i52_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i54_3_lut (.A(a_for_shift_right[22]), .B(a_for_shift_right[23]), 
         .C(\shift_amt[0] ), .Z(n54)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i54_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i23_3_lut (.A(tmp_data[9]), .B(tmp_data[22]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i24_3_lut (.A(tmp_data[8]), .B(tmp_data[23]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i21_3_lut (.A(tmp_data[11]), .B(tmp_data[20]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i22_3_lut (.A(tmp_data[10]), .B(tmp_data[21]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i56_3_lut (.A(a_for_shift_right[24]), .B(a_for_shift_right[25]), 
         .C(\shift_amt[0] ), .Z(n56)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i56_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i58_3_lut (.A(a_for_shift_right[26]), .B(a_for_shift_right[27]), 
         .C(\shift_amt[0] ), .Z(n58)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i58_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i27_3_lut (.A(tmp_data[5]), .B(tmp_data[26]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i28_3_lut (.A(tmp_data[4]), .B(tmp_data[27]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i25_3_lut (.A(tmp_data[7]), .B(tmp_data[24]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i26_3_lut (.A(tmp_data[6]), .B(tmp_data[25]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i60_3_lut (.A(a_for_shift_right[28]), .B(a_for_shift_right[29]), 
         .C(\shift_amt[0] ), .Z(n60)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i60_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i62_3_lut (.A(a_for_shift_right[30]), .B(a_for_shift_right[31]), 
         .C(\shift_amt[0] ), .Z(n62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i62_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i31_3_lut (.A(tmp_data[1]), .B(tmp_data[30]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i32_3_lut (.A(tmp_data[0]), .B(tmp_data[31]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i29_3_lut (.A(tmp_data[3]), .B(tmp_data[28]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i30_3_lut (.A(tmp_data[2]), .B(tmp_data[29]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i105_3_lut (.A(n39), .B(n41), .C(\shift_amt[1] ), 
         .Z(n105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i105_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i32_3_lut (.A(a_for_shift_right[0]), .B(a_for_shift_right[1]), 
         .C(\shift_amt[0] ), .Z(n32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i32_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i101_3_lut (.A(n35), .B(n37), .C(\shift_amt[1] ), 
         .Z(n101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i101_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i1_3_lut (.A(tmp_data[31]), .B(tmp_data[0]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i34_3_lut (.A(a_for_shift_right[2]), .B(a_for_shift_right[3]), 
         .C(\shift_amt[0] ), .Z(n34)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i34_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i3_3_lut (.A(tmp_data[29]), .B(tmp_data[2]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i2_3_lut (.A(tmp_data[30]), .B(tmp_data[1]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i36_3_lut (.A(a_for_shift_right[4]), .B(a_for_shift_right[5]), 
         .C(\shift_amt[0] ), .Z(n36)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i36_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i38_3_lut (.A(a_for_shift_right[6]), .B(a_for_shift_right[7]), 
         .C(\shift_amt[0] ), .Z(n38)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i38_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i33_3_lut (.A(a_for_shift_right[1]), .B(a_for_shift_right[2]), 
         .C(\shift_amt[0] ), .Z(n33)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i33_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i43_3_lut (.A(a_for_shift_right[11]), .B(a_for_shift_right[12]), 
         .C(\shift_amt[0] ), .Z(n43)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i43_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i45_3_lut (.A(a_for_shift_right[13]), .B(a_for_shift_right[14]), 
         .C(\shift_amt[0] ), .Z(n45)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i45_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i47_4_lut (.A(tmp_data[16]), .B(tmp_data[15]), .C(\alu_op_in[2] ), 
         .D(\shift_amt[0] ), .Z(n47)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A !((C (D)+!C !(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i47_4_lut.init = 16'hacca;
    L6MUX21 i21247 (.D0(n23520), .D1(n23521), .SD(shift_amt[4]), .Z(dr_3__N_1595[31]));
    L6MUX21 i21262 (.D0(n23535), .D1(n23536), .SD(shift_amt[4]), .Z(\dr_3__N_1595[32] ));
    L6MUX21 i21277 (.D0(n23550), .D1(n23551), .SD(shift_amt[4]), .Z(\dr_3__N_1595[33] ));
    L6MUX21 i21284 (.D0(n23557), .D1(n23558), .SD(shift_amt[4]), .Z(dr_3__N_1595[34]));
    LUT4 top_bit_I_0_i40_3_lut (.A(a_for_shift_right[8]), .B(a_for_shift_right[9]), 
         .C(\shift_amt[0] ), .Z(n40)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i40_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i42_3_lut (.A(a_for_shift_right[10]), .B(a_for_shift_right[11]), 
         .C(\shift_amt[0] ), .Z(n42)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i42_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i12_3_lut (.A(tmp_data[20]), .B(tmp_data[11]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i44_3_lut (.A(a_for_shift_right[12]), .B(a_for_shift_right[13]), 
         .C(\shift_amt[0] ), .Z(n44)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i44_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i46_3_lut (.A(a_for_shift_right[14]), .B(a_for_shift_right[15]), 
         .C(\shift_amt[0] ), .Z(n46)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i46_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i16_3_lut (.A(tmp_data[16]), .B(tmp_data[15]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i16_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i13_3_lut (.A(tmp_data[19]), .B(tmp_data[12]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i14_3_lut (.A(tmp_data[18]), .B(tmp_data[13]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i15_3_lut (.A(tmp_data[17]), .B(tmp_data[14]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i15_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module tinyqv_registers
//

module tinyqv_registers (rs2, data_rs2, rs1, data_rs1, rd, debug_reg_wen, 
            clk_c, return_addr, debug_rd, \reg_access[4][3] , \reg_access[3][2] , 
            n26608, n26610, \counter_hi[2] , \instr[12] , n25180, 
            any_additional_mem_ops, n3645) /* synthesis syn_module_defined=1 */ ;
    input [3:0]rs2;
    output [3:0]data_rs2;
    input [3:0]rs1;
    output [3:0]data_rs1;
    input [3:0]rd;
    input debug_reg_wen;
    input clk_c;
    output [23:1]return_addr;
    input [3:0]debug_rd;
    output \reg_access[4][3] ;
    output \reg_access[3][2] ;
    input n26608;
    input n26610;
    input \counter_hi[2] ;
    input \instr[12] ;
    input n25180;
    input any_additional_mem_ops;
    output n3645;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n23460, n23461, n23475, n23476, n23490, n23491, n23505, 
        n23506, n23448, n23449, n23456, n25186, n25185, n25184;
    wire [31:0]\registers[14] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[15] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n12;
    wire [31:0]\registers[12] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[13] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n11, n25183;
    wire [31:0]\registers[10] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[11] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n9;
    wire [31:0]\registers[8] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[9] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n8, n12_adj_2331, n11_adj_2332, n9_adj_2333, n8_adj_2334, 
        n23500, n23499, n23463, n23464, n23471, n23498, n23497;
    wire [31:0]\registers[6] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[7] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n23496;
    wire [31:0]\registers[5] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n23495, n23478, n23479, n23486, n23485, n23484, n23483, 
        n23482, n23481, n23493, n23494, n23501, n23480, n23470, 
        n23469;
    wire [31:0]\registers[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_1__2__N_1487, n23468, registers_1__1__N_1488, registers_1__0__N_1489;
    wire [31:0]\registers[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_2__3__N_1490, registers_2__2__N_1493, registers_2__1__N_1494, 
        registers_2__0__N_1495, registers_5__3__N_1496, registers_5__2__N_1499, 
        registers_5__1__N_1500, registers_5__0__N_1501, registers_6__3__N_1502, 
        registers_6__2__N_1505, registers_6__1__N_1506, registers_6__0__N_1507, 
        registers_7__3__N_1508, registers_7__2__N_1511, n23467, registers_7__1__N_1512, 
        registers_7__0__N_1513, registers_8__3__N_1514, registers_8__2__N_1517, 
        registers_8__1__N_1518, registers_8__0__N_1519, registers_9__3__N_1520, 
        registers_9__2__N_1523, registers_9__1__N_1524, registers_9__0__N_1525, 
        registers_10__3__N_1526, registers_10__2__N_1529, registers_10__1__N_1530, 
        registers_10__0__N_1531, registers_11__3__N_1532, registers_11__2__N_1535, 
        registers_11__1__N_1536, registers_11__0__N_1537, registers_12__3__N_1538, 
        registers_12__2__N_1541, registers_12__1__N_1542, registers_12__0__N_1543, 
        registers_13__3__N_1544, registers_13__2__N_1547, registers_13__1__N_1548, 
        registers_13__0__N_1549, registers_14__3__N_1550, registers_14__2__N_1553, 
        registers_14__1__N_1554, registers_14__0__N_1555, registers_15__3__N_1556, 
        registers_15__2__N_1559, registers_15__1__N_1560, registers_15__0__N_1561, 
        registers_1__3__N_1484, n23466, n23465, n23455, n23454, n23453, 
        n23452, n23451, n23450, n25377, n23417, n23418, n12_adj_2335, 
        n25379, n11_adj_2336, n9_adj_2337, n8_adj_2338, n5, n12_adj_2339, 
        n11_adj_2340, n9_adj_2341, n8_adj_2342, n5_adj_2343, n25380, 
        n5_adj_2344, n4, n23568, n5_adj_2345, n4_adj_2346, n23561, 
        n25382, n23457, n23410, n23411, n23567, n23472, n23487, 
        n23502, n23407, n23560, n23413, n23406, n23414, n23408, 
        n23409, n23415, n23416, n23571, n23572, n23564, n23458, 
        n23459, n23473, n23474, n23488, n23489, n23503, n23504, 
        n23562, n23563, n23565, n23569, n23570;
    
    L6MUX21 i21187 (.D0(n23460), .D1(n23461), .SD(rs2[3]), .Z(data_rs2[0]));
    L6MUX21 i21202 (.D0(n23475), .D1(n23476), .SD(rs1[3]), .Z(data_rs1[0]));
    L6MUX21 i21217 (.D0(n23490), .D1(n23491), .SD(rs1[3]), .Z(data_rs1[2]));
    L6MUX21 i21232 (.D0(n23505), .D1(n23506), .SD(rs2[3]), .Z(data_rs2[2]));
    PFUMX i21181 (.BLUT(n23448), .ALUT(n23449), .C0(rs2[1]), .Z(n23456));
    LUT4 i1_2_lut_rep_450_3_lut (.A(rd[1]), .B(rd[0]), .C(debug_reg_wen), 
         .Z(n25186)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_rep_450_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_449_3_lut (.A(rd[1]), .B(debug_reg_wen), .C(rd[0]), 
         .Z(n25185)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_449_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_448_3_lut (.A(rd[1]), .B(rd[0]), .C(debug_reg_wen), 
         .Z(n25184)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_448_3_lut.init = 16'h8080;
    LUT4 rs2_3__I_0_Mux_3_i12_3_lut (.A(\registers[14] [7]), .B(\registers[15] [7]), 
         .C(rs2[0]), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i12_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i11_3_lut (.A(\registers[12] [7]), .B(\registers[13] [7]), 
         .C(rs2[0]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_447_3_lut (.A(rd[1]), .B(debug_reg_wen), .C(rd[0]), 
         .Z(n25183)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_rep_447_3_lut.init = 16'h0404;
    LUT4 rs2_3__I_0_Mux_3_i9_3_lut (.A(\registers[10] [7]), .B(\registers[11] [7]), 
         .C(rs2[0]), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i8_3_lut (.A(\registers[8] [7]), .B(\registers[9] [7]), 
         .C(rs2[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i12_3_lut (.A(\registers[14] [7]), .B(\registers[15] [7]), 
         .C(rs1[0]), .Z(n12_adj_2331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i12_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i11_3_lut (.A(\registers[12] [7]), .B(\registers[13] [7]), 
         .C(rs1[0]), .Z(n11_adj_2332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i9_3_lut (.A(\registers[10] [7]), .B(\registers[11] [7]), 
         .C(rs1[0]), .Z(n9_adj_2333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i8_3_lut (.A(\registers[8] [7]), .B(\registers[9] [7]), 
         .C(rs1[0]), .Z(n8_adj_2334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 i21225_3_lut (.A(\registers[14] [6]), .B(\registers[15] [6]), .C(rs2[0]), 
         .Z(n23500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21225_3_lut.init = 16'hcaca;
    LUT4 i21224_3_lut (.A(\registers[12] [6]), .B(\registers[13] [6]), .C(rs2[0]), 
         .Z(n23499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21224_3_lut.init = 16'hcaca;
    PFUMX i21196 (.BLUT(n23463), .ALUT(n23464), .C0(rs1[1]), .Z(n23471));
    LUT4 i21223_3_lut (.A(\registers[10] [6]), .B(\registers[11] [6]), .C(rs2[0]), 
         .Z(n23498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21223_3_lut.init = 16'hcaca;
    LUT4 i21222_3_lut (.A(\registers[8] [6]), .B(\registers[9] [6]), .C(rs2[0]), 
         .Z(n23497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21222_3_lut.init = 16'hcaca;
    LUT4 i21221_3_lut (.A(\registers[6] [6]), .B(\registers[7] [6]), .C(rs2[0]), 
         .Z(n23496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21221_3_lut.init = 16'hcaca;
    LUT4 i21220_3_lut (.A(\registers[5] [6]), .B(rs2[0]), .Z(n23495)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21220_3_lut.init = 16'h8888;
    PFUMX i21211 (.BLUT(n23478), .ALUT(n23479), .C0(rs1[1]), .Z(n23486));
    LUT4 i21210_3_lut (.A(\registers[14] [6]), .B(\registers[15] [6]), .C(rs1[0]), 
         .Z(n23485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21210_3_lut.init = 16'hcaca;
    LUT4 i21209_3_lut (.A(\registers[12] [6]), .B(\registers[13] [6]), .C(rs1[0]), 
         .Z(n23484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21209_3_lut.init = 16'hcaca;
    LUT4 i21208_3_lut (.A(\registers[10] [6]), .B(\registers[11] [6]), .C(rs1[0]), 
         .Z(n23483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21208_3_lut.init = 16'hcaca;
    LUT4 i21207_3_lut (.A(\registers[8] [6]), .B(\registers[9] [6]), .C(rs1[0]), 
         .Z(n23482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21207_3_lut.init = 16'hcaca;
    LUT4 i21206_3_lut (.A(\registers[6] [6]), .B(\registers[7] [6]), .C(rs1[0]), 
         .Z(n23481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21206_3_lut.init = 16'hcaca;
    PFUMX i21226 (.BLUT(n23493), .ALUT(n23494), .C0(rs2[1]), .Z(n23501));
    LUT4 i21205_3_lut (.A(\registers[5] [6]), .B(rs1[0]), .Z(n23480)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21205_3_lut.init = 16'h8888;
    LUT4 i21195_3_lut (.A(\registers[14] [4]), .B(\registers[15] [4]), .C(rs1[0]), 
         .Z(n23470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21195_3_lut.init = 16'hcaca;
    LUT4 i21194_3_lut (.A(\registers[12] [4]), .B(\registers[13] [4]), .C(rs1[0]), 
         .Z(n23469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21194_3_lut.init = 16'hcaca;
    FD1S3AX \registers_1[[2__504  (.D(registers_1__2__N_1487), .CK(clk_c), 
            .Q(\registers[1] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[2__504 .GSR = "DISABLED";
    LUT4 i21193_3_lut (.A(\registers[10] [4]), .B(\registers[11] [4]), .C(rs1[0]), 
         .Z(n23468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21193_3_lut.init = 16'hcaca;
    FD1S3AX \registers_1[[1__505  (.D(registers_1__1__N_1488), .CK(clk_c), 
            .Q(\registers[1] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[1__505 .GSR = "DISABLED";
    FD1S3AX \registers_1[[0__506  (.D(registers_1__0__N_1489), .CK(clk_c), 
            .Q(\registers[1] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[0__506 .GSR = "DISABLED";
    FD1S3AX \registers_1[[31__507  (.D(\registers[1] [3]), .CK(clk_c), .Q(return_addr[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[31__507 .GSR = "DISABLED";
    FD1S3AX \registers_1[[30__508  (.D(\registers[1] [2]), .CK(clk_c), .Q(return_addr[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[30__508 .GSR = "DISABLED";
    FD1S3AX \registers_1[[29__509  (.D(\registers[1] [1]), .CK(clk_c), .Q(return_addr[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[29__509 .GSR = "DISABLED";
    FD1S3AX \registers_1[[28__510  (.D(\registers[1] [0]), .CK(clk_c), .Q(return_addr[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[28__510 .GSR = "DISABLED";
    FD1S3AX \registers_1[[27__511  (.D(return_addr[23]), .CK(clk_c), .Q(return_addr[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[27__511 .GSR = "DISABLED";
    FD1S3AX \registers_1[[26__512  (.D(return_addr[22]), .CK(clk_c), .Q(return_addr[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[26__512 .GSR = "DISABLED";
    FD1S3AX \registers_1[[25__513  (.D(return_addr[21]), .CK(clk_c), .Q(return_addr[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[25__513 .GSR = "DISABLED";
    FD1S3AX \registers_1[[24__514  (.D(return_addr[20]), .CK(clk_c), .Q(return_addr[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[24__514 .GSR = "DISABLED";
    FD1S3AX \registers_1[[23__515  (.D(return_addr[19]), .CK(clk_c), .Q(return_addr[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[23__515 .GSR = "DISABLED";
    FD1S3AX \registers_1[[22__516  (.D(return_addr[18]), .CK(clk_c), .Q(return_addr[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[22__516 .GSR = "DISABLED";
    FD1S3AX \registers_1[[21__517  (.D(return_addr[17]), .CK(clk_c), .Q(return_addr[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[21__517 .GSR = "DISABLED";
    FD1S3AX \registers_1[[20__518  (.D(return_addr[16]), .CK(clk_c), .Q(return_addr[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[20__518 .GSR = "DISABLED";
    FD1S3AX \registers_1[[19__519  (.D(return_addr[15]), .CK(clk_c), .Q(return_addr[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[19__519 .GSR = "DISABLED";
    FD1S3AX \registers_1[[18__520  (.D(return_addr[14]), .CK(clk_c), .Q(return_addr[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[18__520 .GSR = "DISABLED";
    FD1S3AX \registers_1[[17__521  (.D(return_addr[13]), .CK(clk_c), .Q(return_addr[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[17__521 .GSR = "DISABLED";
    FD1S3AX \registers_1[[16__522  (.D(return_addr[12]), .CK(clk_c), .Q(return_addr[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[16__522 .GSR = "DISABLED";
    FD1S3AX \registers_1[[15__523  (.D(return_addr[11]), .CK(clk_c), .Q(return_addr[7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[15__523 .GSR = "DISABLED";
    FD1S3AX \registers_1[[14__524  (.D(return_addr[10]), .CK(clk_c), .Q(return_addr[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[14__524 .GSR = "DISABLED";
    FD1S3AX \registers_1[[13__525  (.D(return_addr[9]), .CK(clk_c), .Q(return_addr[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[13__525 .GSR = "DISABLED";
    FD1S3AX \registers_1[[12__526  (.D(return_addr[8]), .CK(clk_c), .Q(return_addr[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[12__526 .GSR = "DISABLED";
    FD1S3AX \registers_1[[11__527  (.D(return_addr[7]), .CK(clk_c), .Q(return_addr[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[11__527 .GSR = "DISABLED";
    FD1S3AX \registers_1[[10__528  (.D(return_addr[6]), .CK(clk_c), .Q(return_addr[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[10__528 .GSR = "DISABLED";
    FD1S3AX \registers_1[[9__529  (.D(return_addr[5]), .CK(clk_c), .Q(return_addr[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[9__529 .GSR = "DISABLED";
    FD1S3AX \registers_1[[8__530  (.D(return_addr[4]), .CK(clk_c), .Q(\registers[1] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[8__530 .GSR = "DISABLED";
    FD1S3AX \registers_1[[7__531  (.D(return_addr[3]), .CK(clk_c), .Q(\registers[1] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[7__531 .GSR = "DISABLED";
    FD1S3AX \registers_1[[6__532  (.D(return_addr[2]), .CK(clk_c), .Q(\registers[1] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[6__532 .GSR = "DISABLED";
    FD1S3AX \registers_1[[5__533  (.D(return_addr[1]), .CK(clk_c), .Q(\registers[1] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[5__533 .GSR = "DISABLED";
    FD1S3AX \registers_1[[4__534  (.D(\registers[1] [8]), .CK(clk_c), .Q(\registers[1] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[4__534 .GSR = "DISABLED";
    FD1S3AX \registers_2[[3__535  (.D(registers_2__3__N_1490), .CK(clk_c), 
            .Q(\registers[2] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[3__535 .GSR = "DISABLED";
    FD1S3AX \registers_2[[2__536  (.D(registers_2__2__N_1493), .CK(clk_c), 
            .Q(\registers[2] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[2__536 .GSR = "DISABLED";
    FD1S3AX \registers_2[[1__537  (.D(registers_2__1__N_1494), .CK(clk_c), 
            .Q(\registers[2] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[1__537 .GSR = "DISABLED";
    FD1S3AX \registers_2[[0__538  (.D(registers_2__0__N_1495), .CK(clk_c), 
            .Q(\registers[2] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[0__538 .GSR = "DISABLED";
    FD1S3AX \registers_2[[31__539  (.D(\registers[2] [3]), .CK(clk_c), .Q(\registers[2] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[31__539 .GSR = "DISABLED";
    FD1S3AX \registers_2[[30__540  (.D(\registers[2] [2]), .CK(clk_c), .Q(\registers[2] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[30__540 .GSR = "DISABLED";
    FD1S3AX \registers_2[[29__541  (.D(\registers[2] [1]), .CK(clk_c), .Q(\registers[2] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[29__541 .GSR = "DISABLED";
    FD1S3AX \registers_2[[28__542  (.D(\registers[2] [0]), .CK(clk_c), .Q(\registers[2] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[28__542 .GSR = "DISABLED";
    FD1S3AX \registers_2[[27__543  (.D(\registers[2] [31]), .CK(clk_c), 
            .Q(\registers[2] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[27__543 .GSR = "DISABLED";
    FD1S3AX \registers_2[[26__544  (.D(\registers[2] [30]), .CK(clk_c), 
            .Q(\registers[2] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[26__544 .GSR = "DISABLED";
    FD1S3AX \registers_2[[25__545  (.D(\registers[2] [29]), .CK(clk_c), 
            .Q(\registers[2] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[25__545 .GSR = "DISABLED";
    FD1S3AX \registers_2[[24__546  (.D(\registers[2] [28]), .CK(clk_c), 
            .Q(\registers[2] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[24__546 .GSR = "DISABLED";
    FD1S3AX \registers_2[[23__547  (.D(\registers[2] [27]), .CK(clk_c), 
            .Q(\registers[2] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[23__547 .GSR = "DISABLED";
    FD1S3AX \registers_2[[22__548  (.D(\registers[2] [26]), .CK(clk_c), 
            .Q(\registers[2] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[22__548 .GSR = "DISABLED";
    FD1S3AX \registers_2[[21__549  (.D(\registers[2] [25]), .CK(clk_c), 
            .Q(\registers[2] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[21__549 .GSR = "DISABLED";
    FD1S3AX \registers_2[[20__550  (.D(\registers[2] [24]), .CK(clk_c), 
            .Q(\registers[2] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[20__550 .GSR = "DISABLED";
    FD1S3AX \registers_2[[19__551  (.D(\registers[2] [23]), .CK(clk_c), 
            .Q(\registers[2] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[19__551 .GSR = "DISABLED";
    FD1S3AX \registers_2[[18__552  (.D(\registers[2] [22]), .CK(clk_c), 
            .Q(\registers[2] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[18__552 .GSR = "DISABLED";
    FD1S3AX \registers_2[[17__553  (.D(\registers[2] [21]), .CK(clk_c), 
            .Q(\registers[2] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[17__553 .GSR = "DISABLED";
    FD1S3AX \registers_2[[16__554  (.D(\registers[2] [20]), .CK(clk_c), 
            .Q(\registers[2] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[16__554 .GSR = "DISABLED";
    FD1S3AX \registers_2[[15__555  (.D(\registers[2] [19]), .CK(clk_c), 
            .Q(\registers[2] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[15__555 .GSR = "DISABLED";
    FD1S3AX \registers_2[[14__556  (.D(\registers[2] [18]), .CK(clk_c), 
            .Q(\registers[2] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[14__556 .GSR = "DISABLED";
    FD1S3AX \registers_2[[13__557  (.D(\registers[2] [17]), .CK(clk_c), 
            .Q(\registers[2] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[13__557 .GSR = "DISABLED";
    FD1S3AX \registers_2[[12__558  (.D(\registers[2] [16]), .CK(clk_c), 
            .Q(\registers[2] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[12__558 .GSR = "DISABLED";
    FD1S3AX \registers_2[[11__559  (.D(\registers[2] [15]), .CK(clk_c), 
            .Q(\registers[2] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[11__559 .GSR = "DISABLED";
    FD1S3AX \registers_2[[10__560  (.D(\registers[2] [14]), .CK(clk_c), 
            .Q(\registers[2] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[10__560 .GSR = "DISABLED";
    FD1S3AX \registers_2[[9__561  (.D(\registers[2] [13]), .CK(clk_c), .Q(\registers[2] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[9__561 .GSR = "DISABLED";
    FD1S3AX \registers_2[[8__562  (.D(\registers[2] [12]), .CK(clk_c), .Q(\registers[2] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[8__562 .GSR = "DISABLED";
    FD1S3AX \registers_2[[7__563  (.D(\registers[2] [11]), .CK(clk_c), .Q(\registers[2] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[7__563 .GSR = "DISABLED";
    FD1S3AX \registers_2[[6__564  (.D(\registers[2] [10]), .CK(clk_c), .Q(\registers[2] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[6__564 .GSR = "DISABLED";
    FD1S3AX \registers_2[[5__565  (.D(\registers[2] [9]), .CK(clk_c), .Q(\registers[2] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[5__565 .GSR = "DISABLED";
    FD1S3AX \registers_2[[4__566  (.D(\registers[2] [8]), .CK(clk_c), .Q(\registers[2] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[4__566 .GSR = "DISABLED";
    FD1S3AX \registers_5[[3__567  (.D(registers_5__3__N_1496), .CK(clk_c), 
            .Q(\registers[5] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[3__567 .GSR = "DISABLED";
    FD1S3AX \registers_5[[2__568  (.D(registers_5__2__N_1499), .CK(clk_c), 
            .Q(\registers[5] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[2__568 .GSR = "DISABLED";
    FD1S3AX \registers_5[[1__569  (.D(registers_5__1__N_1500), .CK(clk_c), 
            .Q(\registers[5] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[1__569 .GSR = "DISABLED";
    FD1S3AX \registers_5[[0__570  (.D(registers_5__0__N_1501), .CK(clk_c), 
            .Q(\registers[5] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[0__570 .GSR = "DISABLED";
    FD1S3AX \registers_5[[31__571  (.D(\registers[5] [3]), .CK(clk_c), .Q(\registers[5] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[31__571 .GSR = "DISABLED";
    FD1S3AX \registers_5[[30__572  (.D(\registers[5] [2]), .CK(clk_c), .Q(\registers[5] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[30__572 .GSR = "DISABLED";
    FD1S3AX \registers_5[[29__573  (.D(\registers[5] [1]), .CK(clk_c), .Q(\registers[5] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[29__573 .GSR = "DISABLED";
    FD1S3AX \registers_5[[28__574  (.D(\registers[5] [0]), .CK(clk_c), .Q(\registers[5] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[28__574 .GSR = "DISABLED";
    FD1S3AX \registers_5[[27__575  (.D(\registers[5] [31]), .CK(clk_c), 
            .Q(\registers[5] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[27__575 .GSR = "DISABLED";
    FD1S3AX \registers_5[[26__576  (.D(\registers[5] [30]), .CK(clk_c), 
            .Q(\registers[5] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[26__576 .GSR = "DISABLED";
    FD1S3AX \registers_5[[25__577  (.D(\registers[5] [29]), .CK(clk_c), 
            .Q(\registers[5] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[25__577 .GSR = "DISABLED";
    FD1S3AX \registers_5[[24__578  (.D(\registers[5] [28]), .CK(clk_c), 
            .Q(\registers[5] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[24__578 .GSR = "DISABLED";
    FD1S3AX \registers_5[[23__579  (.D(\registers[5] [27]), .CK(clk_c), 
            .Q(\registers[5] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[23__579 .GSR = "DISABLED";
    FD1S3AX \registers_5[[22__580  (.D(\registers[5] [26]), .CK(clk_c), 
            .Q(\registers[5] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[22__580 .GSR = "DISABLED";
    FD1S3AX \registers_5[[21__581  (.D(\registers[5] [25]), .CK(clk_c), 
            .Q(\registers[5] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[21__581 .GSR = "DISABLED";
    FD1S3AX \registers_5[[20__582  (.D(\registers[5] [24]), .CK(clk_c), 
            .Q(\registers[5] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[20__582 .GSR = "DISABLED";
    FD1S3AX \registers_5[[19__583  (.D(\registers[5] [23]), .CK(clk_c), 
            .Q(\registers[5] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[19__583 .GSR = "DISABLED";
    FD1S3AX \registers_5[[18__584  (.D(\registers[5] [22]), .CK(clk_c), 
            .Q(\registers[5] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[18__584 .GSR = "DISABLED";
    FD1S3AX \registers_5[[17__585  (.D(\registers[5] [21]), .CK(clk_c), 
            .Q(\registers[5] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[17__585 .GSR = "DISABLED";
    FD1S3AX \registers_5[[16__586  (.D(\registers[5] [20]), .CK(clk_c), 
            .Q(\registers[5] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[16__586 .GSR = "DISABLED";
    FD1S3AX \registers_5[[15__587  (.D(\registers[5] [19]), .CK(clk_c), 
            .Q(\registers[5] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[15__587 .GSR = "DISABLED";
    FD1S3AX \registers_5[[14__588  (.D(\registers[5] [18]), .CK(clk_c), 
            .Q(\registers[5] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[14__588 .GSR = "DISABLED";
    FD1S3AX \registers_5[[13__589  (.D(\registers[5] [17]), .CK(clk_c), 
            .Q(\registers[5] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[13__589 .GSR = "DISABLED";
    FD1S3AX \registers_5[[12__590  (.D(\registers[5] [16]), .CK(clk_c), 
            .Q(\registers[5] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[12__590 .GSR = "DISABLED";
    FD1S3AX \registers_5[[11__591  (.D(\registers[5] [15]), .CK(clk_c), 
            .Q(\registers[5] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[11__591 .GSR = "DISABLED";
    FD1S3AX \registers_5[[10__592  (.D(\registers[5] [14]), .CK(clk_c), 
            .Q(\registers[5] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[10__592 .GSR = "DISABLED";
    FD1S3AX \registers_5[[9__593  (.D(\registers[5] [13]), .CK(clk_c), .Q(\registers[5] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[9__593 .GSR = "DISABLED";
    FD1S3AX \registers_5[[8__594  (.D(\registers[5] [12]), .CK(clk_c), .Q(\registers[5] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[8__594 .GSR = "DISABLED";
    FD1S3AX \registers_5[[7__595  (.D(\registers[5] [11]), .CK(clk_c), .Q(\registers[5] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[7__595 .GSR = "DISABLED";
    FD1S3AX \registers_5[[6__596  (.D(\registers[5] [10]), .CK(clk_c), .Q(\registers[5] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[6__596 .GSR = "DISABLED";
    FD1S3AX \registers_5[[5__597  (.D(\registers[5] [9]), .CK(clk_c), .Q(\registers[5] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[5__597 .GSR = "DISABLED";
    FD1S3AX \registers_5[[4__598  (.D(\registers[5] [8]), .CK(clk_c), .Q(\registers[5] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[4__598 .GSR = "DISABLED";
    FD1S3AX \registers_6[[3__599  (.D(registers_6__3__N_1502), .CK(clk_c), 
            .Q(\registers[6] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[3__599 .GSR = "DISABLED";
    FD1S3AX \registers_6[[2__600  (.D(registers_6__2__N_1505), .CK(clk_c), 
            .Q(\registers[6] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[2__600 .GSR = "DISABLED";
    FD1S3AX \registers_6[[1__601  (.D(registers_6__1__N_1506), .CK(clk_c), 
            .Q(\registers[6] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[1__601 .GSR = "DISABLED";
    FD1S3AX \registers_6[[0__602  (.D(registers_6__0__N_1507), .CK(clk_c), 
            .Q(\registers[6] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[0__602 .GSR = "DISABLED";
    FD1S3AX \registers_6[[31__603  (.D(\registers[6] [3]), .CK(clk_c), .Q(\registers[6] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[31__603 .GSR = "DISABLED";
    FD1S3AX \registers_6[[30__604  (.D(\registers[6] [2]), .CK(clk_c), .Q(\registers[6] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[30__604 .GSR = "DISABLED";
    FD1S3AX \registers_6[[29__605  (.D(\registers[6] [1]), .CK(clk_c), .Q(\registers[6] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[29__605 .GSR = "DISABLED";
    FD1S3AX \registers_6[[28__606  (.D(\registers[6] [0]), .CK(clk_c), .Q(\registers[6] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[28__606 .GSR = "DISABLED";
    FD1S3AX \registers_6[[27__607  (.D(\registers[6] [31]), .CK(clk_c), 
            .Q(\registers[6] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[27__607 .GSR = "DISABLED";
    FD1S3AX \registers_6[[26__608  (.D(\registers[6] [30]), .CK(clk_c), 
            .Q(\registers[6] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[26__608 .GSR = "DISABLED";
    FD1S3AX \registers_6[[25__609  (.D(\registers[6] [29]), .CK(clk_c), 
            .Q(\registers[6] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[25__609 .GSR = "DISABLED";
    FD1S3AX \registers_6[[24__610  (.D(\registers[6] [28]), .CK(clk_c), 
            .Q(\registers[6] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[24__610 .GSR = "DISABLED";
    FD1S3AX \registers_6[[23__611  (.D(\registers[6] [27]), .CK(clk_c), 
            .Q(\registers[6] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[23__611 .GSR = "DISABLED";
    FD1S3AX \registers_6[[22__612  (.D(\registers[6] [26]), .CK(clk_c), 
            .Q(\registers[6] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[22__612 .GSR = "DISABLED";
    FD1S3AX \registers_6[[21__613  (.D(\registers[6] [25]), .CK(clk_c), 
            .Q(\registers[6] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[21__613 .GSR = "DISABLED";
    FD1S3AX \registers_6[[20__614  (.D(\registers[6] [24]), .CK(clk_c), 
            .Q(\registers[6] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[20__614 .GSR = "DISABLED";
    FD1S3AX \registers_6[[19__615  (.D(\registers[6] [23]), .CK(clk_c), 
            .Q(\registers[6] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[19__615 .GSR = "DISABLED";
    FD1S3AX \registers_6[[18__616  (.D(\registers[6] [22]), .CK(clk_c), 
            .Q(\registers[6] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[18__616 .GSR = "DISABLED";
    FD1S3AX \registers_6[[17__617  (.D(\registers[6] [21]), .CK(clk_c), 
            .Q(\registers[6] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[17__617 .GSR = "DISABLED";
    FD1S3AX \registers_6[[16__618  (.D(\registers[6] [20]), .CK(clk_c), 
            .Q(\registers[6] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[16__618 .GSR = "DISABLED";
    FD1S3AX \registers_6[[15__619  (.D(\registers[6] [19]), .CK(clk_c), 
            .Q(\registers[6] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[15__619 .GSR = "DISABLED";
    FD1S3AX \registers_6[[14__620  (.D(\registers[6] [18]), .CK(clk_c), 
            .Q(\registers[6] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[14__620 .GSR = "DISABLED";
    FD1S3AX \registers_6[[13__621  (.D(\registers[6] [17]), .CK(clk_c), 
            .Q(\registers[6] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[13__621 .GSR = "DISABLED";
    FD1S3AX \registers_6[[12__622  (.D(\registers[6] [16]), .CK(clk_c), 
            .Q(\registers[6] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[12__622 .GSR = "DISABLED";
    FD1S3AX \registers_6[[11__623  (.D(\registers[6] [15]), .CK(clk_c), 
            .Q(\registers[6] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[11__623 .GSR = "DISABLED";
    FD1S3AX \registers_6[[10__624  (.D(\registers[6] [14]), .CK(clk_c), 
            .Q(\registers[6] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[10__624 .GSR = "DISABLED";
    FD1S3AX \registers_6[[9__625  (.D(\registers[6] [13]), .CK(clk_c), .Q(\registers[6] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[9__625 .GSR = "DISABLED";
    FD1S3AX \registers_6[[8__626  (.D(\registers[6] [12]), .CK(clk_c), .Q(\registers[6] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[8__626 .GSR = "DISABLED";
    FD1S3AX \registers_6[[7__627  (.D(\registers[6] [11]), .CK(clk_c), .Q(\registers[6] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[7__627 .GSR = "DISABLED";
    FD1S3AX \registers_6[[6__628  (.D(\registers[6] [10]), .CK(clk_c), .Q(\registers[6] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[6__628 .GSR = "DISABLED";
    FD1S3AX \registers_6[[5__629  (.D(\registers[6] [9]), .CK(clk_c), .Q(\registers[6] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[5__629 .GSR = "DISABLED";
    FD1S3AX \registers_6[[4__630  (.D(\registers[6] [8]), .CK(clk_c), .Q(\registers[6] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[4__630 .GSR = "DISABLED";
    FD1S3AX \registers_7[[3__631  (.D(registers_7__3__N_1508), .CK(clk_c), 
            .Q(\registers[7] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[3__631 .GSR = "DISABLED";
    FD1S3AX \registers_7[[2__632  (.D(registers_7__2__N_1511), .CK(clk_c), 
            .Q(\registers[7] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[2__632 .GSR = "DISABLED";
    LUT4 i21192_3_lut (.A(\registers[8] [4]), .B(\registers[9] [4]), .C(rs1[0]), 
         .Z(n23467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21192_3_lut.init = 16'hcaca;
    FD1S3AX \registers_7[[1__633  (.D(registers_7__1__N_1512), .CK(clk_c), 
            .Q(\registers[7] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[1__633 .GSR = "DISABLED";
    FD1S3AX \registers_7[[0__634  (.D(registers_7__0__N_1513), .CK(clk_c), 
            .Q(\registers[7] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[0__634 .GSR = "DISABLED";
    FD1S3AX \registers_7[[31__635  (.D(\registers[7] [3]), .CK(clk_c), .Q(\registers[7] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[31__635 .GSR = "DISABLED";
    FD1S3AX \registers_7[[30__636  (.D(\registers[7] [2]), .CK(clk_c), .Q(\registers[7] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[30__636 .GSR = "DISABLED";
    FD1S3AX \registers_7[[29__637  (.D(\registers[7] [1]), .CK(clk_c), .Q(\registers[7] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[29__637 .GSR = "DISABLED";
    FD1S3AX \registers_7[[28__638  (.D(\registers[7] [0]), .CK(clk_c), .Q(\registers[7] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[28__638 .GSR = "DISABLED";
    FD1S3AX \registers_7[[27__639  (.D(\registers[7] [31]), .CK(clk_c), 
            .Q(\registers[7] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[27__639 .GSR = "DISABLED";
    FD1S3AX \registers_7[[26__640  (.D(\registers[7] [30]), .CK(clk_c), 
            .Q(\registers[7] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[26__640 .GSR = "DISABLED";
    FD1S3AX \registers_7[[25__641  (.D(\registers[7] [29]), .CK(clk_c), 
            .Q(\registers[7] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[25__641 .GSR = "DISABLED";
    FD1S3AX \registers_7[[24__642  (.D(\registers[7] [28]), .CK(clk_c), 
            .Q(\registers[7] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[24__642 .GSR = "DISABLED";
    FD1S3AX \registers_7[[23__643  (.D(\registers[7] [27]), .CK(clk_c), 
            .Q(\registers[7] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[23__643 .GSR = "DISABLED";
    FD1S3AX \registers_7[[22__644  (.D(\registers[7] [26]), .CK(clk_c), 
            .Q(\registers[7] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[22__644 .GSR = "DISABLED";
    FD1S3AX \registers_7[[21__645  (.D(\registers[7] [25]), .CK(clk_c), 
            .Q(\registers[7] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[21__645 .GSR = "DISABLED";
    FD1S3AX \registers_7[[20__646  (.D(\registers[7] [24]), .CK(clk_c), 
            .Q(\registers[7] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[20__646 .GSR = "DISABLED";
    FD1S3AX \registers_7[[19__647  (.D(\registers[7] [23]), .CK(clk_c), 
            .Q(\registers[7] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[19__647 .GSR = "DISABLED";
    FD1S3AX \registers_7[[18__648  (.D(\registers[7] [22]), .CK(clk_c), 
            .Q(\registers[7] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[18__648 .GSR = "DISABLED";
    FD1S3AX \registers_7[[17__649  (.D(\registers[7] [21]), .CK(clk_c), 
            .Q(\registers[7] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[17__649 .GSR = "DISABLED";
    FD1S3AX \registers_7[[16__650  (.D(\registers[7] [20]), .CK(clk_c), 
            .Q(\registers[7] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[16__650 .GSR = "DISABLED";
    FD1S3AX \registers_7[[15__651  (.D(\registers[7] [19]), .CK(clk_c), 
            .Q(\registers[7] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[15__651 .GSR = "DISABLED";
    FD1S3AX \registers_7[[14__652  (.D(\registers[7] [18]), .CK(clk_c), 
            .Q(\registers[7] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[14__652 .GSR = "DISABLED";
    FD1S3AX \registers_7[[13__653  (.D(\registers[7] [17]), .CK(clk_c), 
            .Q(\registers[7] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[13__653 .GSR = "DISABLED";
    FD1S3AX \registers_7[[12__654  (.D(\registers[7] [16]), .CK(clk_c), 
            .Q(\registers[7] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[12__654 .GSR = "DISABLED";
    FD1S3AX \registers_7[[11__655  (.D(\registers[7] [15]), .CK(clk_c), 
            .Q(\registers[7] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[11__655 .GSR = "DISABLED";
    FD1S3AX \registers_7[[10__656  (.D(\registers[7] [14]), .CK(clk_c), 
            .Q(\registers[7] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[10__656 .GSR = "DISABLED";
    FD1S3AX \registers_7[[9__657  (.D(\registers[7] [13]), .CK(clk_c), .Q(\registers[7] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[9__657 .GSR = "DISABLED";
    FD1S3AX \registers_7[[8__658  (.D(\registers[7] [12]), .CK(clk_c), .Q(\registers[7] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[8__658 .GSR = "DISABLED";
    FD1S3AX \registers_7[[7__659  (.D(\registers[7] [11]), .CK(clk_c), .Q(\registers[7] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[7__659 .GSR = "DISABLED";
    FD1S3AX \registers_7[[6__660  (.D(\registers[7] [10]), .CK(clk_c), .Q(\registers[7] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[6__660 .GSR = "DISABLED";
    FD1S3AX \registers_7[[5__661  (.D(\registers[7] [9]), .CK(clk_c), .Q(\registers[7] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[5__661 .GSR = "DISABLED";
    FD1S3AX \registers_7[[4__662  (.D(\registers[7] [8]), .CK(clk_c), .Q(\registers[7] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[4__662 .GSR = "DISABLED";
    FD1S3AX \registers_8[[3__663  (.D(registers_8__3__N_1514), .CK(clk_c), 
            .Q(\registers[8] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[3__663 .GSR = "DISABLED";
    FD1S3AX \registers_8[[2__664  (.D(registers_8__2__N_1517), .CK(clk_c), 
            .Q(\registers[8] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[2__664 .GSR = "DISABLED";
    FD1S3AX \registers_8[[1__665  (.D(registers_8__1__N_1518), .CK(clk_c), 
            .Q(\registers[8] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[1__665 .GSR = "DISABLED";
    FD1S3AX \registers_8[[0__666  (.D(registers_8__0__N_1519), .CK(clk_c), 
            .Q(\registers[8] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[0__666 .GSR = "DISABLED";
    FD1S3AX \registers_8[[31__667  (.D(\registers[8] [3]), .CK(clk_c), .Q(\registers[8] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[31__667 .GSR = "DISABLED";
    FD1S3AX \registers_8[[30__668  (.D(\registers[8] [2]), .CK(clk_c), .Q(\registers[8] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[30__668 .GSR = "DISABLED";
    FD1S3AX \registers_8[[29__669  (.D(\registers[8] [1]), .CK(clk_c), .Q(\registers[8] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[29__669 .GSR = "DISABLED";
    FD1S3AX \registers_8[[28__670  (.D(\registers[8] [0]), .CK(clk_c), .Q(\registers[8] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[28__670 .GSR = "DISABLED";
    FD1S3AX \registers_8[[27__671  (.D(\registers[8] [31]), .CK(clk_c), 
            .Q(\registers[8] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[27__671 .GSR = "DISABLED";
    FD1S3AX \registers_8[[26__672  (.D(\registers[8] [30]), .CK(clk_c), 
            .Q(\registers[8] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[26__672 .GSR = "DISABLED";
    FD1S3AX \registers_8[[25__673  (.D(\registers[8] [29]), .CK(clk_c), 
            .Q(\registers[8] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[25__673 .GSR = "DISABLED";
    FD1S3AX \registers_8[[24__674  (.D(\registers[8] [28]), .CK(clk_c), 
            .Q(\registers[8] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[24__674 .GSR = "DISABLED";
    FD1S3AX \registers_8[[23__675  (.D(\registers[8] [27]), .CK(clk_c), 
            .Q(\registers[8] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[23__675 .GSR = "DISABLED";
    FD1S3AX \registers_8[[22__676  (.D(\registers[8] [26]), .CK(clk_c), 
            .Q(\registers[8] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[22__676 .GSR = "DISABLED";
    FD1S3AX \registers_8[[21__677  (.D(\registers[8] [25]), .CK(clk_c), 
            .Q(\registers[8] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[21__677 .GSR = "DISABLED";
    FD1S3AX \registers_8[[20__678  (.D(\registers[8] [24]), .CK(clk_c), 
            .Q(\registers[8] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[20__678 .GSR = "DISABLED";
    FD1S3AX \registers_8[[19__679  (.D(\registers[8] [23]), .CK(clk_c), 
            .Q(\registers[8] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[19__679 .GSR = "DISABLED";
    FD1S3AX \registers_8[[18__680  (.D(\registers[8] [22]), .CK(clk_c), 
            .Q(\registers[8] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[18__680 .GSR = "DISABLED";
    FD1S3AX \registers_8[[17__681  (.D(\registers[8] [21]), .CK(clk_c), 
            .Q(\registers[8] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[17__681 .GSR = "DISABLED";
    FD1S3AX \registers_8[[16__682  (.D(\registers[8] [20]), .CK(clk_c), 
            .Q(\registers[8] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[16__682 .GSR = "DISABLED";
    FD1S3AX \registers_8[[15__683  (.D(\registers[8] [19]), .CK(clk_c), 
            .Q(\registers[8] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[15__683 .GSR = "DISABLED";
    FD1S3AX \registers_8[[14__684  (.D(\registers[8] [18]), .CK(clk_c), 
            .Q(\registers[8] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[14__684 .GSR = "DISABLED";
    FD1S3AX \registers_8[[13__685  (.D(\registers[8] [17]), .CK(clk_c), 
            .Q(\registers[8] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[13__685 .GSR = "DISABLED";
    FD1S3AX \registers_8[[12__686  (.D(\registers[8] [16]), .CK(clk_c), 
            .Q(\registers[8] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[12__686 .GSR = "DISABLED";
    FD1S3AX \registers_8[[11__687  (.D(\registers[8] [15]), .CK(clk_c), 
            .Q(\registers[8] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[11__687 .GSR = "DISABLED";
    FD1S3AX \registers_8[[10__688  (.D(\registers[8] [14]), .CK(clk_c), 
            .Q(\registers[8] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[10__688 .GSR = "DISABLED";
    FD1S3AX \registers_8[[9__689  (.D(\registers[8] [13]), .CK(clk_c), .Q(\registers[8] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[9__689 .GSR = "DISABLED";
    FD1S3AX \registers_8[[8__690  (.D(\registers[8] [12]), .CK(clk_c), .Q(\registers[8] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[8__690 .GSR = "DISABLED";
    FD1S3AX \registers_8[[7__691  (.D(\registers[8] [11]), .CK(clk_c), .Q(\registers[8] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[7__691 .GSR = "DISABLED";
    FD1S3AX \registers_8[[6__692  (.D(\registers[8] [10]), .CK(clk_c), .Q(\registers[8] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[6__692 .GSR = "DISABLED";
    FD1S3AX \registers_8[[5__693  (.D(\registers[8] [9]), .CK(clk_c), .Q(\registers[8] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[5__693 .GSR = "DISABLED";
    FD1S3AX \registers_8[[4__694  (.D(\registers[8] [8]), .CK(clk_c), .Q(\registers[8] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[4__694 .GSR = "DISABLED";
    FD1S3AX \registers_9[[3__695  (.D(registers_9__3__N_1520), .CK(clk_c), 
            .Q(\registers[9] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[3__695 .GSR = "DISABLED";
    FD1S3AX \registers_9[[2__696  (.D(registers_9__2__N_1523), .CK(clk_c), 
            .Q(\registers[9] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[2__696 .GSR = "DISABLED";
    FD1S3AX \registers_9[[1__697  (.D(registers_9__1__N_1524), .CK(clk_c), 
            .Q(\registers[9] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[1__697 .GSR = "DISABLED";
    FD1S3AX \registers_9[[0__698  (.D(registers_9__0__N_1525), .CK(clk_c), 
            .Q(\registers[9] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[0__698 .GSR = "DISABLED";
    FD1S3AX \registers_9[[31__699  (.D(\registers[9] [3]), .CK(clk_c), .Q(\registers[9] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[31__699 .GSR = "DISABLED";
    FD1S3AX \registers_9[[30__700  (.D(\registers[9] [2]), .CK(clk_c), .Q(\registers[9] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[30__700 .GSR = "DISABLED";
    FD1S3AX \registers_9[[29__701  (.D(\registers[9] [1]), .CK(clk_c), .Q(\registers[9] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[29__701 .GSR = "DISABLED";
    FD1S3AX \registers_9[[28__702  (.D(\registers[9] [0]), .CK(clk_c), .Q(\registers[9] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[28__702 .GSR = "DISABLED";
    FD1S3AX \registers_9[[27__703  (.D(\registers[9] [31]), .CK(clk_c), 
            .Q(\registers[9] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[27__703 .GSR = "DISABLED";
    FD1S3AX \registers_9[[26__704  (.D(\registers[9] [30]), .CK(clk_c), 
            .Q(\registers[9] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[26__704 .GSR = "DISABLED";
    FD1S3AX \registers_9[[25__705  (.D(\registers[9] [29]), .CK(clk_c), 
            .Q(\registers[9] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[25__705 .GSR = "DISABLED";
    FD1S3AX \registers_9[[24__706  (.D(\registers[9] [28]), .CK(clk_c), 
            .Q(\registers[9] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[24__706 .GSR = "DISABLED";
    FD1S3AX \registers_9[[23__707  (.D(\registers[9] [27]), .CK(clk_c), 
            .Q(\registers[9] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[23__707 .GSR = "DISABLED";
    FD1S3AX \registers_9[[22__708  (.D(\registers[9] [26]), .CK(clk_c), 
            .Q(\registers[9] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[22__708 .GSR = "DISABLED";
    FD1S3AX \registers_9[[21__709  (.D(\registers[9] [25]), .CK(clk_c), 
            .Q(\registers[9] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[21__709 .GSR = "DISABLED";
    FD1S3AX \registers_9[[20__710  (.D(\registers[9] [24]), .CK(clk_c), 
            .Q(\registers[9] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[20__710 .GSR = "DISABLED";
    FD1S3AX \registers_9[[19__711  (.D(\registers[9] [23]), .CK(clk_c), 
            .Q(\registers[9] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[19__711 .GSR = "DISABLED";
    FD1S3AX \registers_9[[18__712  (.D(\registers[9] [22]), .CK(clk_c), 
            .Q(\registers[9] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[18__712 .GSR = "DISABLED";
    FD1S3AX \registers_9[[17__713  (.D(\registers[9] [21]), .CK(clk_c), 
            .Q(\registers[9] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[17__713 .GSR = "DISABLED";
    FD1S3AX \registers_9[[16__714  (.D(\registers[9] [20]), .CK(clk_c), 
            .Q(\registers[9] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[16__714 .GSR = "DISABLED";
    FD1S3AX \registers_9[[15__715  (.D(\registers[9] [19]), .CK(clk_c), 
            .Q(\registers[9] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[15__715 .GSR = "DISABLED";
    FD1S3AX \registers_9[[14__716  (.D(\registers[9] [18]), .CK(clk_c), 
            .Q(\registers[9] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[14__716 .GSR = "DISABLED";
    FD1S3AX \registers_9[[13__717  (.D(\registers[9] [17]), .CK(clk_c), 
            .Q(\registers[9] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[13__717 .GSR = "DISABLED";
    FD1S3AX \registers_9[[12__718  (.D(\registers[9] [16]), .CK(clk_c), 
            .Q(\registers[9] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[12__718 .GSR = "DISABLED";
    FD1S3AX \registers_9[[11__719  (.D(\registers[9] [15]), .CK(clk_c), 
            .Q(\registers[9] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[11__719 .GSR = "DISABLED";
    FD1S3AX \registers_9[[10__720  (.D(\registers[9] [14]), .CK(clk_c), 
            .Q(\registers[9] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[10__720 .GSR = "DISABLED";
    FD1S3AX \registers_9[[9__721  (.D(\registers[9] [13]), .CK(clk_c), .Q(\registers[9] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[9__721 .GSR = "DISABLED";
    FD1S3AX \registers_9[[8__722  (.D(\registers[9] [12]), .CK(clk_c), .Q(\registers[9] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[8__722 .GSR = "DISABLED";
    FD1S3AX \registers_9[[7__723  (.D(\registers[9] [11]), .CK(clk_c), .Q(\registers[9] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[7__723 .GSR = "DISABLED";
    FD1S3AX \registers_9[[6__724  (.D(\registers[9] [10]), .CK(clk_c), .Q(\registers[9] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[6__724 .GSR = "DISABLED";
    FD1S3AX \registers_9[[5__725  (.D(\registers[9] [9]), .CK(clk_c), .Q(\registers[9] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[5__725 .GSR = "DISABLED";
    FD1S3AX \registers_9[[4__726  (.D(\registers[9] [8]), .CK(clk_c), .Q(\registers[9] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[4__726 .GSR = "DISABLED";
    FD1S3AX \registers_10[[3__727  (.D(registers_10__3__N_1526), .CK(clk_c), 
            .Q(\registers[10] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[3__727 .GSR = "DISABLED";
    FD1S3AX \registers_10[[2__728  (.D(registers_10__2__N_1529), .CK(clk_c), 
            .Q(\registers[10] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[2__728 .GSR = "DISABLED";
    FD1S3AX \registers_10[[1__729  (.D(registers_10__1__N_1530), .CK(clk_c), 
            .Q(\registers[10] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[1__729 .GSR = "DISABLED";
    FD1S3AX \registers_10[[0__730  (.D(registers_10__0__N_1531), .CK(clk_c), 
            .Q(\registers[10] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[0__730 .GSR = "DISABLED";
    FD1S3AX \registers_10[[31__731  (.D(\registers[10] [3]), .CK(clk_c), 
            .Q(\registers[10] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[31__731 .GSR = "DISABLED";
    FD1S3AX \registers_10[[30__732  (.D(\registers[10] [2]), .CK(clk_c), 
            .Q(\registers[10] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[30__732 .GSR = "DISABLED";
    FD1S3AX \registers_10[[29__733  (.D(\registers[10] [1]), .CK(clk_c), 
            .Q(\registers[10] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[29__733 .GSR = "DISABLED";
    FD1S3AX \registers_10[[28__734  (.D(\registers[10] [0]), .CK(clk_c), 
            .Q(\registers[10] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[28__734 .GSR = "DISABLED";
    FD1S3AX \registers_10[[27__735  (.D(\registers[10] [31]), .CK(clk_c), 
            .Q(\registers[10] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[27__735 .GSR = "DISABLED";
    FD1S3AX \registers_10[[26__736  (.D(\registers[10] [30]), .CK(clk_c), 
            .Q(\registers[10] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[26__736 .GSR = "DISABLED";
    FD1S3AX \registers_10[[25__737  (.D(\registers[10] [29]), .CK(clk_c), 
            .Q(\registers[10] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[25__737 .GSR = "DISABLED";
    FD1S3AX \registers_10[[24__738  (.D(\registers[10] [28]), .CK(clk_c), 
            .Q(\registers[10] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[24__738 .GSR = "DISABLED";
    FD1S3AX \registers_10[[23__739  (.D(\registers[10] [27]), .CK(clk_c), 
            .Q(\registers[10] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[23__739 .GSR = "DISABLED";
    FD1S3AX \registers_10[[22__740  (.D(\registers[10] [26]), .CK(clk_c), 
            .Q(\registers[10] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[22__740 .GSR = "DISABLED";
    FD1S3AX \registers_10[[21__741  (.D(\registers[10] [25]), .CK(clk_c), 
            .Q(\registers[10] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[21__741 .GSR = "DISABLED";
    FD1S3AX \registers_10[[20__742  (.D(\registers[10] [24]), .CK(clk_c), 
            .Q(\registers[10] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[20__742 .GSR = "DISABLED";
    FD1S3AX \registers_10[[19__743  (.D(\registers[10] [23]), .CK(clk_c), 
            .Q(\registers[10] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[19__743 .GSR = "DISABLED";
    FD1S3AX \registers_10[[18__744  (.D(\registers[10] [22]), .CK(clk_c), 
            .Q(\registers[10] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[18__744 .GSR = "DISABLED";
    FD1S3AX \registers_10[[17__745  (.D(\registers[10] [21]), .CK(clk_c), 
            .Q(\registers[10] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[17__745 .GSR = "DISABLED";
    FD1S3AX \registers_10[[16__746  (.D(\registers[10] [20]), .CK(clk_c), 
            .Q(\registers[10] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[16__746 .GSR = "DISABLED";
    FD1S3AX \registers_10[[15__747  (.D(\registers[10] [19]), .CK(clk_c), 
            .Q(\registers[10] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[15__747 .GSR = "DISABLED";
    FD1S3AX \registers_10[[14__748  (.D(\registers[10] [18]), .CK(clk_c), 
            .Q(\registers[10] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[14__748 .GSR = "DISABLED";
    FD1S3AX \registers_10[[13__749  (.D(\registers[10] [17]), .CK(clk_c), 
            .Q(\registers[10] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[13__749 .GSR = "DISABLED";
    FD1S3AX \registers_10[[12__750  (.D(\registers[10] [16]), .CK(clk_c), 
            .Q(\registers[10] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[12__750 .GSR = "DISABLED";
    FD1S3AX \registers_10[[11__751  (.D(\registers[10] [15]), .CK(clk_c), 
            .Q(\registers[10] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[11__751 .GSR = "DISABLED";
    FD1S3AX \registers_10[[10__752  (.D(\registers[10] [14]), .CK(clk_c), 
            .Q(\registers[10] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[10__752 .GSR = "DISABLED";
    FD1S3AX \registers_10[[9__753  (.D(\registers[10] [13]), .CK(clk_c), 
            .Q(\registers[10] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[9__753 .GSR = "DISABLED";
    FD1S3AX \registers_10[[8__754  (.D(\registers[10] [12]), .CK(clk_c), 
            .Q(\registers[10] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[8__754 .GSR = "DISABLED";
    FD1S3AX \registers_10[[7__755  (.D(\registers[10] [11]), .CK(clk_c), 
            .Q(\registers[10] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[7__755 .GSR = "DISABLED";
    FD1S3AX \registers_10[[6__756  (.D(\registers[10] [10]), .CK(clk_c), 
            .Q(\registers[10] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[6__756 .GSR = "DISABLED";
    FD1S3AX \registers_10[[5__757  (.D(\registers[10] [9]), .CK(clk_c), 
            .Q(\registers[10] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[5__757 .GSR = "DISABLED";
    FD1S3AX \registers_10[[4__758  (.D(\registers[10] [8]), .CK(clk_c), 
            .Q(\registers[10] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[4__758 .GSR = "DISABLED";
    FD1S3AX \registers_11[[3__759  (.D(registers_11__3__N_1532), .CK(clk_c), 
            .Q(\registers[11] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[3__759 .GSR = "DISABLED";
    FD1S3AX \registers_11[[2__760  (.D(registers_11__2__N_1535), .CK(clk_c), 
            .Q(\registers[11] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[2__760 .GSR = "DISABLED";
    FD1S3AX \registers_11[[1__761  (.D(registers_11__1__N_1536), .CK(clk_c), 
            .Q(\registers[11] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[1__761 .GSR = "DISABLED";
    FD1S3AX \registers_11[[0__762  (.D(registers_11__0__N_1537), .CK(clk_c), 
            .Q(\registers[11] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[0__762 .GSR = "DISABLED";
    FD1S3AX \registers_11[[31__763  (.D(\registers[11] [3]), .CK(clk_c), 
            .Q(\registers[11] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[31__763 .GSR = "DISABLED";
    FD1S3AX \registers_11[[30__764  (.D(\registers[11] [2]), .CK(clk_c), 
            .Q(\registers[11] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[30__764 .GSR = "DISABLED";
    FD1S3AX \registers_11[[29__765  (.D(\registers[11] [1]), .CK(clk_c), 
            .Q(\registers[11] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[29__765 .GSR = "DISABLED";
    FD1S3AX \registers_11[[28__766  (.D(\registers[11] [0]), .CK(clk_c), 
            .Q(\registers[11] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[28__766 .GSR = "DISABLED";
    FD1S3AX \registers_11[[27__767  (.D(\registers[11] [31]), .CK(clk_c), 
            .Q(\registers[11] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[27__767 .GSR = "DISABLED";
    FD1S3AX \registers_11[[26__768  (.D(\registers[11] [30]), .CK(clk_c), 
            .Q(\registers[11] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[26__768 .GSR = "DISABLED";
    FD1S3AX \registers_11[[25__769  (.D(\registers[11] [29]), .CK(clk_c), 
            .Q(\registers[11] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[25__769 .GSR = "DISABLED";
    FD1S3AX \registers_11[[24__770  (.D(\registers[11] [28]), .CK(clk_c), 
            .Q(\registers[11] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[24__770 .GSR = "DISABLED";
    FD1S3AX \registers_11[[23__771  (.D(\registers[11] [27]), .CK(clk_c), 
            .Q(\registers[11] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[23__771 .GSR = "DISABLED";
    FD1S3AX \registers_11[[22__772  (.D(\registers[11] [26]), .CK(clk_c), 
            .Q(\registers[11] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[22__772 .GSR = "DISABLED";
    FD1S3AX \registers_11[[21__773  (.D(\registers[11] [25]), .CK(clk_c), 
            .Q(\registers[11] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[21__773 .GSR = "DISABLED";
    FD1S3AX \registers_11[[20__774  (.D(\registers[11] [24]), .CK(clk_c), 
            .Q(\registers[11] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[20__774 .GSR = "DISABLED";
    FD1S3AX \registers_11[[19__775  (.D(\registers[11] [23]), .CK(clk_c), 
            .Q(\registers[11] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[19__775 .GSR = "DISABLED";
    FD1S3AX \registers_11[[18__776  (.D(\registers[11] [22]), .CK(clk_c), 
            .Q(\registers[11] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[18__776 .GSR = "DISABLED";
    FD1S3AX \registers_11[[17__777  (.D(\registers[11] [21]), .CK(clk_c), 
            .Q(\registers[11] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[17__777 .GSR = "DISABLED";
    FD1S3AX \registers_11[[16__778  (.D(\registers[11] [20]), .CK(clk_c), 
            .Q(\registers[11] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[16__778 .GSR = "DISABLED";
    FD1S3AX \registers_11[[15__779  (.D(\registers[11] [19]), .CK(clk_c), 
            .Q(\registers[11] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[15__779 .GSR = "DISABLED";
    FD1S3AX \registers_11[[14__780  (.D(\registers[11] [18]), .CK(clk_c), 
            .Q(\registers[11] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[14__780 .GSR = "DISABLED";
    FD1S3AX \registers_11[[13__781  (.D(\registers[11] [17]), .CK(clk_c), 
            .Q(\registers[11] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[13__781 .GSR = "DISABLED";
    FD1S3AX \registers_11[[12__782  (.D(\registers[11] [16]), .CK(clk_c), 
            .Q(\registers[11] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[12__782 .GSR = "DISABLED";
    FD1S3AX \registers_11[[11__783  (.D(\registers[11] [15]), .CK(clk_c), 
            .Q(\registers[11] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[11__783 .GSR = "DISABLED";
    FD1S3AX \registers_11[[10__784  (.D(\registers[11] [14]), .CK(clk_c), 
            .Q(\registers[11] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[10__784 .GSR = "DISABLED";
    FD1S3AX \registers_11[[9__785  (.D(\registers[11] [13]), .CK(clk_c), 
            .Q(\registers[11] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[9__785 .GSR = "DISABLED";
    FD1S3AX \registers_11[[8__786  (.D(\registers[11] [12]), .CK(clk_c), 
            .Q(\registers[11] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[8__786 .GSR = "DISABLED";
    FD1S3AX \registers_11[[7__787  (.D(\registers[11] [11]), .CK(clk_c), 
            .Q(\registers[11] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[7__787 .GSR = "DISABLED";
    FD1S3AX \registers_11[[6__788  (.D(\registers[11] [10]), .CK(clk_c), 
            .Q(\registers[11] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[6__788 .GSR = "DISABLED";
    FD1S3AX \registers_11[[5__789  (.D(\registers[11] [9]), .CK(clk_c), 
            .Q(\registers[11] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[5__789 .GSR = "DISABLED";
    FD1S3AX \registers_11[[4__790  (.D(\registers[11] [8]), .CK(clk_c), 
            .Q(\registers[11] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[4__790 .GSR = "DISABLED";
    FD1S3AX \registers_12[[3__791  (.D(registers_12__3__N_1538), .CK(clk_c), 
            .Q(\registers[12] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[3__791 .GSR = "DISABLED";
    FD1S3AX \registers_12[[2__792  (.D(registers_12__2__N_1541), .CK(clk_c), 
            .Q(\registers[12] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[2__792 .GSR = "DISABLED";
    FD1S3AX \registers_12[[1__793  (.D(registers_12__1__N_1542), .CK(clk_c), 
            .Q(\registers[12] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[1__793 .GSR = "DISABLED";
    FD1S3AX \registers_12[[0__794  (.D(registers_12__0__N_1543), .CK(clk_c), 
            .Q(\registers[12] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[0__794 .GSR = "DISABLED";
    FD1S3AX \registers_12[[31__795  (.D(\registers[12] [3]), .CK(clk_c), 
            .Q(\registers[12] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[31__795 .GSR = "DISABLED";
    FD1S3AX \registers_12[[30__796  (.D(\registers[12] [2]), .CK(clk_c), 
            .Q(\registers[12] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[30__796 .GSR = "DISABLED";
    FD1S3AX \registers_12[[29__797  (.D(\registers[12] [1]), .CK(clk_c), 
            .Q(\registers[12] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[29__797 .GSR = "DISABLED";
    FD1S3AX \registers_12[[28__798  (.D(\registers[12] [0]), .CK(clk_c), 
            .Q(\registers[12] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[28__798 .GSR = "DISABLED";
    FD1S3AX \registers_12[[27__799  (.D(\registers[12] [31]), .CK(clk_c), 
            .Q(\registers[12] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[27__799 .GSR = "DISABLED";
    FD1S3AX \registers_12[[26__800  (.D(\registers[12] [30]), .CK(clk_c), 
            .Q(\registers[12] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[26__800 .GSR = "DISABLED";
    FD1S3AX \registers_12[[25__801  (.D(\registers[12] [29]), .CK(clk_c), 
            .Q(\registers[12] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[25__801 .GSR = "DISABLED";
    FD1S3AX \registers_12[[24__802  (.D(\registers[12] [28]), .CK(clk_c), 
            .Q(\registers[12] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[24__802 .GSR = "DISABLED";
    FD1S3AX \registers_12[[23__803  (.D(\registers[12] [27]), .CK(clk_c), 
            .Q(\registers[12] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[23__803 .GSR = "DISABLED";
    FD1S3AX \registers_12[[22__804  (.D(\registers[12] [26]), .CK(clk_c), 
            .Q(\registers[12] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[22__804 .GSR = "DISABLED";
    FD1S3AX \registers_12[[21__805  (.D(\registers[12] [25]), .CK(clk_c), 
            .Q(\registers[12] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[21__805 .GSR = "DISABLED";
    FD1S3AX \registers_12[[20__806  (.D(\registers[12] [24]), .CK(clk_c), 
            .Q(\registers[12] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[20__806 .GSR = "DISABLED";
    FD1S3AX \registers_12[[19__807  (.D(\registers[12] [23]), .CK(clk_c), 
            .Q(\registers[12] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[19__807 .GSR = "DISABLED";
    FD1S3AX \registers_12[[18__808  (.D(\registers[12] [22]), .CK(clk_c), 
            .Q(\registers[12] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[18__808 .GSR = "DISABLED";
    FD1S3AX \registers_12[[17__809  (.D(\registers[12] [21]), .CK(clk_c), 
            .Q(\registers[12] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[17__809 .GSR = "DISABLED";
    FD1S3AX \registers_12[[16__810  (.D(\registers[12] [20]), .CK(clk_c), 
            .Q(\registers[12] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[16__810 .GSR = "DISABLED";
    FD1S3AX \registers_12[[15__811  (.D(\registers[12] [19]), .CK(clk_c), 
            .Q(\registers[12] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[15__811 .GSR = "DISABLED";
    FD1S3AX \registers_12[[14__812  (.D(\registers[12] [18]), .CK(clk_c), 
            .Q(\registers[12] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[14__812 .GSR = "DISABLED";
    FD1S3AX \registers_12[[13__813  (.D(\registers[12] [17]), .CK(clk_c), 
            .Q(\registers[12] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[13__813 .GSR = "DISABLED";
    FD1S3AX \registers_12[[12__814  (.D(\registers[12] [16]), .CK(clk_c), 
            .Q(\registers[12] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[12__814 .GSR = "DISABLED";
    FD1S3AX \registers_12[[11__815  (.D(\registers[12] [15]), .CK(clk_c), 
            .Q(\registers[12] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[11__815 .GSR = "DISABLED";
    FD1S3AX \registers_12[[10__816  (.D(\registers[12] [14]), .CK(clk_c), 
            .Q(\registers[12] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[10__816 .GSR = "DISABLED";
    FD1S3AX \registers_12[[9__817  (.D(\registers[12] [13]), .CK(clk_c), 
            .Q(\registers[12] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[9__817 .GSR = "DISABLED";
    FD1S3AX \registers_12[[8__818  (.D(\registers[12] [12]), .CK(clk_c), 
            .Q(\registers[12] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[8__818 .GSR = "DISABLED";
    FD1S3AX \registers_12[[7__819  (.D(\registers[12] [11]), .CK(clk_c), 
            .Q(\registers[12] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[7__819 .GSR = "DISABLED";
    FD1S3AX \registers_12[[6__820  (.D(\registers[12] [10]), .CK(clk_c), 
            .Q(\registers[12] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[6__820 .GSR = "DISABLED";
    FD1S3AX \registers_12[[5__821  (.D(\registers[12] [9]), .CK(clk_c), 
            .Q(\registers[12] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[5__821 .GSR = "DISABLED";
    FD1S3AX \registers_12[[4__822  (.D(\registers[12] [8]), .CK(clk_c), 
            .Q(\registers[12] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[4__822 .GSR = "DISABLED";
    FD1S3AX \registers_13[[3__823  (.D(registers_13__3__N_1544), .CK(clk_c), 
            .Q(\registers[13] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[3__823 .GSR = "DISABLED";
    FD1S3AX \registers_13[[2__824  (.D(registers_13__2__N_1547), .CK(clk_c), 
            .Q(\registers[13] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[2__824 .GSR = "DISABLED";
    FD1S3AX \registers_13[[1__825  (.D(registers_13__1__N_1548), .CK(clk_c), 
            .Q(\registers[13] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[1__825 .GSR = "DISABLED";
    FD1S3AX \registers_13[[0__826  (.D(registers_13__0__N_1549), .CK(clk_c), 
            .Q(\registers[13] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[0__826 .GSR = "DISABLED";
    FD1S3AX \registers_13[[31__827  (.D(\registers[13] [3]), .CK(clk_c), 
            .Q(\registers[13] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[31__827 .GSR = "DISABLED";
    FD1S3AX \registers_13[[30__828  (.D(\registers[13] [2]), .CK(clk_c), 
            .Q(\registers[13] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[30__828 .GSR = "DISABLED";
    FD1S3AX \registers_13[[29__829  (.D(\registers[13] [1]), .CK(clk_c), 
            .Q(\registers[13] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[29__829 .GSR = "DISABLED";
    FD1S3AX \registers_13[[28__830  (.D(\registers[13] [0]), .CK(clk_c), 
            .Q(\registers[13] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[28__830 .GSR = "DISABLED";
    FD1S3AX \registers_13[[27__831  (.D(\registers[13] [31]), .CK(clk_c), 
            .Q(\registers[13] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[27__831 .GSR = "DISABLED";
    FD1S3AX \registers_13[[26__832  (.D(\registers[13] [30]), .CK(clk_c), 
            .Q(\registers[13] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[26__832 .GSR = "DISABLED";
    FD1S3AX \registers_13[[25__833  (.D(\registers[13] [29]), .CK(clk_c), 
            .Q(\registers[13] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[25__833 .GSR = "DISABLED";
    FD1S3AX \registers_13[[24__834  (.D(\registers[13] [28]), .CK(clk_c), 
            .Q(\registers[13] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[24__834 .GSR = "DISABLED";
    FD1S3AX \registers_13[[23__835  (.D(\registers[13] [27]), .CK(clk_c), 
            .Q(\registers[13] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[23__835 .GSR = "DISABLED";
    FD1S3AX \registers_13[[22__836  (.D(\registers[13] [26]), .CK(clk_c), 
            .Q(\registers[13] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[22__836 .GSR = "DISABLED";
    FD1S3AX \registers_13[[21__837  (.D(\registers[13] [25]), .CK(clk_c), 
            .Q(\registers[13] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[21__837 .GSR = "DISABLED";
    FD1S3AX \registers_13[[20__838  (.D(\registers[13] [24]), .CK(clk_c), 
            .Q(\registers[13] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[20__838 .GSR = "DISABLED";
    FD1S3AX \registers_13[[19__839  (.D(\registers[13] [23]), .CK(clk_c), 
            .Q(\registers[13] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[19__839 .GSR = "DISABLED";
    FD1S3AX \registers_13[[18__840  (.D(\registers[13] [22]), .CK(clk_c), 
            .Q(\registers[13] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[18__840 .GSR = "DISABLED";
    FD1S3AX \registers_13[[17__841  (.D(\registers[13] [21]), .CK(clk_c), 
            .Q(\registers[13] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[17__841 .GSR = "DISABLED";
    FD1S3AX \registers_13[[16__842  (.D(\registers[13] [20]), .CK(clk_c), 
            .Q(\registers[13] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[16__842 .GSR = "DISABLED";
    FD1S3AX \registers_13[[15__843  (.D(\registers[13] [19]), .CK(clk_c), 
            .Q(\registers[13] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[15__843 .GSR = "DISABLED";
    FD1S3AX \registers_13[[14__844  (.D(\registers[13] [18]), .CK(clk_c), 
            .Q(\registers[13] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[14__844 .GSR = "DISABLED";
    FD1S3AX \registers_13[[13__845  (.D(\registers[13] [17]), .CK(clk_c), 
            .Q(\registers[13] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[13__845 .GSR = "DISABLED";
    FD1S3AX \registers_13[[12__846  (.D(\registers[13] [16]), .CK(clk_c), 
            .Q(\registers[13] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[12__846 .GSR = "DISABLED";
    FD1S3AX \registers_13[[11__847  (.D(\registers[13] [15]), .CK(clk_c), 
            .Q(\registers[13] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[11__847 .GSR = "DISABLED";
    FD1S3AX \registers_13[[10__848  (.D(\registers[13] [14]), .CK(clk_c), 
            .Q(\registers[13] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[10__848 .GSR = "DISABLED";
    FD1S3AX \registers_13[[9__849  (.D(\registers[13] [13]), .CK(clk_c), 
            .Q(\registers[13] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[9__849 .GSR = "DISABLED";
    FD1S3AX \registers_13[[8__850  (.D(\registers[13] [12]), .CK(clk_c), 
            .Q(\registers[13] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[8__850 .GSR = "DISABLED";
    FD1S3AX \registers_13[[7__851  (.D(\registers[13] [11]), .CK(clk_c), 
            .Q(\registers[13] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[7__851 .GSR = "DISABLED";
    FD1S3AX \registers_13[[6__852  (.D(\registers[13] [10]), .CK(clk_c), 
            .Q(\registers[13] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[6__852 .GSR = "DISABLED";
    FD1S3AX \registers_13[[5__853  (.D(\registers[13] [9]), .CK(clk_c), 
            .Q(\registers[13] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[5__853 .GSR = "DISABLED";
    FD1S3AX \registers_13[[4__854  (.D(\registers[13] [8]), .CK(clk_c), 
            .Q(\registers[13] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[4__854 .GSR = "DISABLED";
    FD1S3AX \registers_14[[3__855  (.D(registers_14__3__N_1550), .CK(clk_c), 
            .Q(\registers[14] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[3__855 .GSR = "DISABLED";
    FD1S3AX \registers_14[[2__856  (.D(registers_14__2__N_1553), .CK(clk_c), 
            .Q(\registers[14] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[2__856 .GSR = "DISABLED";
    FD1S3AX \registers_14[[1__857  (.D(registers_14__1__N_1554), .CK(clk_c), 
            .Q(\registers[14] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[1__857 .GSR = "DISABLED";
    FD1S3AX \registers_14[[0__858  (.D(registers_14__0__N_1555), .CK(clk_c), 
            .Q(\registers[14] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[0__858 .GSR = "DISABLED";
    FD1S3AX \registers_14[[31__859  (.D(\registers[14] [3]), .CK(clk_c), 
            .Q(\registers[14] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[31__859 .GSR = "DISABLED";
    FD1S3AX \registers_14[[30__860  (.D(\registers[14] [2]), .CK(clk_c), 
            .Q(\registers[14] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[30__860 .GSR = "DISABLED";
    FD1S3AX \registers_14[[29__861  (.D(\registers[14] [1]), .CK(clk_c), 
            .Q(\registers[14] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[29__861 .GSR = "DISABLED";
    FD1S3AX \registers_14[[28__862  (.D(\registers[14] [0]), .CK(clk_c), 
            .Q(\registers[14] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[28__862 .GSR = "DISABLED";
    FD1S3AX \registers_14[[27__863  (.D(\registers[14] [31]), .CK(clk_c), 
            .Q(\registers[14] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[27__863 .GSR = "DISABLED";
    FD1S3AX \registers_14[[26__864  (.D(\registers[14] [30]), .CK(clk_c), 
            .Q(\registers[14] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[26__864 .GSR = "DISABLED";
    FD1S3AX \registers_14[[25__865  (.D(\registers[14] [29]), .CK(clk_c), 
            .Q(\registers[14] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[25__865 .GSR = "DISABLED";
    FD1S3AX \registers_14[[24__866  (.D(\registers[14] [28]), .CK(clk_c), 
            .Q(\registers[14] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[24__866 .GSR = "DISABLED";
    FD1S3AX \registers_14[[23__867  (.D(\registers[14] [27]), .CK(clk_c), 
            .Q(\registers[14] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[23__867 .GSR = "DISABLED";
    FD1S3AX \registers_14[[22__868  (.D(\registers[14] [26]), .CK(clk_c), 
            .Q(\registers[14] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[22__868 .GSR = "DISABLED";
    FD1S3AX \registers_14[[21__869  (.D(\registers[14] [25]), .CK(clk_c), 
            .Q(\registers[14] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[21__869 .GSR = "DISABLED";
    FD1S3AX \registers_14[[20__870  (.D(\registers[14] [24]), .CK(clk_c), 
            .Q(\registers[14] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[20__870 .GSR = "DISABLED";
    FD1S3AX \registers_14[[19__871  (.D(\registers[14] [23]), .CK(clk_c), 
            .Q(\registers[14] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[19__871 .GSR = "DISABLED";
    FD1S3AX \registers_14[[18__872  (.D(\registers[14] [22]), .CK(clk_c), 
            .Q(\registers[14] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[18__872 .GSR = "DISABLED";
    FD1S3AX \registers_14[[17__873  (.D(\registers[14] [21]), .CK(clk_c), 
            .Q(\registers[14] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[17__873 .GSR = "DISABLED";
    FD1S3AX \registers_14[[16__874  (.D(\registers[14] [20]), .CK(clk_c), 
            .Q(\registers[14] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[16__874 .GSR = "DISABLED";
    FD1S3AX \registers_14[[15__875  (.D(\registers[14] [19]), .CK(clk_c), 
            .Q(\registers[14] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[15__875 .GSR = "DISABLED";
    FD1S3AX \registers_14[[14__876  (.D(\registers[14] [18]), .CK(clk_c), 
            .Q(\registers[14] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[14__876 .GSR = "DISABLED";
    FD1S3AX \registers_14[[13__877  (.D(\registers[14] [17]), .CK(clk_c), 
            .Q(\registers[14] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[13__877 .GSR = "DISABLED";
    FD1S3AX \registers_14[[12__878  (.D(\registers[14] [16]), .CK(clk_c), 
            .Q(\registers[14] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[12__878 .GSR = "DISABLED";
    FD1S3AX \registers_14[[11__879  (.D(\registers[14] [15]), .CK(clk_c), 
            .Q(\registers[14] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[11__879 .GSR = "DISABLED";
    FD1S3AX \registers_14[[10__880  (.D(\registers[14] [14]), .CK(clk_c), 
            .Q(\registers[14] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[10__880 .GSR = "DISABLED";
    FD1S3AX \registers_14[[9__881  (.D(\registers[14] [13]), .CK(clk_c), 
            .Q(\registers[14] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[9__881 .GSR = "DISABLED";
    FD1S3AX \registers_14[[8__882  (.D(\registers[14] [12]), .CK(clk_c), 
            .Q(\registers[14] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[8__882 .GSR = "DISABLED";
    FD1S3AX \registers_14[[7__883  (.D(\registers[14] [11]), .CK(clk_c), 
            .Q(\registers[14] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[7__883 .GSR = "DISABLED";
    FD1S3AX \registers_14[[6__884  (.D(\registers[14] [10]), .CK(clk_c), 
            .Q(\registers[14] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[6__884 .GSR = "DISABLED";
    FD1S3AX \registers_14[[5__885  (.D(\registers[14] [9]), .CK(clk_c), 
            .Q(\registers[14] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[5__885 .GSR = "DISABLED";
    FD1S3AX \registers_14[[4__886  (.D(\registers[14] [8]), .CK(clk_c), 
            .Q(\registers[14] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[4__886 .GSR = "DISABLED";
    FD1S3AX \registers_15[[3__887  (.D(registers_15__3__N_1556), .CK(clk_c), 
            .Q(\registers[15] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[3__887 .GSR = "DISABLED";
    FD1S3AX \registers_15[[2__888  (.D(registers_15__2__N_1559), .CK(clk_c), 
            .Q(\registers[15] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[2__888 .GSR = "DISABLED";
    FD1S3AX \registers_15[[1__889  (.D(registers_15__1__N_1560), .CK(clk_c), 
            .Q(\registers[15] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[1__889 .GSR = "DISABLED";
    FD1S3AX \registers_15[[0__890  (.D(registers_15__0__N_1561), .CK(clk_c), 
            .Q(\registers[15] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[0__890 .GSR = "DISABLED";
    FD1S3AX \registers_15[[31__891  (.D(\registers[15] [3]), .CK(clk_c), 
            .Q(\registers[15] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[31__891 .GSR = "DISABLED";
    FD1S3AX \registers_15[[30__892  (.D(\registers[15] [2]), .CK(clk_c), 
            .Q(\registers[15] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[30__892 .GSR = "DISABLED";
    FD1S3AX \registers_15[[29__893  (.D(\registers[15] [1]), .CK(clk_c), 
            .Q(\registers[15] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[29__893 .GSR = "DISABLED";
    FD1S3AX \registers_15[[28__894  (.D(\registers[15] [0]), .CK(clk_c), 
            .Q(\registers[15] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[28__894 .GSR = "DISABLED";
    FD1S3AX \registers_15[[27__895  (.D(\registers[15] [31]), .CK(clk_c), 
            .Q(\registers[15] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[27__895 .GSR = "DISABLED";
    FD1S3AX \registers_15[[26__896  (.D(\registers[15] [30]), .CK(clk_c), 
            .Q(\registers[15] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[26__896 .GSR = "DISABLED";
    FD1S3AX \registers_15[[25__897  (.D(\registers[15] [29]), .CK(clk_c), 
            .Q(\registers[15] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[25__897 .GSR = "DISABLED";
    FD1S3AX \registers_15[[24__898  (.D(\registers[15] [28]), .CK(clk_c), 
            .Q(\registers[15] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[24__898 .GSR = "DISABLED";
    FD1S3AX \registers_15[[23__899  (.D(\registers[15] [27]), .CK(clk_c), 
            .Q(\registers[15] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[23__899 .GSR = "DISABLED";
    FD1S3AX \registers_15[[22__900  (.D(\registers[15] [26]), .CK(clk_c), 
            .Q(\registers[15] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[22__900 .GSR = "DISABLED";
    FD1S3AX \registers_15[[21__901  (.D(\registers[15] [25]), .CK(clk_c), 
            .Q(\registers[15] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[21__901 .GSR = "DISABLED";
    FD1S3AX \registers_15[[20__902  (.D(\registers[15] [24]), .CK(clk_c), 
            .Q(\registers[15] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[20__902 .GSR = "DISABLED";
    FD1S3AX \registers_15[[19__903  (.D(\registers[15] [23]), .CK(clk_c), 
            .Q(\registers[15] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[19__903 .GSR = "DISABLED";
    FD1S3AX \registers_15[[18__904  (.D(\registers[15] [22]), .CK(clk_c), 
            .Q(\registers[15] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[18__904 .GSR = "DISABLED";
    FD1S3AX \registers_15[[17__905  (.D(\registers[15] [21]), .CK(clk_c), 
            .Q(\registers[15] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[17__905 .GSR = "DISABLED";
    FD1S3AX \registers_15[[16__906  (.D(\registers[15] [20]), .CK(clk_c), 
            .Q(\registers[15] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[16__906 .GSR = "DISABLED";
    FD1S3AX \registers_15[[15__907  (.D(\registers[15] [19]), .CK(clk_c), 
            .Q(\registers[15] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[15__907 .GSR = "DISABLED";
    FD1S3AX \registers_15[[14__908  (.D(\registers[15] [18]), .CK(clk_c), 
            .Q(\registers[15] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[14__908 .GSR = "DISABLED";
    FD1S3AX \registers_15[[13__909  (.D(\registers[15] [17]), .CK(clk_c), 
            .Q(\registers[15] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[13__909 .GSR = "DISABLED";
    FD1S3AX \registers_15[[12__910  (.D(\registers[15] [16]), .CK(clk_c), 
            .Q(\registers[15] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[12__910 .GSR = "DISABLED";
    FD1S3AX \registers_15[[11__911  (.D(\registers[15] [15]), .CK(clk_c), 
            .Q(\registers[15] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[11__911 .GSR = "DISABLED";
    FD1S3AX \registers_15[[10__912  (.D(\registers[15] [14]), .CK(clk_c), 
            .Q(\registers[15] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[10__912 .GSR = "DISABLED";
    FD1S3AX \registers_15[[9__913  (.D(\registers[15] [13]), .CK(clk_c), 
            .Q(\registers[15] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[9__913 .GSR = "DISABLED";
    FD1S3AX \registers_15[[8__914  (.D(\registers[15] [12]), .CK(clk_c), 
            .Q(\registers[15] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[8__914 .GSR = "DISABLED";
    FD1S3AX \registers_15[[7__915  (.D(\registers[15] [11]), .CK(clk_c), 
            .Q(\registers[15] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[7__915 .GSR = "DISABLED";
    FD1S3AX \registers_15[[6__916  (.D(\registers[15] [10]), .CK(clk_c), 
            .Q(\registers[15] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[6__916 .GSR = "DISABLED";
    FD1S3AX \registers_15[[5__917  (.D(\registers[15] [9]), .CK(clk_c), 
            .Q(\registers[15] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[5__917 .GSR = "DISABLED";
    FD1S3AX \registers_15[[4__918  (.D(\registers[15] [8]), .CK(clk_c), 
            .Q(\registers[15] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[4__918 .GSR = "DISABLED";
    FD1S3AX \registers_1[[3__503  (.D(registers_1__3__N_1484), .CK(clk_c), 
            .Q(\registers[1] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[3__503 .GSR = "DISABLED";
    LUT4 i21191_3_lut (.A(\registers[6] [4]), .B(\registers[7] [4]), .C(rs1[0]), 
         .Z(n23466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21191_3_lut.init = 16'hcaca;
    LUT4 i21190_3_lut (.A(\registers[5] [4]), .B(rs1[0]), .Z(n23465)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21190_3_lut.init = 16'h8888;
    LUT4 i21180_3_lut (.A(\registers[14] [4]), .B(\registers[15] [4]), .C(rs2[0]), 
         .Z(n23455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21180_3_lut.init = 16'hcaca;
    LUT4 i21179_3_lut (.A(\registers[12] [4]), .B(\registers[13] [4]), .C(rs2[0]), 
         .Z(n23454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21179_3_lut.init = 16'hcaca;
    LUT4 i21178_3_lut (.A(\registers[10] [4]), .B(\registers[11] [4]), .C(rs2[0]), 
         .Z(n23453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21178_3_lut.init = 16'hcaca;
    LUT4 i21177_3_lut (.A(\registers[8] [4]), .B(\registers[9] [4]), .C(rs2[0]), 
         .Z(n23452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21177_3_lut.init = 16'hcaca;
    LUT4 i21176_3_lut (.A(\registers[6] [4]), .B(\registers[7] [4]), .C(rs2[0]), 
         .Z(n23451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21176_3_lut.init = 16'hcaca;
    LUT4 i21175_3_lut (.A(\registers[5] [4]), .B(rs2[0]), .Z(n23450)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21175_3_lut.init = 16'h8888;
    LUT4 registers_15__7__I_0_3_lut_4_lut (.A(n25377), .B(n25184), .C(debug_rd[3]), 
         .D(\registers[15] [7]), .Z(registers_15__3__N_1556)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_15__6__I_0_3_lut_4_lut (.A(n25377), .B(n25184), .C(debug_rd[2]), 
         .D(\registers[15] [6]), .Z(registers_15__2__N_1559)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_15__5__I_0_3_lut_4_lut (.A(n25377), .B(n25184), .C(debug_rd[1]), 
         .D(\registers[15] [5]), .Z(registers_15__1__N_1560)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_15__4__I_0_3_lut_4_lut (.A(n25377), .B(n25184), .C(debug_rd[0]), 
         .D(\registers[15] [4]), .Z(registers_15__0__N_1561)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__7__I_0_3_lut_4_lut (.A(n25377), .B(n25185), .C(debug_rd[3]), 
         .D(\registers[14] [7]), .Z(registers_14__3__N_1550)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__6__I_0_3_lut_4_lut (.A(n25377), .B(n25185), .C(debug_rd[2]), 
         .D(\registers[14] [6]), .Z(registers_14__2__N_1553)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__5__I_0_3_lut_4_lut (.A(n25377), .B(n25185), .C(debug_rd[1]), 
         .D(\registers[14] [5]), .Z(registers_14__1__N_1554)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_14__4__I_0_3_lut_4_lut (.A(n25377), .B(n25185), .C(debug_rd[0]), 
         .D(\registers[14] [4]), .Z(registers_14__0__N_1555)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i21144_3_lut (.A(n23417), .B(n23418), .C(rs1[3]), .Z(data_rs1[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21144_3_lut.init = 16'hcaca;
    LUT4 registers_13__7__I_0_3_lut_4_lut (.A(n25377), .B(n25186), .C(debug_rd[3]), 
         .D(\registers[13] [7]), .Z(registers_13__3__N_1544)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__6__I_0_3_lut_4_lut (.A(n25377), .B(n25186), .C(debug_rd[2]), 
         .D(\registers[13] [6]), .Z(registers_13__2__N_1547)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__5__I_0_3_lut_4_lut (.A(n25377), .B(n25186), .C(debug_rd[1]), 
         .D(\registers[13] [5]), .Z(registers_13__1__N_1548)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__4__I_0_3_lut_4_lut (.A(n25377), .B(n25186), .C(debug_rd[0]), 
         .D(\registers[13] [4]), .Z(registers_13__0__N_1549)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__7__I_0_3_lut_4_lut (.A(n25377), .B(n25183), .C(debug_rd[3]), 
         .D(\registers[12] [7]), .Z(registers_12__3__N_1538)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__6__I_0_3_lut_4_lut (.A(n25377), .B(n25183), .C(debug_rd[2]), 
         .D(\registers[12] [6]), .Z(registers_12__2__N_1541)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__5__I_0_3_lut_4_lut (.A(n25377), .B(n25183), .C(debug_rd[1]), 
         .D(\registers[12] [5]), .Z(registers_12__1__N_1542)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 rs1_3__I_0_Mux_1_i12_3_lut (.A(\registers[14] [5]), .B(\registers[15] [5]), 
         .C(rs1[0]), .Z(n12_adj_2335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i12_3_lut.init = 16'hcaca;
    LUT4 registers_12__4__I_0_3_lut_4_lut (.A(n25377), .B(n25183), .C(debug_rd[0]), 
         .D(\registers[12] [4]), .Z(registers_12__0__N_1543)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_11__7__I_0_3_lut_4_lut (.A(n25379), .B(n25184), .C(debug_rd[3]), 
         .D(\registers[11] [7]), .Z(registers_11__3__N_1532)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__6__I_0_3_lut_4_lut (.A(n25379), .B(n25184), .C(debug_rd[2]), 
         .D(\registers[11] [6]), .Z(registers_11__2__N_1535)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs1_3__I_0_Mux_1_i11_3_lut (.A(\registers[12] [5]), .B(\registers[13] [5]), 
         .C(rs1[0]), .Z(n11_adj_2336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i11_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i9_3_lut (.A(\registers[10] [5]), .B(\registers[11] [5]), 
         .C(rs1[0]), .Z(n9_adj_2337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i8_3_lut (.A(\registers[8] [5]), .B(\registers[9] [5]), 
         .C(rs1[0]), .Z(n8_adj_2338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i8_3_lut.init = 16'hcaca;
    LUT4 registers_11__5__I_0_3_lut_4_lut (.A(n25379), .B(n25184), .C(debug_rd[1]), 
         .D(\registers[11] [5]), .Z(registers_11__1__N_1536)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__4__I_0_3_lut_4_lut (.A(n25379), .B(n25184), .C(debug_rd[0]), 
         .D(\registers[11] [4]), .Z(registers_11__0__N_1537)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs1_3__I_0_Mux_1_i5_3_lut (.A(\registers[6] [5]), .B(\registers[7] [5]), 
         .C(rs1[0]), .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 registers_10__7__I_0_3_lut_4_lut (.A(n25379), .B(n25185), .C(debug_rd[3]), 
         .D(\registers[10] [7]), .Z(registers_10__3__N_1526)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__6__I_0_3_lut_4_lut (.A(n25379), .B(n25185), .C(debug_rd[2]), 
         .D(\registers[10] [6]), .Z(registers_10__2__N_1529)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs2_3__I_0_Mux_1_i12_3_lut (.A(\registers[14] [5]), .B(\registers[15] [5]), 
         .C(rs2[0]), .Z(n12_adj_2339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i12_3_lut.init = 16'hcaca;
    LUT4 registers_10__5__I_0_3_lut_4_lut (.A(n25379), .B(n25185), .C(debug_rd[1]), 
         .D(\registers[10] [5]), .Z(registers_10__1__N_1530)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs2_3__I_0_Mux_1_i11_3_lut (.A(\registers[12] [5]), .B(\registers[13] [5]), 
         .C(rs2[0]), .Z(n11_adj_2340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i11_3_lut.init = 16'hcaca;
    LUT4 registers_10__4__I_0_3_lut_4_lut (.A(n25379), .B(n25185), .C(debug_rd[0]), 
         .D(\registers[10] [4]), .Z(registers_10__0__N_1531)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__7__I_0_3_lut_4_lut (.A(n25379), .B(n25186), .C(debug_rd[3]), 
         .D(\registers[9] [7]), .Z(registers_9__3__N_1520)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs2_3__I_0_Mux_1_i9_3_lut (.A(\registers[10] [5]), .B(\registers[11] [5]), 
         .C(rs2[0]), .Z(n9_adj_2341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i8_3_lut (.A(\registers[8] [5]), .B(\registers[9] [5]), 
         .C(rs2[0]), .Z(n8_adj_2342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i8_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i5_3_lut (.A(\registers[6] [5]), .B(\registers[7] [5]), 
         .C(rs2[0]), .Z(n5_adj_2343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 registers_9__6__I_0_3_lut_4_lut (.A(n25379), .B(n25186), .C(debug_rd[2]), 
         .D(\registers[9] [6]), .Z(registers_9__2__N_1523)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__5__I_0_3_lut_4_lut (.A(n25379), .B(n25186), .C(debug_rd[1]), 
         .D(\registers[9] [5]), .Z(registers_9__1__N_1524)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__4__I_0_3_lut_4_lut (.A(n25379), .B(n25186), .C(debug_rd[0]), 
         .D(\registers[9] [4]), .Z(registers_9__0__N_1525)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__7__I_0_3_lut_4_lut (.A(n25379), .B(n25183), .C(debug_rd[3]), 
         .D(\registers[8] [7]), .Z(registers_8__3__N_1514)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__6__I_0_3_lut_4_lut (.A(n25379), .B(n25183), .C(debug_rd[2]), 
         .D(\registers[8] [6]), .Z(registers_8__2__N_1517)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__5__I_0_3_lut_4_lut (.A(n25379), .B(n25183), .C(debug_rd[1]), 
         .D(\registers[8] [5]), .Z(registers_8__1__N_1518)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__4__I_0_3_lut_4_lut (.A(n25379), .B(n25183), .C(debug_rd[0]), 
         .D(\registers[8] [4]), .Z(registers_8__0__N_1519)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__7__I_0_3_lut_4_lut (.A(n25380), .B(n25184), .C(debug_rd[3]), 
         .D(\registers[7] [7]), .Z(registers_7__3__N_1508)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__6__I_0_3_lut_4_lut (.A(n25380), .B(n25184), .C(debug_rd[2]), 
         .D(\registers[7] [6]), .Z(registers_7__2__N_1511)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__5__I_0_3_lut_4_lut (.A(n25380), .B(n25184), .C(debug_rd[1]), 
         .D(\registers[7] [5]), .Z(registers_7__1__N_1512)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__4__I_0_3_lut_4_lut (.A(n25380), .B(n25184), .C(debug_rd[0]), 
         .D(\registers[7] [4]), .Z(registers_7__0__N_1513)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__7__I_0_3_lut_4_lut (.A(n25380), .B(n25185), .C(debug_rd[3]), 
         .D(\registers[6] [7]), .Z(registers_6__3__N_1502)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__6__I_0_3_lut_4_lut (.A(n25380), .B(n25185), .C(debug_rd[2]), 
         .D(\registers[6] [6]), .Z(registers_6__2__N_1505)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__5__I_0_3_lut_4_lut (.A(n25380), .B(n25185), .C(debug_rd[1]), 
         .D(\registers[6] [5]), .Z(registers_6__1__N_1506)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__4__I_0_3_lut_4_lut (.A(n25380), .B(n25185), .C(debug_rd[0]), 
         .D(\registers[6] [4]), .Z(registers_6__0__N_1507)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__6__I_0_3_lut_4_lut (.A(n25380), .B(n25186), .C(debug_rd[2]), 
         .D(\registers[5] [6]), .Z(registers_5__2__N_1499)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__4__I_0_3_lut_4_lut (.A(n25380), .B(n25186), .C(debug_rd[0]), 
         .D(\registers[5] [4]), .Z(registers_5__0__N_1501)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 rs2_3__I_0_Mux_3_i5_3_lut (.A(\registers[6] [7]), .B(\registers[7] [7]), 
         .C(rs2[0]), .Z(n5_adj_2344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i4_3_lut (.A(\reg_access[4][3] ), .B(\registers[5] [7]), 
         .C(rs2[0]), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i4_3_lut.init = 16'hcaca;
    LUT4 i21388_3_lut (.A(n4), .B(n5_adj_2344), .C(rs2[1]), .Z(n23568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21388_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i5_3_lut (.A(\registers[6] [7]), .B(\registers[7] [7]), 
         .C(rs1[0]), .Z(n5_adj_2345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i4_3_lut (.A(\reg_access[4][3] ), .B(\registers[5] [7]), 
         .C(rs1[0]), .Z(n4_adj_2346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i4_3_lut.init = 16'hcaca;
    LUT4 i21390_3_lut (.A(n4_adj_2346), .B(n5_adj_2345), .C(rs1[1]), .Z(n23561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21390_3_lut.init = 16'hcaca;
    LUT4 registers_5__5__I_0_3_lut_4_lut (.A(n25380), .B(n25186), .C(debug_rd[1]), 
         .D(\registers[5] [5]), .Z(registers_5__1__N_1500)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__7__I_0_3_lut_4_lut (.A(n25380), .B(n25186), .C(debug_rd[3]), 
         .D(\registers[5] [7]), .Z(registers_5__3__N_1496)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_2__6__I_0_3_lut_4_lut (.A(n25185), .B(n25382), .C(debug_rd[2]), 
         .D(\registers[2] [6]), .Z(registers_2__2__N_1493)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__4__I_0_3_lut_4_lut (.A(n25185), .B(n25382), .C(debug_rd[0]), 
         .D(\registers[2] [4]), .Z(registers_2__0__N_1495)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__4__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__5__I_0_3_lut_4_lut (.A(n25185), .B(n25382), .C(debug_rd[1]), 
         .D(\registers[2] [5]), .Z(registers_2__1__N_1494)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__7__I_0_3_lut_4_lut (.A(n25185), .B(n25382), .C(debug_rd[3]), 
         .D(\registers[2] [7]), .Z(registers_2__3__N_1490)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__7__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__5__I_0_3_lut_4_lut (.A(n25186), .B(n25382), .C(debug_rd[1]), 
         .D(\registers[1] [5]), .Z(registers_1__1__N_1488)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__7__I_0_3_lut_4_lut (.A(n25186), .B(n25382), .C(debug_rd[3]), 
         .D(\registers[1] [7]), .Z(registers_1__3__N_1484)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__7__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__4__I_0_3_lut_4_lut (.A(n25186), .B(n25382), .C(debug_rd[0]), 
         .D(\registers[1] [4]), .Z(registers_1__0__N_1489)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__4__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__6__I_0_3_lut_4_lut (.A(n25186), .B(n25382), .C(debug_rd[2]), 
         .D(\registers[1] [6]), .Z(registers_1__2__N_1487)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11656_2_lut_rep_641 (.A(rd[2]), .B(rd[3]), .Z(n25377)) /* synthesis lut_function=(A (B)) */ ;
    defparam i11656_2_lut_rep_641.init = 16'h8888;
    LUT4 equal_134_i6_2_lut_rep_643 (.A(rd[2]), .B(rd[3]), .Z(n25379)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam equal_134_i6_2_lut_rep_643.init = 16'hbbbb;
    LUT4 i21219_3_lut (.A(\registers[2] [6]), .B(\reg_access[3][2] ), .C(rs2[0]), 
         .Z(n23494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21219_3_lut.init = 16'hcaca;
    LUT4 equal_129_i6_2_lut_rep_644 (.A(rd[2]), .B(rd[3]), .Z(n25380)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam equal_129_i6_2_lut_rep_644.init = 16'hdddd;
    LUT4 i12008_2_lut_rep_646 (.A(rd[3]), .B(rd[2]), .Z(n25382)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12008_2_lut_rep_646.init = 16'heeee;
    L6MUX21 i21185 (.D0(n23456), .D1(n23457), .SD(rs2[2]), .Z(n23460));
    LUT4 i21137_3_lut (.A(n23410), .B(n23411), .C(rs2[3]), .Z(data_rs2[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21137_3_lut.init = 16'hcaca;
    LUT4 i21292_4_lut_4_lut (.A(\registers[2] [7]), .B(rs2[0]), .C(rs2[1]), 
         .D(\registers[1] [7]), .Z(n23567)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i21292_4_lut_4_lut.init = 16'h2c20;
    L6MUX21 i21200 (.D0(n23471), .D1(n23472), .SD(rs1[2]), .Z(n23475));
    L6MUX21 i21215 (.D0(n23486), .D1(n23487), .SD(rs1[2]), .Z(n23490));
    L6MUX21 i21230 (.D0(n23501), .D1(n23502), .SD(rs2[2]), .Z(n23505));
    LUT4 i21344_3_lut_4_lut (.A(\registers[5] [5]), .B(rs2[0]), .C(rs2[1]), 
         .D(n5_adj_2343), .Z(n23407)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i21344_3_lut_4_lut.init = 16'hf808;
    LUT4 i21285_4_lut_4_lut (.A(\registers[2] [7]), .B(rs1[0]), .C(rs1[1]), 
         .D(\registers[1] [7]), .Z(n23560)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i21285_4_lut_4_lut.init = 16'h2c20;
    LUT4 i21138_4_lut_4_lut (.A(\registers[2] [5]), .B(rs1[0]), .C(rs1[1]), 
         .D(\registers[1] [5]), .Z(n23413)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i21138_4_lut_4_lut.init = 16'h2c20;
    LUT4 i21131_4_lut_4_lut (.A(\registers[2] [5]), .B(rs2[0]), .C(rs2[1]), 
         .D(\registers[1] [5]), .Z(n23406)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i21131_4_lut_4_lut.init = 16'h2c20;
    LUT4 i21341_3_lut_4_lut (.A(\registers[5] [5]), .B(rs1[0]), .C(rs1[1]), 
         .D(n5), .Z(n23414)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i21341_3_lut_4_lut.init = 16'hf808;
    LUT4 i21775_3_lut (.A(n26608), .B(n26610), .C(\counter_hi[2] ), .Z(\reg_access[4][3] )) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(40[41:55])
    defparam i21775_3_lut.init = 16'h0808;
    LUT4 mux_2187_i1_3_lut_4_lut_4_lut (.A(rd[0]), .B(\instr[12] ), .C(n25180), 
         .D(any_additional_mem_ops), .Z(n3645)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B+(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam mux_2187_i1_3_lut_4_lut_4_lut.init = 16'h5ccc;
    PFUMX i21135 (.BLUT(n23406), .ALUT(n23407), .C0(rs2[2]), .Z(n23410));
    L6MUX21 i21136 (.D0(n23408), .D1(n23409), .SD(rs2[2]), .Z(n23411));
    PFUMX i21142 (.BLUT(n23413), .ALUT(n23414), .C0(rs1[2]), .Z(n23417));
    L6MUX21 i21143 (.D0(n23415), .D1(n23416), .SD(rs1[2]), .Z(n23418));
    LUT4 i21298_3_lut (.A(n23571), .B(n23572), .C(rs2[3]), .Z(data_rs2[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21298_3_lut.init = 16'hcaca;
    PFUMX i21289 (.BLUT(n23560), .ALUT(n23561), .C0(rs1[2]), .Z(n23564));
    L6MUX21 i21186 (.D0(n23458), .D1(n23459), .SD(rs2[2]), .Z(n23461));
    L6MUX21 i21201 (.D0(n23473), .D1(n23474), .SD(rs1[2]), .Z(n23476));
    L6MUX21 i21216 (.D0(n23488), .D1(n23489), .SD(rs1[2]), .Z(n23491));
    L6MUX21 i21231 (.D0(n23503), .D1(n23504), .SD(rs2[2]), .Z(n23506));
    L6MUX21 i21290 (.D0(n23562), .D1(n23563), .SD(rs1[2]), .Z(n23565));
    L6MUX21 i21297 (.D0(n23569), .D1(n23570), .SD(rs2[2]), .Z(n23572));
    LUT4 i21291_3_lut (.A(n23564), .B(n23565), .C(rs1[3]), .Z(data_rs1[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21291_3_lut.init = 16'hcaca;
    PFUMX i21296 (.BLUT(n23567), .ALUT(n23568), .C0(rs2[2]), .Z(n23571));
    PFUMX i21133 (.BLUT(n8_adj_2342), .ALUT(n9_adj_2341), .C0(rs2[1]), 
          .Z(n23408));
    PFUMX i21134 (.BLUT(n11_adj_2340), .ALUT(n12_adj_2339), .C0(rs2[1]), 
          .Z(n23409));
    PFUMX i21140 (.BLUT(n8_adj_2338), .ALUT(n9_adj_2337), .C0(rs1[1]), 
          .Z(n23415));
    LUT4 i21218_3_lut (.A(\registers[1] [6]), .B(rs2[0]), .Z(n23493)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21218_3_lut.init = 16'h8888;
    PFUMX i21141 (.BLUT(n11_adj_2336), .ALUT(n12_adj_2335), .C0(rs1[1]), 
          .Z(n23416));
    LUT4 i21778_3_lut (.A(\counter_hi[2] ), .B(n26610), .C(n26608), .Z(\reg_access[3][2] )) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(38[47:61])
    defparam i21778_3_lut.init = 16'h0404;
    LUT4 i21204_3_lut (.A(\registers[2] [6]), .B(\reg_access[3][2] ), .C(rs1[0]), 
         .Z(n23479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21204_3_lut.init = 16'hcaca;
    LUT4 i21203_3_lut (.A(\registers[1] [6]), .B(rs1[0]), .Z(n23478)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21203_3_lut.init = 16'h8888;
    LUT4 i21189_3_lut (.A(\registers[2] [4]), .B(\reg_access[4][3] ), .C(rs1[0]), 
         .Z(n23464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21189_3_lut.init = 16'hcaca;
    LUT4 i21188_3_lut (.A(\registers[1] [4]), .B(rs1[0]), .Z(n23463)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21188_3_lut.init = 16'h8888;
    PFUMX i21182 (.BLUT(n23450), .ALUT(n23451), .C0(rs2[1]), .Z(n23457));
    PFUMX i21183 (.BLUT(n23452), .ALUT(n23453), .C0(rs2[1]), .Z(n23458));
    PFUMX i21184 (.BLUT(n23454), .ALUT(n23455), .C0(rs2[1]), .Z(n23459));
    PFUMX i21197 (.BLUT(n23465), .ALUT(n23466), .C0(rs1[1]), .Z(n23472));
    PFUMX i21198 (.BLUT(n23467), .ALUT(n23468), .C0(rs1[1]), .Z(n23473));
    PFUMX i21199 (.BLUT(n23469), .ALUT(n23470), .C0(rs1[1]), .Z(n23474));
    PFUMX i21212 (.BLUT(n23480), .ALUT(n23481), .C0(rs1[1]), .Z(n23487));
    LUT4 i21174_3_lut (.A(\registers[2] [4]), .B(\reg_access[4][3] ), .C(rs2[0]), 
         .Z(n23449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21174_3_lut.init = 16'hcaca;
    LUT4 i21173_3_lut (.A(\registers[1] [4]), .B(rs2[0]), .Z(n23448)) /* synthesis lut_function=(A (B)) */ ;
    defparam i21173_3_lut.init = 16'h8888;
    PFUMX i21213 (.BLUT(n23482), .ALUT(n23483), .C0(rs1[1]), .Z(n23488));
    PFUMX i21214 (.BLUT(n23484), .ALUT(n23485), .C0(rs1[1]), .Z(n23489));
    PFUMX i21227 (.BLUT(n23495), .ALUT(n23496), .C0(rs2[1]), .Z(n23502));
    PFUMX i21228 (.BLUT(n23497), .ALUT(n23498), .C0(rs2[1]), .Z(n23503));
    PFUMX i21229 (.BLUT(n23499), .ALUT(n23500), .C0(rs2[1]), .Z(n23504));
    PFUMX i21287 (.BLUT(n8_adj_2334), .ALUT(n9_adj_2333), .C0(rs1[1]), 
          .Z(n23562));
    PFUMX i21288 (.BLUT(n11_adj_2332), .ALUT(n12_adj_2331), .C0(rs1[1]), 
          .Z(n23563));
    PFUMX i21294 (.BLUT(n8), .ALUT(n9), .C0(rs2[1]), .Z(n23569));
    PFUMX i21295 (.BLUT(n11), .ALUT(n12), .C0(rs2[1]), .Z(n23570));
    
endmodule
//
// Verilog Description of module tinyqv_counter_U0
//

module tinyqv_counter_U0 (cy, clk_c, n25424, \increment_result_3__N_1656[0] , 
            instrret_count, n25294, n25308) /* synthesis syn_module_defined=1 */ ;
    output cy;
    input clk_c;
    input n25424;
    input \increment_result_3__N_1656[0] ;
    output [3:0]instrret_count;
    input n25294;
    input n25308;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [4:0]increment_result_3__N_1656;
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    
    FD1S3IX cy_51 (.D(increment_result_3__N_1656[4]), .CK(clk_c), .CD(n25424), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3IX register_2__48 (.D(increment_result_3__N_1656[2]), .CK(clk_c), 
            .CD(n25424), .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result_3__N_1656[1]), .CK(clk_c), 
            .CD(n25424), .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(\increment_result_3__N_1656[0] ), .CK(clk_c), 
            .CD(n25424), .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(register[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(register[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(register[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(instrret_count[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(register[10]), .CK(clk_c), .Q(instrret_count[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(register[9]), .CK(clk_c), .Q(instrret_count[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(register[8]), .CK(clk_c), .Q(instrret_count[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result_3__N_1656[3]), .CK(clk_c), 
            .CD(n25424), .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 i3968_2_lut_3_lut_4_lut (.A(instrret_count[1]), .B(n25294), .C(instrret_count[3]), 
         .D(instrret_count[2]), .Z(increment_result_3__N_1656[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i3968_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i3970_2_lut_3_lut_4_lut (.A(instrret_count[1]), .B(n25294), .C(instrret_count[3]), 
         .D(instrret_count[2]), .Z(increment_result_3__N_1656[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i3970_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i3954_2_lut_3_lut (.A(instrret_count[0]), .B(n25308), .C(instrret_count[1]), 
         .Z(increment_result_3__N_1656[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i3954_2_lut_3_lut.init = 16'h7878;
    LUT4 i3961_2_lut_3_lut_4_lut (.A(instrret_count[0]), .B(n25308), .C(instrret_count[2]), 
         .D(instrret_count[1]), .Z(increment_result_3__N_1656[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i3961_2_lut_3_lut_4_lut.init = 16'h78f0;
    
endmodule
//
// Verilog Description of module \tinyqv_counter(OUTPUT_WIDTH=7) 
//

module \tinyqv_counter(OUTPUT_WIDTH=7)  (cy, clk_c, n25424, \increment_result_3__N_1642[1] , 
            \increment_result_3__N_1642[0] , cycle_count_wide, n25298, 
            n25315, n25246) /* synthesis syn_module_defined=1 */ ;
    output cy;
    input clk_c;
    input n25424;
    input \increment_result_3__N_1642[1] ;
    input \increment_result_3__N_1642[0] ;
    output [6:0]cycle_count_wide;
    input n25298;
    input n25315;
    output n25246;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [4:0]increment_result_3__N_1642;
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    
    FD1S3IX cy_51 (.D(increment_result_3__N_1642[4]), .CK(clk_c), .CD(n25424), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3IX register_2__48 (.D(increment_result_3__N_1642[2]), .CK(clk_c), 
            .CD(n25424), .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(\increment_result_3__N_1642[1] ), .CK(clk_c), 
            .CD(n25424), .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(\increment_result_3__N_1642[0] ), .CK(clk_c), 
            .CD(n25424), .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(cycle_count_wide[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(cycle_count_wide[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(cycle_count_wide[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(cycle_count_wide[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(cycle_count_wide[6]), .CK(clk_c), .Q(cycle_count_wide[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(cycle_count_wide[5]), .CK(clk_c), .Q(cycle_count_wide[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(cycle_count_wide[4]), .CK(clk_c), .Q(cycle_count_wide[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result_3__N_1642[3]), .CK(clk_c), 
            .CD(n25424), .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 i3942_2_lut_3_lut_4_lut (.A(cycle_count_wide[1]), .B(n25298), .C(cycle_count_wide[3]), 
         .D(cycle_count_wide[2]), .Z(increment_result_3__N_1642[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i3942_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i3940_2_lut_3_lut_4_lut (.A(cycle_count_wide[1]), .B(n25298), .C(cycle_count_wide[3]), 
         .D(cycle_count_wide[2]), .Z(increment_result_3__N_1642[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i3940_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i3935_2_lut_rep_510_3_lut_4_lut (.A(cycle_count_wide[0]), .B(n25315), 
         .C(cycle_count_wide[2]), .D(cycle_count_wide[1]), .Z(n25246)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i3935_2_lut_rep_510_3_lut_4_lut.init = 16'h8000;
    LUT4 i3933_2_lut_3_lut_4_lut (.A(cycle_count_wide[0]), .B(n25315), .C(cycle_count_wide[2]), 
         .D(cycle_count_wide[1]), .Z(increment_result_3__N_1642[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i3933_2_lut_3_lut_4_lut.init = 16'h78f0;
    
endmodule
//
// Verilog Description of module tinyqv_alu
//

module tinyqv_alu (n22558, \alu_op_in[2] , n25254, alu_a_in, n25218, 
            n25274, alu_b_in, n21812, n25251, cy_out, n24569, n25250, 
            n25352, n25318, n25357, n24571, n4411, n25358, alu_out) /* synthesis syn_module_defined=1 */ ;
    input n22558;
    input \alu_op_in[2] ;
    input n25254;
    input [3:0]alu_a_in;
    input n25218;
    input n25274;
    input [3:0]alu_b_in;
    input n21812;
    input n25251;
    output cy_out;
    output n24569;
    input n25250;
    input n25352;
    input n25318;
    input n25357;
    output n24571;
    input [3:0]n4411;
    input n25358;
    output [3:0]alu_out;
    
    wire [3:0]a_xor_b;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[16:23])
    wire [3:0]n4421;
    
    wire n22498, n25285, n25200, n25217, n26595, n22464, n25188, 
        n22442, n6, cmp_res_N_1586, n25187, n26594, n24570, n25192;
    wire [3:0]n4430;
    
    LUT4 mux_2677_i1_4_lut (.A(n22558), .B(a_xor_b[0]), .C(\alu_op_in[2] ), 
         .D(n25254), .Z(n4421[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_2677_i1_4_lut.init = 16'hc5ca;
    LUT4 mux_2677_i2_4_lut (.A(n22498), .B(n25285), .C(\alu_op_in[2] ), 
         .D(n25200), .Z(n4421[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_2677_i2_4_lut.init = 16'hc5ca;
    LUT4 i4611_4_lut_rep_703 (.A(alu_a_in[1]), .B(n25218), .C(n25217), 
         .D(n25274), .Z(n26595)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4611_4_lut_rep_703.init = 16'haaa8;
    LUT4 mux_2677_i3_4_lut (.A(n22464), .B(a_xor_b[2]), .C(\alu_op_in[2] ), 
         .D(n25188), .Z(n4421[2])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_2677_i3_4_lut.init = 16'hc5ca;
    LUT4 a_3__I_0_29_i3_2_lut (.A(alu_a_in[2]), .B(alu_b_in[2]), .Z(a_xor_b[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i3_2_lut.init = 16'h6666;
    LUT4 a_3__I_0_29_i4_2_lut (.A(alu_a_in[3]), .B(alu_b_in[3]), .Z(a_xor_b[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i4_2_lut.init = 16'h6666;
    LUT4 a_3__I_0_29_i1_2_lut (.A(alu_a_in[0]), .B(alu_b_in[0]), .Z(a_xor_b[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i1_2_lut.init = 16'h6666;
    LUT4 mux_2677_i4_4_lut (.A(n22442), .B(a_xor_b[3]), .C(\alu_op_in[2] ), 
         .D(n6), .Z(n4421[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_2677_i4_4_lut.init = 16'hc5ca;
    LUT4 i1_4_lut (.A(a_xor_b[2]), .B(a_xor_b[3]), .C(a_xor_b[0]), .D(n21812), 
         .Z(cmp_res_N_1586)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    LUT4 i3882_2_lut_rep_452_3_lut_4_lut_4_lut (.A(alu_a_in[1]), .B(n25218), 
         .C(n25217), .D(n25274), .Z(n25188)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i3882_2_lut_rep_452_3_lut_4_lut_4_lut.init = 16'hfea8;
    LUT4 i3896_4_lut_4_lut (.A(alu_a_in[3]), .B(n25187), .C(n26594), .D(n25251), 
         .Z(cy_out)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i3896_4_lut_4_lut.init = 16'hfea8;
    LUT4 alu_op_in_0__bdd_4_lut (.A(n25187), .B(n26594), .C(n25251), .D(alu_a_in[3]), 
         .Z(n24569)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C (D))))) */ ;
    defparam alu_op_in_0__bdd_4_lut.init = 16'h011f;
    LUT4 n5915_bdd_4_lut (.A(n25187), .B(n26594), .C(n25251), .D(alu_a_in[3]), 
         .Z(n24570)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+(D)))) */ ;
    defparam n5915_bdd_4_lut.init = 16'hf110;
    LUT4 i4590_rep_702 (.A(alu_a_in[2]), .B(n26595), .C(n25192), .D(n25250), 
         .Z(n26594)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4590_rep_702.init = 16'haaa8;
    LUT4 i1_2_lut_3_lut (.A(alu_b_in[2]), .B(n25352), .C(alu_a_in[2]), 
         .Z(n22464)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_adj_203 (.A(alu_b_in[3]), .B(n25352), .C(alu_a_in[3]), 
         .Z(n22442)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut_adj_203.init = 16'h9696;
    LUT4 i4612_3_lut_rep_481_4_lut (.A(alu_b_in[0]), .B(n25352), .C(n25318), 
         .D(alu_a_in[0]), .Z(n25217)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i4612_3_lut_rep_481_4_lut.init = 16'hf600;
    LUT4 i3887_2_lut_rep_451_3_lut_4_lut (.A(n25274), .B(n25200), .C(n25250), 
         .D(n26595), .Z(n25187)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i3887_2_lut_rep_451_3_lut_4_lut.init = 16'hf080;
    LUT4 i3875_2_lut_rep_464_4_lut_3_lut_4_lut (.A(alu_b_in[0]), .B(n25352), 
         .C(alu_a_in[0]), .D(n25318), .Z(n25200)) /* synthesis lut_function=(A (B (C (D))+!B (C+(D)))+!A (B (C+(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i3875_2_lut_rep_464_4_lut_3_lut_4_lut.init = 16'hf660;
    PFUMX i22178 (.BLUT(cmp_res_N_1586), .ALUT(n24570), .C0(n25357), .Z(n24571));
    LUT4 i3889_2_lut_3_lut_4_lut_4_lut (.A(alu_a_in[2]), .B(n26595), .C(n25192), 
         .D(n25250), .Z(n6)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i3889_2_lut_3_lut_4_lut_4_lut.init = 16'hfea8;
    PFUMX mux_2682_i4 (.BLUT(n4421[3]), .ALUT(n4411[3]), .C0(n25357), 
          .Z(n4430[3]));
    PFUMX mux_2682_i3 (.BLUT(n4421[2]), .ALUT(n4411[2]), .C0(n25357), 
          .Z(n4430[2]));
    LUT4 i1_2_lut_3_lut_adj_204 (.A(alu_b_in[1]), .B(n25352), .C(alu_a_in[1]), 
         .Z(n22498)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut_adj_204.init = 16'h9696;
    PFUMX mux_2682_i2 (.BLUT(n4421[1]), .ALUT(n4411[1]), .C0(n25357), 
          .Z(n4430[1]));
    LUT4 i11994_2_lut_4_lut (.A(n25358), .B(\alu_op_in[2] ), .C(n25357), 
         .D(n4430[1]), .Z(alu_out[1])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i11994_2_lut_4_lut.init = 16'hc500;
    LUT4 i11768_2_lut_4_lut (.A(n25358), .B(\alu_op_in[2] ), .C(n25357), 
         .D(n4430[0]), .Z(alu_out[0])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i11768_2_lut_4_lut.init = 16'hc500;
    LUT4 i11996_2_lut_4_lut (.A(n25358), .B(\alu_op_in[2] ), .C(n25357), 
         .D(n4430[3]), .Z(alu_out[3])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i11996_2_lut_4_lut.init = 16'hc500;
    LUT4 i11995_2_lut_4_lut (.A(n25358), .B(\alu_op_in[2] ), .C(n25357), 
         .D(n4430[2]), .Z(alu_out[2])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i11995_2_lut_4_lut.init = 16'hc500;
    PFUMX mux_2682_i1 (.BLUT(n4421[0]), .ALUT(n4411[0]), .C0(n25357), 
          .Z(n4430[0]));
    LUT4 a_3__I_0_29_i2_2_lut_rep_549 (.A(alu_a_in[1]), .B(alu_b_in[1]), 
         .Z(n25285)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i2_2_lut_rep_549.init = 16'h6666;
    LUT4 i3880_2_lut_rep_456_3_lut_4_lut (.A(n25254), .B(n25318), .C(n25274), 
         .D(n25217), .Z(n25192)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i3880_2_lut_rep_456_3_lut_4_lut.init = 16'hf080;
    
endmodule
