// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Thu Jan 08 21:50:47 2026
//
// Verilog Description of module tinyQV_top
//

module tinyQV_top (clk, rst_n, ui_in, uo_out) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(8[8:18])
    input clk;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    input rst_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(10[20:25])
    input [7:0]ui_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    output [7:0]uo_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    wire GND_net, VCC_net, rst_n_c, ui_in_c_7, ui_in_c_6, ui_in_c_5, 
        ui_in_c_4, ui_in_c_3, ui_in_c_2, ui_in_c_1, ui_in_c_0, uo_out_c_7, 
        uo_out_c_6, uo_out_c_5, uo_out_c_4, uo_out_c_3, uo_out_c_2, 
        uo_out_c_1, uo_out_c_0, rst_reg_n;
    wire [3:0]qspi_data_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(34[16:28])
    
    wire n31717;
    wire [3:0]qspi_data_oe;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(36[16:28])
    
    wire qspi_ram_a_select, qspi_ram_b_select;
    wire [27:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    wire [31:0]data_to_write;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(56[17:30])
    wire [31:0]data_from_read;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(59[16:30])
    wire [3:0]debug_rd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(75[16:24])
    
    wire debug_uart_txd;
    wire [7:6]gpio_out_sel;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(79[16:28])
    
    wire debug_register_data;
    wire [3:0]debug_rd_r;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(85[15:25])
    
    wire debug_uart_tx_start;
    wire [7:0]peri_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(95[16:24])
    
    wire n23720;
    wire [31:0]peri_data_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(96[17:30])
    wire [7:0]ui_in_sync0;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(101[15:26])
    wire [7:0]ui_in_sync;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(102[15:25])
    wire [7:0]time_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(238[15:25])
    wire [3:0]qspi_data_in_3__N_1;
    wire [3:0]qspi_data_out_3__N_5;
    wire [1:0]gpio_out_sel_7__N_13;
    wire [24:0]addr_adj_3335;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(23[16:20])
    
    wire n51;
    wire [31:0]addr_24__N_228;
    wire [31:0]writing_N_164;
    
    wire debug_instr_valid, debug_stop_txn;
    wire [23:1]instr_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(56[15:25])
    wire [15:0]instr_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(61[15:25])
    
    wire rst_reg_n_adj_3274, data_out_hold, data_ready_r, n29752, n29751, 
        n29201, n51_adj_3275, n54, n29750, n29749, n29747, n29199, 
        n41, n40, n15604, n27030, clk_c_enable_186, clk_c_enable_324, 
        clk_c_enable_452, n84, n39, n38, n26266, clk_c_enable_395, 
        n23719, n23718, n23717, n23653, n23716;
    wire [7:0]\uo_out_from_user_peri[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(59[17:38])
    wire [7:0]\uo_out_from_user_peri[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(59[17:38])
    wire [12:0]baud_divider_adj_3392;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(36[31:43])
    
    wire n23715, n60, n48, n23652, n23714, n23651, n31819, n23713, 
        n4263, n45, n63, n33, n29198, n33_adj_3276, n23712, n23711;
    wire [4:0]\gpio_out_func_sel[0] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    wire [4:0]\gpio_out_func_sel[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    wire [4:0]\gpio_out_func_sel[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    wire [4:0]\gpio_out_func_sel[3] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    wire [4:0]\gpio_out_func_sel[4] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    wire [4:0]\gpio_out_func_sel[5] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    wire [4:0]\gpio_out_func_sel[6] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    wire [4:0]\gpio_out_func_sel[7] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    
    wire led_out, data_ready_r_N_2792, n39_adj_3277, n23650, n8819, 
        n6228, n6232, n42, n23710, n23709;
    wire [12:0]cycle_counter;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(43[25:38])
    wire [3:0]fsm_state;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(47[11:20])
    
    wire next_bit, n23649, uart_txd_N_2974, n26036, is_ret_de;
    wire [31:0]imm;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(100[16:19])
    wire [2:1]instr_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(113[15:24])
    wire [3:0]rs1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(117[15:18])
    wire [3:0]rs2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(118[15:18])
    wire [3:0]rd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(119[15:17])
    wire [31:0]pc;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(128[17:19])
    wire [31:0]next_pc_for_core;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(129[17:33])
    wire [4:2]counter_hi;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(139[15:25])
    wire [3:1]instr_write_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(152[15:33])
    
    wire was_early_branch;
    wire [3:0]data_out_slice;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(230[16:30])
    wire [15:0]\instr_data[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]\instr_data[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]\instr_data[3] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [23:1]early_branch_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[17:34])
    
    wire n4, n31064, n10500, n31063, n31062, n31061, n31742, n31060, 
        n57, n10499, n31059, n42_adj_3278, n30, n8, clk_c_enable_360, 
        n8135, n80, n23648, clk_c_enable_349;
    wire [59:0]debug_rd_3__N_405;
    
    wire clk_c_enable_259, n23647, n26116, n23705, n10573, n42_adj_3279, 
        n23704;
    wire [22:0]instr_addr_23__N_318;
    
    wire clk_c_enable_357, n1724, n57_adj_3280, data_stall, instr_active_N_2106, 
        n23703, n29633, clk_c_enable_273, n28276, n7884, n23702, 
        continue_txn_N_2131, data_stall_N_2158, n31798, n23701, n23700, 
        n23699, n23698, n23697, n28246, n23696, n23646, n28242, 
        n23695, n23694, n31716, n54_adj_3281, n45_adj_3282, clk_c_enable_387, 
        n28230, n2524, n2514, n2152, n2136, n23645, n23693, n2565, 
        clk_c_enable_231, n23692, n18086, n23690, n2208, n23689, 
        n2504;
    wire [1:0]cycle;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(58[15:20])
    wire [3:0]alu_b_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[16:24])
    wire [3:0]mul_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(138[16:23])
    
    wire n23688, alu_b_in_3__N_1504, n31735, instr_complete_N_1647, 
        n23687, clk_c_enable_234, n66, n44, n43, n23686, n9, n23685, 
        data_out_3__N_1385, clk_c_enable_542, n39_adj_3283, n23684, 
        n23683, n23682, n23681, n60_adj_3284, n31713, n28964, n23633, 
        n32077;
    wire [3:0]csr_read_3__N_1447;
    
    wire clk_c_enable_376, n66_adj_3285, n23632, n23634, n63_adj_3286, 
        n32055, n27620, n30906, n3, n30905, n30904, clk_c_enable_239, 
        clk_c_enable_445, n32035, n32034, n32033, n5171, n27183, 
        n32031, n32027, n27421, n29162, n32022, n32021, n18241, 
        n23670, n23669, n32019;
    wire [2:0]fsm_state_adj_3443;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(82[15:24])
    
    wire is_writing;
    wire [23:0]addr_adj_3444;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(84[31:35])
    wire [2:0]nibbles_remaining;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(86[15:32])
    
    wire stop_txn_reg, stop_txn_now_N_2363, n32017, is_writing_N_2331, 
        n32016, n32013, n10467, n23637, n23668, n32003, n31593, 
        n48_adj_3288, n6210, n31997, clk_c_enable_531, n30_adj_3289, 
        clk_c_enable_534, n4_adj_3290, n1084, n45_adj_3291, n36, n28850;
    wire [12:0]cycle_counter_adj_3465;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(43[25:38])
    wire [3:0]fsm_state_adj_3466;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(47[11:20])
    
    wire next_bit_adj_3308, n26282, n23667, n28840, n26205, n31978, 
        n31977, n12, n23666, n23665, clk_c_enable_36;
    wire [12:0]cycle_counter_adj_3488;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(39[25:38])
    wire [3:0]fsm_state_adj_3489;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(47[11:20])
    
    wire next_bit_adj_3326, n23664, n31971;
    wire [31:0]next_fsm_state_3__N_3015;
    
    wire n23635, n11, n23663, n23636, n23662, n23631, n23661, 
        n1160, n31967, n23660;
    wire [31:0]\registers[5] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[6] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[7] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n36_adj_3327, n31964, n31963, n31962, n31961;
    wire [15:0]accum;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(104[22:27])
    wire [19:0]next_accum;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[23:33])
    wire [19:0]d_3__N_1868;
    
    wire n31958, n23659, n23658, n23657, n23732, n23731, n1, n31950, 
        n23730, n28800, n23729, n780, n31944, n33479, n23656, 
        n26216, n23728, n23727, n28760, n31936, n23725, n31935, 
        n31934, clk_c_enable_268, n31932, n24, n23724, n23723, n23722, 
        n31389, n31388, n31930, n31929, n9_adj_3328, n8_adj_3329, 
        n31927, n23721, n31925, n27081, n31923, n31922, n31761, 
        n31906, n31905, n31904, n28686, n31902, n31901, n28950, 
        n31900, n28626, n28624, n31885, n19, n4_adj_3330, n31883, 
        n31880, n31879, n32105, n32104, n14, n32103, n28966, n14_adj_3331, 
        n28968, n32101, n32100, n32088, n29004, n10, n32087, n31869, 
        n31868, n31867, n28538, n3_adj_3332, n31865, n31864, n31863, 
        n31712, n27464, n27347, n31860, clk_c_enable_390, n31855, 
        clk_c_enable_355, n31853, n31849, n31847, n31844, n31164, 
        n31163, n31841, n31162, n31828;
    
    VHI i2 (.Z(VCC_net));
    INV i29333 (.A(clk_c), .Z(clk_N_45));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    FD1S3AX debug_rd_r_i0 (.D(debug_rd[0]), .CK(clk_c), .Q(debug_rd_r[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(257[12] 259[8])
    defparam debug_rd_r_i0.GSR = "DISABLED";
    FD1S3AX rst_reg_n_53 (.D(rst_n_c), .CK(clk_N_45), .Q(rst_reg_n));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(31[12:46])
    defparam rst_reg_n_53.GSR = "DISABLED";
    CCU2C _add_1_5116_add_4_5 (.A0(early_branch_addr[5]), .B0(was_early_branch), 
          .C0(pc[5]), .D0(VCC_net), .A1(early_branch_addr[6]), .B1(was_early_branch), 
          .C1(pc[6]), .D1(VCC_net), .CIN(n23710), .COUT(n23711), .S0(instr_addr_23__N_318[4]), 
          .S1(instr_addr_23__N_318[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_5.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_5.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_10 (.A0(accum[8]), .B0(d_3__N_1868[8]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[9]), .B1(d_3__N_1868[9]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23648), .COUT(n23649), .S0(next_accum[8]), 
          .S1(next_accum[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_5116_add_4_3 (.A0(pc[3]), .B0(was_early_branch), .C0(early_branch_addr[3]), 
          .D0(instr_write_offset[3]), .A1(early_branch_addr[4]), .B1(was_early_branch), 
          .C1(pc[4]), .D1(VCC_net), .CIN(n23709), .COUT(n23710), .S0(instr_addr_23__N_318[2]), 
          .S1(instr_addr_23__N_318[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_3.INIT0 = 16'hd1e2;
    defparam _add_1_5116_add_4_3.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5116_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(was_early_branch), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n23709));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5116_add_4_1.INIT1 = 16'hffff;
    defparam _add_1_5116_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_5127_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23705), .S0(next_bit_adj_3308));
    defparam _add_1_5127_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_5127_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_5127_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_5127_add_4_cout.INJECT1_1 = "NO";
    \peripherals_min(CLOCK_MHZ=14)  i_peripherals (.\peri_data_out[4] (peri_data_out[4]), 
            .clk_c(clk_c), .clk_c_enable_387(clk_c_enable_387), .\peri_data_out[3] (peri_data_out[3]), 
            .\peri_data_out[0] (peri_data_out[0]), .\peri_data_out[2] (peri_data_out[2]), 
            .\peri_data_out[1] (peri_data_out[1]), .\gpio_out_func_sel[5] ({\gpio_out_func_sel[5] }), 
            .clk_c_enable_445(clk_c_enable_445), .\data_to_write[2] (data_to_write[2]), 
            .clk_c_enable_349(clk_c_enable_349), .\data_to_write[4] (data_to_write[4]), 
            .data_out_hold(data_out_hold), .n31883(n31883), .clk_c_enable_360(clk_c_enable_360), 
            .\data_to_write[3] (data_to_write[3]), .\gpio_out_func_sel[3] ({Open_0, 
            \gpio_out_func_sel[3] [3], Open_1, Open_2, Open_3}), .clk_c_enable_357(clk_c_enable_357), 
            .clk_c_enable_259(clk_c_enable_259), .\data_to_write[1] (data_to_write[1]), 
            .clk_c_enable_273(clk_c_enable_273), .\gpio_out_func_sel[7][3] (\gpio_out_func_sel[7] [3]), 
            .n32035(n32035), .n26282(n26282), .\addr[6] (addr[6]), .\addr[9] (addr[9]), 
            .n31934(n31934), .n32034(n32034), .ui_in_sync({ui_in_sync}), 
            .n32019(n32019), .\gpio_out_func_sel[1][3] (\gpio_out_func_sel[1] [3]), 
            .\data_to_write[0] (data_to_write[0]), .\addr[2] (addr[2]), 
            .\addr[3] (addr[3]), .\gpio_out_func_sel[4][3] (\gpio_out_func_sel[4] [3]), 
            .\gpio_out_func_sel[7][4] (\gpio_out_func_sel[7] [4]), .\gpio_out_func_sel[7][2] (\gpio_out_func_sel[7] [2]), 
            .baud_divider({baud_divider_adj_3392}), .n31922(n31922), .\gpio_out_func_sel[2][3] (\gpio_out_func_sel[2] [3]), 
            .\uo_out_from_user_peri[1][5] (\uo_out_from_user_peri[1] [5]), 
            .n32003(n32003), .n26205(n26205), .\gpio_out_func_sel[6][3] (\gpio_out_func_sel[6] [3]), 
            .\gpio_out_func_sel[0][3] (\gpio_out_func_sel[0] [3]), .data_ready_r(data_ready_r), 
            .rst_reg_n(rst_reg_n), .data_ready_r_N_2792(data_ready_r_N_2792), 
            .\peri_data_out[12] (peri_data_out[12]), .\peri_data_out[11] (peri_data_out[11]), 
            .\peri_data_out[10] (peri_data_out[10]), .\peri_data_out[9] (peri_data_out[9]), 
            .\peri_data_out[8] (peri_data_out[8]), .\peri_data_out[7] (peri_data_out[7]), 
            .\peri_data_out[6] (peri_data_out[6]), .\peri_data_out[5] (peri_data_out[5]), 
            .led_out(led_out), .\addr[10] (addr[10]), .\addr[4] (addr[4]), 
            .\addr[8] (addr[8]), .n4(n4_adj_3290), .n28840(n28840), .\uo_out_from_user_peri[1][3] (\uo_out_from_user_peri[1] [3]), 
            .\data_to_write[5] (data_to_write[5]), .\data_to_write[6] (data_to_write[6]), 
            .\data_to_write[7] (data_to_write[7]), .\addr[7] (addr[7]), 
            .n31967(n31967), .n32017(n32017), .n8819(n8819), .n31962(n31962), 
            .n31935(n31935), .n18241(n18241), .n31936(n31936), .\debug_rd_r[0] (debug_rd_r[0]), 
            .debug_register_data(debug_register_data), .uo_out_c_2(uo_out_c_2), 
            .\debug_rd_r[1] (debug_rd_r[1]), .uo_out_c_3(uo_out_c_3), .\uo_out_from_user_peri[2][7] (\uo_out_from_user_peri[2] [7]), 
            .n26266(n26266), .clk_c_enable_268(clk_c_enable_268), .n31901(n31901), 
            .n80(n80), .n31900(n31900), .n1(n1), .\debug_rd_r[2] (debug_rd_r[2]), 
            .uo_out_c_4(uo_out_c_4), .\peri_out[6] (peri_out[6]), .n3(n3), 
            .uo_out_c_0(uo_out_c_0), .uo_out_c_1(uo_out_c_1), .clk_c_enable_542(clk_c_enable_542), 
            .clk_c_enable_390(clk_c_enable_390), .clk_c_enable_395(clk_c_enable_395), 
            .\data_to_write[8] (data_to_write[8]), .\data_to_write[9] (data_to_write[9]), 
            .\data_to_write[10] (data_to_write[10]), .\data_to_write[11] (data_to_write[11]), 
            .\data_to_write[12] (data_to_write[12]), .\next_fsm_state_3__N_3015[3] (next_fsm_state_3__N_3015[3]), 
            .n27347(n27347), .n31932(n31932), .n26116(n26116), .n26216(n26216), 
            .n31905(n31905), .n32033(n32033), .n31929(n31929), .\imm[6] (imm[6]), 
            .\csr_read_3__N_1447[2] (csr_read_3__N_1447[2]), .n29162(n29162), 
            .cycle_counter({cycle_counter_adj_3465}), .n72({n30, n33, 
            n36_adj_3327, n39_adj_3283, n42_adj_3279, n45, n48, n51, 
            n54_adj_3281, n57_adj_3280, n60, n63_adj_3286, n66}), 
            .fsm_state({fsm_state_adj_3466}), .n31855(n31855), .next_bit(next_bit_adj_3308), 
            .n31963(n31963), .fsm_state_adj_72({fsm_state_adj_3489}), .next_bit_adj_56(next_bit_adj_3326), 
            .cycle_counter_adj_73({cycle_counter_adj_3488}), .n28760(n28760), 
            .GND_net(GND_net), .VCC_net(VCC_net), .n31902(n31902), .n31925(n31925), 
            .n31923(n31923), .next_bit_adj_70(next_bit), .n31828(n31828), 
            .uart_txd_N_2974(uart_txd_N_2974), .clk_c_enable_534(clk_c_enable_534), 
            .debug_stop_txn(debug_stop_txn), .instr_active_N_2106(instr_active_N_2106), 
            .n32013(n32013), .\fsm_state[0]_adj_71 (fsm_state[0]), .clk_c_enable_376(clk_c_enable_376), 
            .n28686(n28686), .n31880(n31880), .clk_c_enable_355(clk_c_enable_355), 
            .n1084(n1084), .stop_txn_reg(stop_txn_reg), .stop_txn_now_N_2363(stop_txn_now_N_2363), 
            .clk_c_enable_239(clk_c_enable_239), .n31971(n31971), .n33479(n33479), 
            .\qspi_data_in[1] (qspi_data_in[1]), .n31593(n31593), .n31927(n31927), 
            .n27620(n27620), .n31906(n31906), .n27081(n27081), .n6210(n6210), 
            .n31819(n31819), .n28800(n28800), .n32027(n32027), .clk_c_enable_531(clk_c_enable_531), 
            .n31950(n31950), .n31977(n31977), .n8135(n8135), .n10499(n10499), 
            .n10500(n10500), .clk_c_enable_186(clk_c_enable_186), .n32021(n32021), 
            .n31997(n31997), .\addr[27] (addr[27]), .n31930(n31930), .n32022(n32022), 
            .n31958(n31958), .n26036(n26036), .instr_complete_N_1647(instr_complete_N_1647), 
            .n28276(n28276), .n31717(n31717), .n29201(n29201)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(161[46] 180[6])
    CCU2C _add_1_add_4_add_4_8 (.A0(accum[6]), .B0(d_3__N_1868[6]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[7]), .B1(d_3__N_1868[7]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23647), .COUT(n23648), .S0(next_accum[6]), 
          .S1(next_accum[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_5127_add_4_14 (.A0(baud_divider_adj_3392[11]), .B0(cycle_counter_adj_3465[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[12]), 
          .B1(cycle_counter_adj_3465[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23704), .COUT(n23705));
    defparam _add_1_5127_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_5127_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_5127_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_5127_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_5127_add_4_12 (.A0(baud_divider_adj_3392[9]), .B0(cycle_counter_adj_3465[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[10]), 
          .B1(cycle_counter_adj_3465[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23703), .COUT(n23704));
    defparam _add_1_5127_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_5127_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_5127_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_5127_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_5127_add_4_10 (.A0(baud_divider_adj_3392[7]), .B0(cycle_counter_adj_3465[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[8]), .B1(cycle_counter_adj_3465[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23702), .COUT(n23703));
    defparam _add_1_5127_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_5127_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_5127_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_5127_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_5127_add_4_8 (.A0(baud_divider_adj_3392[5]), .B0(cycle_counter_adj_3465[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[6]), .B1(cycle_counter_adj_3465[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23701), .COUT(n23702));
    defparam _add_1_5127_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_5127_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_5127_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_5127_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_5127_add_4_6 (.A0(baud_divider_adj_3392[3]), .B0(cycle_counter_adj_3465[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[4]), .B1(cycle_counter_adj_3465[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23700), .COUT(n23701));
    defparam _add_1_5127_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_5127_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_5127_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_5127_add_4_6.INJECT1_1 = "NO";
    LUT4 i27755_2_lut (.A(n10573), .B(rst_reg_n), .Z(n780)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i27755_2_lut.init = 16'h7777;
    CCU2C _add_1_5127_add_4_4 (.A0(baud_divider_adj_3392[1]), .B0(cycle_counter_adj_3465[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[2]), .B1(cycle_counter_adj_3465[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23699), .COUT(n23700));
    defparam _add_1_5127_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_5127_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_5127_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_5127_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_5127_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(baud_divider_adj_3392[0]), .B1(cycle_counter_adj_3465[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n23699));
    defparam _add_1_5127_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_5127_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_5127_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_5127_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_5119_add_4_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23698), .S0(next_bit_adj_3326));
    defparam _add_1_5119_add_4_cout.INIT0 = 16'h0000;
    defparam _add_1_5119_add_4_cout.INIT1 = 16'h0000;
    defparam _add_1_5119_add_4_cout.INJECT1_0 = "NO";
    defparam _add_1_5119_add_4_cout.INJECT1_1 = "NO";
    CCU2C _add_1_5119_add_4_14 (.A0(baud_divider_adj_3392[11]), .B0(cycle_counter_adj_3488[11]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[12]), 
          .B1(cycle_counter_adj_3488[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23697), .COUT(n23698));
    defparam _add_1_5119_add_4_14.INIT0 = 16'h9995;
    defparam _add_1_5119_add_4_14.INIT1 = 16'h9995;
    defparam _add_1_5119_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_5119_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_6 (.A0(accum[4]), .B0(d_3__N_1868[4]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[5]), .B1(d_3__N_1868[5]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23646), .COUT(n23647), .S0(next_accum[4]), 
          .S1(next_accum[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_4 (.A0(accum[2]), .B0(d_3__N_1868[2]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[3]), .B1(d_3__N_1868[3]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23645), .COUT(n23646), .S0(mul_out[2]), 
          .S1(mul_out[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_2 (.A0(accum[0]), .B0(d_3__N_1868[0]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[1]), .B1(d_3__N_1868[1]), .C1(GND_net), 
          .D1(VCC_net), .COUT(n23645), .S1(mul_out[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_add_4_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_7 (.A0(addr_adj_3335[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3335[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23633), .COUT(n23634), .S0(addr_24__N_228[5]), 
          .S1(addr_24__N_228[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5104_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_13 (.A0(addr_adj_3335[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3335[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23636), .COUT(n23637), .S0(addr_24__N_228[11]), 
          .S1(addr_24__N_228[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5104_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_3 (.A0(addr_adj_3335[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3335[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23631), .COUT(n23632), .S0(addr_24__N_228[1]), 
          .S1(addr_24__N_228[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5104_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(addr_adj_3335[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n23631), .S1(addr_24__N_228[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5104_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5104_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_5104_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_5104_add_4_15 (.A0(addr_adj_3335[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3335[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23637), .S0(addr_24__N_228[13]), .S1(addr_24__N_228[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5104_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_5119_add_4_12 (.A0(baud_divider_adj_3392[9]), .B0(cycle_counter_adj_3488[9]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[10]), 
          .B1(cycle_counter_adj_3488[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23696), .COUT(n23697));
    defparam _add_1_5119_add_4_12.INIT0 = 16'h9995;
    defparam _add_1_5119_add_4_12.INIT1 = 16'h9995;
    defparam _add_1_5119_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_5119_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_5119_add_4_10 (.A0(baud_divider_adj_3392[7]), .B0(cycle_counter_adj_3488[7]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[8]), .B1(cycle_counter_adj_3488[8]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23695), .COUT(n23696));
    defparam _add_1_5119_add_4_10.INIT0 = 16'h9995;
    defparam _add_1_5119_add_4_10.INIT1 = 16'h9995;
    defparam _add_1_5119_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_5119_add_4_10.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync0_i5 (.D(ui_in_c_5), .CK(clk_c), .Q(ui_in_sync0[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i5.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n28626), .B(n28950), .C(time_count[0]), .D(n28624), 
         .Z(n10573)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut.init = 16'hffbf;
    GSR GSR_INST (.GSR(n32031));
    LUT4 i1_3_lut (.A(time_count[4]), .B(time_count[7]), .C(time_count[6]), 
         .Z(n28626)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 n31661_bdd_4_lut_then_4_lut (.A(is_writing), .B(fsm_state_adj_3443[1]), 
         .C(fsm_state_adj_3443[0]), .D(instr_data[13]), .Z(n32088)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam n31661_bdd_4_lut_then_4_lut.init = 16'h0020;
    LUT4 n31661_bdd_4_lut_else_4_lut (.A(fsm_state_adj_3443[1]), .B(addr_adj_3444[21]), 
         .C(fsm_state_adj_3443[0]), .D(nibbles_remaining[0]), .Z(n32087)) /* synthesis lut_function=(!(A (B+(C))+!A !(C (D)))) */ ;
    defparam n31661_bdd_4_lut_else_4_lut.init = 16'h5202;
    LUT4 i26392_2_lut (.A(time_count[2]), .B(time_count[3]), .Z(n28950)) /* synthesis lut_function=(A (B)) */ ;
    defparam i26392_2_lut.init = 16'h8888;
    FD1S3IX time_count_3561__i0 (.D(n45_adj_3282), .CK(clk_c), .CD(n780), 
            .Q(time_count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561__i0.GSR = "DISABLED";
    LUT4 i3851_4_lut_then_3_lut (.A(n31841), .B(counter_hi[4]), .C(counter_hi[3]), 
         .Z(n32101)) /* synthesis lut_function=(A+!((C)+!B)) */ ;
    defparam i3851_4_lut_then_3_lut.init = 16'haeae;
    LUT4 i3851_4_lut_else_3_lut (.A(n31841), .B(counter_hi[4]), .C(counter_hi[3]), 
         .D(counter_hi[2]), .Z(n32100)) /* synthesis lut_function=(A+!((C+!(D))+!B)) */ ;
    defparam i3851_4_lut_else_3_lut.init = 16'haeaa;
    LUT4 i23945_4_lut_then_3_lut (.A(fsm_state_adj_3443[1]), .B(instr_data[15]), 
         .C(fsm_state_adj_3443[2]), .Z(n32104)) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam i23945_4_lut_then_3_lut.init = 16'h1515;
    LUT4 i23945_4_lut_else_3_lut (.A(fsm_state_adj_3443[1]), .B(nibbles_remaining[0]), 
         .C(fsm_state_adj_3443[2]), .Z(n32103)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i23945_4_lut_else_3_lut.init = 16'h0404;
    LUT4 i1_2_lut (.A(time_count[5]), .B(time_count[1]), .Z(n28624)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 n8_bdd_4_lut (.A(n8_adj_3329), .B(n27030), .C(fsm_state_adj_3443[0]), 
         .D(qspi_data_oe[0]), .Z(qspi_data_in_3__N_1[2])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n8_bdd_4_lut.init = 16'hca00;
    LUT4 i27135_3_lut (.A(n29749), .B(n29750), .C(rs2[2]), .Z(n29752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27135_3_lut.init = 16'hcaca;
    LUT4 i15490_2_lut (.A(qspi_data_in[3]), .B(rst_reg_n), .Z(qspi_data_out_3__N_5[3])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(127[22:56])
    defparam i15490_2_lut.init = 16'h8888;
    FD1S3AX debug_rd_r_i3 (.D(debug_rd[3]), .CK(clk_c), .Q(debug_rd_r[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(257[12] 259[8])
    defparam debug_rd_r_i3.GSR = "DISABLED";
    CCU2C _add_1_5104_add_4_5 (.A0(addr_adj_3335[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3335[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23632), .COUT(n23633), .S0(addr_24__N_228[3]), 
          .S1(addr_24__N_228[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5104_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_5.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync0_i4 (.D(ui_in_c_4), .CK(clk_c), .Q(ui_in_sync0[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i4.GSR = "DISABLED";
    OB uo_out_pad_2 (.I(uo_out_c_2), .O(uo_out[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    LUT4 i27319_3_lut (.A(n29747), .B(n30906), .C(rs2[2]), .Z(n29751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27319_3_lut.init = 16'hcaca;
    FD1S3AX debug_rd_r_i2 (.D(debug_rd[2]), .CK(clk_c), .Q(debug_rd_r[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(257[12] 259[8])
    defparam debug_rd_r_i2.GSR = "DISABLED";
    LUT4 i3856_4_lut (.A(n27464), .B(n31717), .C(n6228), .D(n31712), 
         .Z(clk_c_enable_231)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C))) */ ;
    defparam i3856_4_lut.init = 16'hfcdc;
    OB uo_out_pad_3 (.I(uo_out_c_3), .O(uo_out[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    FD1S3AX debug_rd_r_i1 (.D(debug_rd[1]), .CK(clk_c), .Q(debug_rd_r[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(257[12] 259[8])
    defparam debug_rd_r_i1.GSR = "DISABLED";
    CCU2C _add_1_5119_add_4_8 (.A0(baud_divider_adj_3392[5]), .B0(cycle_counter_adj_3488[5]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[6]), .B1(cycle_counter_adj_3488[6]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23694), .COUT(n23695));
    defparam _add_1_5119_add_4_8.INIT0 = 16'h9995;
    defparam _add_1_5119_add_4_8.INIT1 = 16'h9995;
    defparam _add_1_5119_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_5119_add_4_8.INJECT1_1 = "NO";
    OB uo_out_pad_4 (.I(uo_out_c_4), .O(uo_out[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    FD1S3AX ui_in_sync0_i3 (.D(ui_in_c_3), .CK(clk_c), .Q(ui_in_sync0[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i3.GSR = "DISABLED";
    FD1P3AX gpio_out_sel_i7 (.D(gpio_out_sel_7__N_13[1]), .SP(clk_c_enable_531), 
            .CK(clk_c), .Q(gpio_out_sel[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(204[12] 211[8])
    defparam gpio_out_sel_i7.GSR = "DISABLED";
    OB uo_out_pad_5 (.I(uo_out_c_5), .O(uo_out[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_6 (.I(uo_out_c_6), .O(uo_out[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    LUT4 i1841_4_lut (.A(pc[2]), .B(n2208), .C(debug_instr_valid), .D(pc[1]), 
         .Z(n2504)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i1841_4_lut.init = 16'hc5c0;
    LUT4 n32087_bdd_4_lut (.A(n32087), .B(n32088), .C(fsm_state_adj_3443[2]), 
         .D(qspi_data_oe[0]), .Z(qspi_data_in_3__N_1[1])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;
    defparam n32087_bdd_4_lut.init = 16'h3500;
    tinyQV i_tinyqv (.rst_reg_n_adj_17(rst_reg_n_adj_3274), .clk_c(clk_c), 
           .rst_reg_n(rst_reg_n), .data_out_hold(data_out_hold), .data_ready_r_N_2792(data_ready_r_N_2792), 
           .n31883(n31883), .clk_c_enable_387(clk_c_enable_387), .\addr[10] (addr[10]), 
           .n26205(n26205), .n8819(n8819), .\addr[8] (addr[8]), .clk_c_enable_36(clk_c_enable_36), 
           .n31958(n31958), .n28276(n28276), .n26216(n26216), .n31936(n31936), 
           .clk_c_enable_395(clk_c_enable_395), .\addr[2] (addr[2]), .\addr[9] (addr[9]), 
           .n32033(n32033), .n10467(n10467), .n31934(n31934), .n31880(n31880), 
           .data_ready_r(data_ready_r), .n18241(n18241), .n31977(n31977), 
           .n26036(n26036), .data_stall(data_stall), .n29198(n29198), 
           .n31930(n31930), .clk_c_enable_445(clk_c_enable_445), .is_writing(is_writing), 
           .stop_txn_now_N_2363(stop_txn_now_N_2363), .n31713(n31713), .\instr_addr_23__N_318[7] (instr_addr_23__N_318[7]), 
           .\instr_addr_23__N_318[11] (instr_addr_23__N_318[11]), .instr_active_N_2106(instr_active_N_2106), 
           .\instr_addr_23__N_318[9] (instr_addr_23__N_318[9]), .\instr_addr_23__N_318[12] (instr_addr_23__N_318[12]), 
           .n10500(n10500), .\instr_addr_23__N_318[13] (instr_addr_23__N_318[13]), 
           .\instr_addr_23__N_318[3] (instr_addr_23__N_318[3]), .\addr[4] (addr[4]), 
           .\instr_addr_23__N_318[22] (instr_addr_23__N_318[22]), .\instr_addr_23__N_318[10] (instr_addr_23__N_318[10]), 
           .\instr_addr_23__N_318[4] (instr_addr_23__N_318[4]), .\addr[5] (addr[5]), 
           .\instr_data[15] (instr_data[15]), .\instr_data[13] (instr_data[13]), 
           .\instr_addr_23__N_318[8] (instr_addr_23__N_318[8]), .\instr_addr_23__N_318[6] (instr_addr_23__N_318[6]), 
           .\addr[7] (addr[7]), .\instr_addr_23__N_318[5] (instr_addr_23__N_318[5]), 
           .\addr[6] (addr[6]), .\instr_addr_23__N_318[14] (instr_addr_23__N_318[14]), 
           .\instr_addr_23__N_318[15] (instr_addr_23__N_318[15]), .\instr_addr_23__N_318[16] (instr_addr_23__N_318[16]), 
           .\instr_addr_23__N_318[17] (instr_addr_23__N_318[17]), .\instr_addr_23__N_318[18] (instr_addr_23__N_318[18]), 
           .\instr_addr_23__N_318[19] (instr_addr_23__N_318[19]), .\instr_addr_23__N_318[20] (instr_addr_23__N_318[20]), 
           .\instr_addr_23__N_318[21] (instr_addr_23__N_318[21]), .\instr_addr_23__N_318[2] (instr_addr_23__N_318[2]), 
           .\addr[3] (addr[3]), .\instr_addr[1] (instr_addr[1]), .data_stall_N_2158(data_stall_N_2158), 
           .continue_txn_N_2131(continue_txn_N_2131), .n10499(n10499), .data_to_write({Open_4, 
           Open_5, Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, 
           Open_12, Open_13, Open_14, Open_15, Open_16, Open_17, 
           Open_18, Open_19, Open_20, Open_21, Open_22, Open_23, 
           Open_24, Open_25, Open_26, Open_27, Open_28, Open_29, 
           Open_30, Open_31, Open_32, Open_33, Open_34, data_to_write[0]}), 
           .\data_to_write[12] (data_to_write[12]), .\data_to_write[11] (data_to_write[11]), 
           .\data_to_write[10] (data_to_write[10]), .\data_to_write[9] (data_to_write[9]), 
           .\data_to_write[8] (data_to_write[8]), .\data_to_write[7] (data_to_write[7]), 
           .\data_to_write[6] (data_to_write[6]), .\data_to_write[5] (data_to_write[5]), 
           .\data_to_write[4] (data_to_write[4]), .\data_to_write[3] (data_to_write[3]), 
           .\data_to_write[2] (data_to_write[2]), .\data_to_write[1] (data_to_write[1]), 
           .n31716(n31716), .is_writing_N_2331(is_writing_N_2331), .n33479(n33479), 
           .fsm_state({fsm_state_adj_3443}), .clk_c_enable_231(clk_c_enable_231), 
           .n31717(n31717), .clk_c_enable_186(clk_c_enable_186), .qspi_ram_b_select(qspi_ram_b_select), 
           .clk_c_enable_239(clk_c_enable_239), .qspi_ram_a_select(qspi_ram_a_select), 
           .n29199(n29199), .\qspi_data_out_3__N_5[0] (qspi_data_out_3__N_5[0]), 
           .\nibbles_remaining[0] (nibbles_remaining[0]), .n32077(n32077), 
           .clk_c_enable_452(clk_c_enable_452), .n31906(n31906), .n6228(n6228), 
           .n1084(n1084), .\writing_N_164[3] (writing_N_164[3]), .n31971(n31971), 
           .n27464(n27464), .clk_N_45(clk_N_45), .\qspi_data_out_3__N_5[2] (qspi_data_out_3__N_5[2]), 
           .n27081(n27081), .\qspi_data_oe[0] (qspi_data_oe[0]), .clk_c_enable_324(clk_c_enable_324), 
           .stop_txn_reg(stop_txn_reg), .n8135(n8135), .debug_stop_txn(debug_stop_txn), 
           .n31950(n31950), .\qspi_data_in[0] (qspi_data_in[0]), .\qspi_data_out_3__N_5[3] (qspi_data_out_3__N_5[3]), 
           .\qspi_data_in_3__N_1[0] (qspi_data_in_3__N_1[0]), .\addr[21] (addr_adj_3444[21]), 
           .spi_clk_pos_derived_59(spi_clk_pos_derived_59), .qspi_clk_N_56(qspi_clk_N_56), 
           .n31712(n31712), .n27030(n27030), .n8(n8_adj_3329), .n3(n3_adj_3332), 
           .n6232(n6232), .n27620(n27620), .n27183(n27183), .\qspi_data_in[2] (qspi_data_in[2]), 
           .\qspi_data_in[3] (qspi_data_in[3]), .\instr_addr_23__N_318[0] (instr_addr_23__N_318[0]), 
           .n31593(n31593), .\data_from_read[2] (data_from_read[2]), .counter_hi({counter_hi}), 
           .was_early_branch(was_early_branch), .\rd[0] (rd[0]), .\rs1[0] (rs1[0]), 
           .\addr[27] (addr[27]), .\instr_write_offset[3] (instr_write_offset[3]), 
           .n31860(n31860), .rs2({rs2}), .\instr_len[2] (instr_len[2]), 
           .n31869(n31869), .debug_instr_valid(debug_instr_valid), .\pc[1] (pc[1]), 
           .\pc[2] (pc[2]), .n2565(n2565), .n2208(n2208), .n31742(n31742), 
           .\data_out_slice[3] (data_out_slice[3]), .n31879(n31879), .n19(n19), 
           .n31885(n31885), .\peri_data_out[9] (peri_data_out[9]), .n4(n4_adj_3330), 
           .n31865(n31865), .n31944(n31944), .n2524(n2524), .n2504(n2504), 
           .VCC_net(VCC_net), .n31997(n31997), .n31902(n31902), .\pc[5] (pc[5]), 
           .\pc[13] (pc[13]), .n28964(n28964), .\peri_data_out[6] (peri_data_out[6]), 
           .n31867(n31867), .n4_adj_18(n4_adj_3290), .n4263(n4263), .\pc[9] (pc[9]), 
           .\imm[23] (imm[23]), .\imm[22] (imm[22]), .\imm[21] (imm[21]), 
           .\imm[20] (imm[20]), .\imm[19] (imm[19]), .\imm[18] (imm[18]), 
           .\imm[17] (imm[17]), .\imm[16] (imm[16]), .\imm[15] (imm[15]), 
           .\imm[14] (imm[14]), .\imm[13] (imm[13]), .\imm[12] (imm[12]), 
           .\imm[11] (imm[11]), .\imm[10] (imm[10]), .\imm[9] (imm[9]), 
           .\imm[8] (imm[8]), .\imm[7] (imm[7]), .\imm[6] (imm[6]), .\imm[5] (imm[5]), 
           .\imm[4] (imm[4]), .\imm[3] (imm[3]), .\imm[2] (imm[2]), .\imm[1] (imm[1]), 
           .n32035(n32035), .n32019(n32019), .n31900(n31900), .n26266(n26266), 
           .n31901(n31901), .n80(n80), .n31868(n31868), .n31978(n31978), 
           .n31847(n31847), .instr_complete_N_1647(instr_complete_N_1647), 
           .n2152(n2152), .\early_branch_addr[2] (early_branch_addr[2]), 
           .n31863(n31863), .\instr_data[1][7] (\instr_data[1] [7]), .\instr_data[2][7] (\instr_data[2] [7]), 
           .n31853(n31853), .n31849(n31849), .\instr_data[3][7] (\instr_data[3] [7]), 
           .n32055(n32055), .\debug_rd_3__N_405[31] (debug_rd_3__N_405[31]), 
           .\next_pc_for_core[6] (next_pc_for_core[6]), .n2136(n2136), .n2514(n2514), 
           .\next_pc_for_core[4] (next_pc_for_core[4]), .\next_pc_for_core[9] (next_pc_for_core[9]), 
           .\next_pc_for_core[13] (next_pc_for_core[13]), .\next_pc_for_core[10] (next_pc_for_core[10]), 
           .\next_pc_for_core[14] (next_pc_for_core[14]), .\peri_data_out[10] (peri_data_out[10]), 
           .n31761(n31761), .\cycle[0] (cycle[0]), .data_out_3__N_1385(data_out_3__N_1385), 
           .is_ret_de(is_ret_de), .n32027(n32027), .clk_c_enable_268(clk_c_enable_268), 
           .\next_pc_for_core[8] (next_pc_for_core[8]), .\next_pc_for_core[12] (next_pc_for_core[12]), 
           .n31905(n31905), .n28760(n28760), .\next_pc_for_core[3] (next_pc_for_core[3]), 
           .\pc[23] (pc[23]), .\pc[22] (pc[22]), .\pc[21] (pc[21]), .\pc[20] (pc[20]), 
           .\pc[19] (pc[19]), .\pc[18] (pc[18]), .\pc[17] (pc[17]), .\pc[16] (pc[16]), 
           .\pc[15] (pc[15]), .\pc[14] (pc[14]), .\pc[12] (pc[12]), .\pc[11] (pc[11]), 
           .\pc[10] (pc[10]), .\pc[8] (pc[8]), .\pc[7] (pc[7]), .\next_pc_for_core[5] (next_pc_for_core[5]), 
           .\pc[6] (pc[6]), .\pc[4] (pc[4]), .\next_pc_for_core[7] (next_pc_for_core[7]), 
           .n84(n84), .\next_pc_for_core[11] (next_pc_for_core[11]), .\next_pc_for_core[15] (next_pc_for_core[15]), 
           .\pc[3] (pc[3]), .\early_branch_addr[5] (early_branch_addr[5]), 
           .n32016(n32016), .\next_pc_for_core[16] (next_pc_for_core[16]), 
           .\early_branch_addr[6] (early_branch_addr[6]), .\next_pc_for_core[17] (next_pc_for_core[17]), 
           .\next_pc_for_core[18] (next_pc_for_core[18]), .\next_pc_for_core[19] (next_pc_for_core[19]), 
           .\next_pc_for_core[20] (next_pc_for_core[20]), .\early_branch_addr[4] (early_branch_addr[4]), 
           .\early_branch_addr[3] (early_branch_addr[3]), .\early_branch_addr[7] (early_branch_addr[7]), 
           .\early_branch_addr[8] (early_branch_addr[8]), .\early_branch_addr[9] (early_branch_addr[9]), 
           .\early_branch_addr[10] (early_branch_addr[10]), .\next_pc_for_core[21] (next_pc_for_core[21]), 
           .\early_branch_addr[11] (early_branch_addr[11]), .\early_branch_addr[12] (early_branch_addr[12]), 
           .\early_branch_addr[13] (early_branch_addr[13]), .\early_branch_addr[14] (early_branch_addr[14]), 
           .\early_branch_addr[15] (early_branch_addr[15]), .\next_pc_for_core[22] (next_pc_for_core[22]), 
           .\early_branch_addr[16] (early_branch_addr[16]), .\early_branch_addr[17] (early_branch_addr[17]), 
           .\next_pc_for_core[23] (next_pc_for_core[23]), .n32034(n32034), 
           .\gpio_out_sel_7__N_13[0] (gpio_out_sel_7__N_13[0]), .\early_branch_addr[18] (early_branch_addr[18]), 
           .\early_branch_addr[19] (early_branch_addr[19]), .\early_branch_addr[20] (early_branch_addr[20]), 
           .\early_branch_addr[21] (early_branch_addr[21]), .\early_branch_addr[22] (early_branch_addr[22]), 
           .\early_branch_addr[23] (early_branch_addr[23]), .n31864(n31864), 
           .n1724(n1724), .n31935(n31935), .n32021(n32021), .n32022(n32022), 
           .n31962(n31962), .n31925(n31925), .n31927(n31927), .n26282(n26282), 
           .n31964(n31964), .n31967(n31967), .n31735(n31735), .n31164(n31164), 
           .n32017(n32017), .n31163(n31163), .clk_c_enable_390(clk_c_enable_390), 
           .\data_from_read[7] (data_from_read[7]), .\data_from_read[3] (data_from_read[3]), 
           .\data_from_read[0] (data_from_read[0]), .\data_from_read[4] (data_from_read[4]), 
           .\data_from_read[8] (data_from_read[8]), .\data_from_read[12] (data_from_read[12]), 
           .\data_from_read[1] (data_from_read[1]), .\data_from_read[5] (data_from_read[5]), 
           .n31932(n31932), .n31922(n31922), .n31819(n31819), .\peri_data_out[11] (peri_data_out[11]), 
           .gpio_out_sel({gpio_out_sel}), .n14(n14_adj_3331), .n14_adj_19(n14), 
           .n31961(n31961), .n5171(n5171), .n28686(n28686), .clk_c_enable_273(clk_c_enable_273), 
           .clk_c_enable_357(clk_c_enable_357), .clk_c_enable_349(clk_c_enable_349), 
           .n32003(n32003), .clk_c_enable_259(clk_c_enable_259), .clk_c_enable_360(clk_c_enable_360), 
           .n31904(n31904), .n10573(n10573), .n31841(n31841), .n15604(n15604), 
           .n29004(n29004), .n31798(n31798), .clk_c_enable_234(clk_c_enable_234), 
           .\ui_in_sync[0] (ui_in_sync[0]), .n1160(n1160), .\alu_b_in[3] (alu_b_in[3]), 
           .debug_rd({debug_rd}), .\ui_in_sync[1] (ui_in_sync[1]), .\next_fsm_state_3__N_3015[3] (next_fsm_state_3__N_3015[3]), 
           .fsm_state_adj_25({fsm_state_adj_3466}), .accum({accum}), .d_3__N_1868({d_3__N_1868}), 
           .n31929(n31929), .\mul_out[1] (mul_out[1]), .\mul_out[2] (mul_out[2]), 
           .\mul_out[3] (mul_out[3]), .n31963(n31963), .next_bit(next_bit_adj_3308), 
           .n28800(n28800), .n31389(n31389), .alu_b_in_3__N_1504(alu_b_in_3__N_1504), 
           .n29162(n29162), .n18086(n18086), .\csr_read_3__N_1447[2] (csr_read_3__N_1447[2]), 
           .GND_net(GND_net), .\next_accum[5] (next_accum[5]), .\next_accum[6] (next_accum[6]), 
           .\next_accum[7] (next_accum[7]), .\next_accum[8] (next_accum[8]), 
           .\next_accum[9] (next_accum[9]), .\next_accum[10] (next_accum[10]), 
           .\next_accum[11] (next_accum[11]), .\next_accum[12] (next_accum[12]), 
           .\next_accum[13] (next_accum[13]), .\next_accum[14] (next_accum[14]), 
           .\next_accum[15] (next_accum[15]), .\next_accum[16] (next_accum[16]), 
           .\next_accum[17] (next_accum[17]), .\next_accum[18] (next_accum[18]), 
           .\next_accum[19] (next_accum[19]), .\next_accum[4] (next_accum[4]), 
           .n12(n12), .n11(n11), .n9(n9), .n8_adj_23(n8), .\registers[5][7] (\registers[5] [7]), 
           .\registers[6][7] (\registers[6] [7]), .\registers[7][7] (\registers[7] [7]), 
           .n29747(n29747), .n4_adj_24(n4)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(111[12] 150[6])
    LUT4 n15604_bdd_3_lut_28129 (.A(\registers[7] [7]), .B(\registers[6] [7]), 
         .C(rs2[0]), .Z(n30904)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n15604_bdd_3_lut_28129.init = 16'hacac;
    FD1S3AX ui_in_sync_i7 (.D(ui_in_sync0[7]), .CK(clk_c), .Q(ui_in_sync[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i7.GSR = "DISABLED";
    LUT4 i27016_3_lut (.A(\gpio_out_func_sel[6] [3]), .B(\gpio_out_func_sel[7] [3]), 
         .C(addr[2]), .Z(n29633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27016_3_lut.init = 16'hcaca;
    CCU2C _add_1_5104_add_4_11 (.A0(addr_adj_3335[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3335[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23635), .COUT(n23636), .S0(addr_24__N_228[9]), 
          .S1(addr_24__N_228[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5104_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_11.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync0_i2 (.D(ui_in_c_2), .CK(clk_c), .Q(ui_in_sync0[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i2.GSR = "DISABLED";
    FD1S3AX ui_in_sync_i6 (.D(ui_in_sync0[6]), .CK(clk_c), .Q(ui_in_sync[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i6.GSR = "DISABLED";
    CCU2C _add_1_5119_add_4_6 (.A0(baud_divider_adj_3392[3]), .B0(cycle_counter_adj_3488[3]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[4]), .B1(cycle_counter_adj_3488[4]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23693), .COUT(n23694));
    defparam _add_1_5119_add_4_6.INIT0 = 16'h9995;
    defparam _add_1_5119_add_4_6.INIT1 = 16'h9995;
    defparam _add_1_5119_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_5119_add_4_6.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_604 (.A(addr[6]), .B(\uo_out_from_user_peri[1] [3]), 
         .C(n24), .D(n31922), .Z(n1)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i1_4_lut_adj_604.init = 16'ha088;
    FD1S3AX ui_in_sync_i5 (.D(ui_in_sync0[5]), .CK(clk_c), .Q(ui_in_sync[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i5.GSR = "DISABLED";
    FD1S3AX ui_in_sync0_i1 (.D(ui_in_c_1), .CK(clk_c), .Q(ui_in_sync0[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i1.GSR = "DISABLED";
    IB ui_in_pad_0 (.I(ui_in[0]), .O(ui_in_c_0));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    FD1S3AX ui_in_sync_i4 (.D(ui_in_sync0[4]), .CK(clk_c), .Q(ui_in_sync[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i4.GSR = "DISABLED";
    OB uo_out_pad_7 (.I(uo_out_c_7), .O(uo_out[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    IB ui_in_pad_1 (.I(ui_in[1]), .O(ui_in_c_1));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_2 (.I(ui_in[2]), .O(ui_in_c_2));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_3 (.I(ui_in[3]), .O(ui_in_c_3));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_4 (.I(ui_in[4]), .O(ui_in_c_4));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_5 (.I(ui_in[5]), .O(ui_in_c_5));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_6 (.I(ui_in[6]), .O(ui_in_c_6));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB ui_in_pad_7 (.I(ui_in[7]), .O(ui_in_c_7));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(12[26:31])
    IB rst_n_pad (.I(rst_n), .O(rst_n_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(10[20:25])
    IB clk_pad (.I(clk), .O(clk_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    OB uo_out_pad_0 (.I(uo_out_c_0), .O(uo_out[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    OB uo_out_pad_1 (.I(uo_out_c_1), .O(uo_out[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(13[27:33])
    CCU2C _add_1_5119_add_4_4 (.A0(baud_divider_adj_3392[1]), .B0(cycle_counter_adj_3488[1]), 
          .C0(GND_net), .D0(VCC_net), .A1(baud_divider_adj_3392[2]), .B1(cycle_counter_adj_3488[2]), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23692), .COUT(n23693));
    defparam _add_1_5119_add_4_4.INIT0 = 16'h9995;
    defparam _add_1_5119_add_4_4.INIT1 = 16'h9995;
    defparam _add_1_5119_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_5119_add_4_4.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync0_i0 (.D(ui_in_c_0), .CK(clk_c), .Q(ui_in_sync0[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i0.GSR = "DISABLED";
    FD1P3AX debug_register_data_58 (.D(n7884), .SP(clk_c_enable_355), .CK(clk_c), 
            .Q(debug_register_data));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(250[12] 255[8])
    defparam debug_register_data_58.GSR = "DISABLED";
    LUT4 n15604_bdd_3_lut_28567 (.A(n15604), .B(\registers[5] [7]), .C(rs2[0]), 
         .Z(n30905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n15604_bdd_3_lut_28567.init = 16'hcaca;
    CCU2C _add_1_5119_add_4_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(baud_divider_adj_3392[0]), .B1(cycle_counter_adj_3488[0]), 
          .C1(GND_net), .D1(VCC_net), .COUT(n23692));
    defparam _add_1_5119_add_4_2.INIT0 = 16'h000f;
    defparam _add_1_5119_add_4_2.INIT1 = 16'h9995;
    defparam _add_1_5119_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_5119_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_21 (.A0(pc[22]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[23]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23690), .S0(next_pc_for_core[22]), .S1(next_pc_for_core[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_21.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync_i3 (.D(ui_in_sync0[3]), .CK(clk_c), .Q(ui_in_sync[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i3.GSR = "DISABLED";
    CCU2C _add_1_5110_add_4_19 (.A0(pc[20]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[21]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23689), .COUT(n23690), .S0(next_pc_for_core[20]), .S1(next_pc_for_core[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_19.INJECT1_1 = "NO";
    FD1S3AX ui_in_sync_i2 (.D(ui_in_sync0[2]), .CK(clk_c), .Q(ui_in_sync[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i2.GSR = "DISABLED";
    FD1S3AX ui_in_sync_i1 (.D(ui_in_sync0[1]), .CK(clk_c), .Q(ui_in_sync[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i1.GSR = "DISABLED";
    FD1S3AX ui_in_sync0_i7 (.D(ui_in_c_7), .CK(clk_c), .Q(ui_in_sync0[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i7.GSR = "DISABLED";
    FD1S3AX ui_in_sync0_i6 (.D(ui_in_c_6), .CK(clk_c), .Q(ui_in_sync0[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync0_i6.GSR = "DISABLED";
    CCU2C _add_1_5110_add_4_17 (.A0(pc[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[19]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23688), .COUT(n23689), .S0(next_pc_for_core[18]), .S1(next_pc_for_core[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_17.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_639_4_lut (.A(clk_c_enable_268), .B(n31904), .C(n32027), 
         .D(n32034), .Z(n31844)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_3_lut_rep_639_4_lut.init = 16'h0020;
    LUT4 i1_4_lut_adj_605 (.A(n28230), .B(n29004), .C(n28246), .D(n31867), 
         .Z(is_ret_de)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_605.init = 16'h0020;
    LUT4 i1_3_lut_adj_606 (.A(n31869), .B(n31868), .C(n31864), .Z(n28230)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_606.init = 16'h4040;
    LUT4 i1_4_lut_adj_607 (.A(n28242), .B(n31863), .C(n31847), .D(n31860), 
         .Z(n28246)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_607.init = 16'h0200;
    CCU2C _add_1_5110_add_4_15 (.A0(pc[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[17]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23687), .COUT(n23688), .S0(next_pc_for_core[16]), .S1(next_pc_for_core[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_15.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_608 (.A(n31853), .B(n31798), .C(n31849), .D(n31865), 
         .Z(n28242)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_608.init = 16'h0004;
    LUT4 i1_4_lut_adj_609 (.A(n31879), .B(n19), .C(peri_data_out[2]), 
         .D(n4_adj_3330), .Z(data_from_read[2])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_609.init = 16'heeec;
    LUT4 i1_4_lut_adj_610 (.A(n31879), .B(n19), .C(peri_data_out[5]), 
         .D(n4_adj_3330), .Z(data_from_read[5])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_610.init = 16'heeec;
    LUT4 i1_4_lut_adj_611 (.A(n31879), .B(n19), .C(peri_data_out[1]), 
         .D(n4_adj_3330), .Z(data_from_read[1])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_611.init = 16'heeec;
    LUT4 i1_4_lut_adj_612 (.A(n31879), .B(n19), .C(peri_data_out[12]), 
         .D(n4_adj_3330), .Z(data_from_read[12])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_612.init = 16'heeec;
    CCU2C _add_1_5110_add_4_13 (.A0(pc[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[15]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23686), .COUT(n23687), .S0(next_pc_for_core[14]), .S1(next_pc_for_core[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_13.INJECT1_1 = "NO";
    FD1S3IX time_count_3561__i1 (.D(n44), .CK(clk_c), .CD(n780), .Q(time_count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561__i1.GSR = "DISABLED";
    LUT4 i15121_3_lut (.A(\instr_data[2] [7]), .B(\instr_data[3] [7]), .C(n2524), 
         .Z(n9_adj_3328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15121_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_613 (.A(n31879), .B(n19), .C(peri_data_out[8]), 
         .D(n4_adj_3330), .Z(data_from_read[8])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_613.init = 16'heeec;
    LUT4 i1_4_lut_adj_614 (.A(n31879), .B(n19), .C(peri_data_out[4]), 
         .D(n4_adj_3330), .Z(data_from_read[4])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_614.init = 16'heeec;
    LUT4 i15425_4_lut (.A(n5171), .B(data_from_read[31]), .C(peri_data_out[0]), 
         .D(n31879), .Z(data_from_read[0])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i15425_4_lut.init = 16'hfcee;
    LUT4 i1_4_lut_adj_615 (.A(n31879), .B(n19), .C(peri_data_out[3]), 
         .D(n4_adj_3330), .Z(data_from_read[3])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_615.init = 16'heeec;
    LUT4 i1_4_lut_adj_616 (.A(next_fsm_state_3__N_3015[3]), .B(rst_reg_n), 
         .C(n28850), .D(fsm_state_adj_3489[2]), .Z(n27347)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_616.init = 16'h0040;
    LUT4 i1_3_lut_adj_617 (.A(fsm_state_adj_3489[0]), .B(fsm_state_adj_3489[3]), 
         .C(fsm_state_adj_3489[1]), .Z(n28850)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_617.init = 16'h8080;
    CCU2C _add_1_5110_add_4_11 (.A0(pc[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[13]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23685), .COUT(n23686), .S0(next_pc_for_core[12]), .S1(next_pc_for_core[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_618 (.A(peri_data_out[7]), .B(n28966), .C(n31879), 
         .D(n10467), .Z(data_from_read[7])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i1_4_lut_adj_618.init = 16'hffec;
    CCU2C _add_1_5110_add_4_9 (.A0(pc[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[11]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23684), .COUT(n23685), .S0(next_pc_for_core[10]), .S1(next_pc_for_core[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_7 (.A0(pc[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[9]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23683), .COUT(n23684), .S0(next_pc_for_core[8]), .S1(next_pc_for_core[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_7.INJECT1_1 = "NO";
    FD1S3IX time_count_3561__i2 (.D(n43), .CK(clk_c), .CD(n780), .Q(time_count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561__i2.GSR = "DISABLED";
    FD1S3IX time_count_3561__i3 (.D(n42_adj_3278), .CK(clk_c), .CD(n780), 
            .Q(time_count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561__i3.GSR = "DISABLED";
    FD1S3IX time_count_3561__i4 (.D(n41), .CK(clk_c), .CD(n780), .Q(time_count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561__i4.GSR = "DISABLED";
    FD1S3IX time_count_3561__i5 (.D(n40), .CK(clk_c), .CD(n780), .Q(time_count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561__i5.GSR = "DISABLED";
    FD1S3IX time_count_3561__i6 (.D(n39), .CK(clk_c), .CD(n780), .Q(time_count[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561__i6.GSR = "DISABLED";
    FD1S3IX time_count_3561__i7 (.D(n38), .CK(clk_c), .CD(n780), .Q(time_count[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561__i7.GSR = "DISABLED";
    CCU2C _add_1_5110_add_4_5 (.A0(pc[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[7]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23682), .COUT(n23683), .S0(next_pc_for_core[6]), .S1(next_pc_for_core[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_5110_add_4_3 (.A0(pc[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[5]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23681), .COUT(n23682), .S0(next_pc_for_core[4]), .S1(next_pc_for_core[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_5110_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_5110_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_3.INJECT1_1 = "NO";
    LUT4 n29633_bdd_3_lut_28369 (.A(\gpio_out_func_sel[4] [3]), .B(addr[2]), 
         .C(\gpio_out_func_sel[5] [3]), .Z(n31059)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n29633_bdd_3_lut_28369.init = 16'he2e2;
    CCU2C _add_1_5110_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pc[3]), .B1(n32055), .C1(instr_len[2]), 
          .D1(pc[2]), .COUT(n23681), .S1(next_pc_for_core[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(377[27:85])
    defparam _add_1_5110_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5110_add_4_1.INIT1 = 16'h566a;
    defparam _add_1_5110_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5110_add_4_1.INJECT1_1 = "NO";
    LUT4 i1836_4_lut (.A(pc[2]), .B(n2565), .C(debug_instr_valid), .D(pc[1]), 
         .Z(n2524)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i1836_4_lut.init = 16'hcac0;
    LUT4 \gpio_out_func_sel_0[[3__bdd_3_lut_28226  (.A(\gpio_out_func_sel[2] [3]), 
         .B(addr[2]), .C(\gpio_out_func_sel[3] [3]), .Z(n31061)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam \gpio_out_func_sel_0[[3__bdd_3_lut_28226 .init = 16'he2e2;
    LUT4 \gpio_out_func_sel_0[[3__bdd_3_lut_28370  (.A(\gpio_out_func_sel[0] [3]), 
         .B(\gpio_out_func_sel[1] [3]), .C(addr[2]), .Z(n31062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \gpio_out_func_sel_0[[3__bdd_3_lut_28370 .init = 16'hcaca;
    PFUMX i28300 (.BLUT(n31163), .ALUT(n31162), .C0(n2136), .Z(n31164));
    VLO i1 (.Z(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i27780_3_lut (.A(n31879), .B(n19), .C(n31885), .Z(data_from_read[31])) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i27780_3_lut.init = 16'hcece;
    CCU2C _add_1_5104_add_4_9 (.A0(addr_adj_3335[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(addr_adj_3335[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23634), .COUT(n23635), .S0(addr_24__N_228[7]), 
          .S1(addr_24__N_228[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(87[25:33])
    defparam _add_1_5104_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_5104_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_5104_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5104_add_4_9.INJECT1_1 = "NO";
    FD1P3AX gpio_out_sel_i6 (.D(gpio_out_sel_7__N_13[0]), .SP(clk_c_enable_531), 
            .CK(clk_c), .Q(gpio_out_sel[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(204[12] 211[8])
    defparam gpio_out_sel_i6.GSR = "DISABLED";
    LUT4 i26408_4_lut (.A(n31934), .B(n32027), .C(addr[4]), .D(n14_adj_3331), 
         .Z(n28966)) /* synthesis lut_function=(!(A+(B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i26408_4_lut.init = 16'h1511;
    LUT4 i26406_4_lut (.A(n31934), .B(n32027), .C(addr[4]), .D(n14), 
         .Z(n28964)) /* synthesis lut_function=(!(A+(B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(193[9] 198[16])
    defparam i26406_4_lut.init = 16'h1511;
    LUT4 i21233_2_lut_rep_811 (.A(imm[1]), .B(pc[1]), .Z(n32016)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i21233_2_lut_rep_811.init = 16'h6666;
    LUT4 instr_addr_23__I_0_i1_3_lut_4_lut (.A(imm[1]), .B(pc[1]), .C(was_early_branch), 
         .D(instr_addr_23__N_318[0]), .Z(instr_addr[1])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam instr_addr_23__I_0_i1_3_lut_4_lut.init = 16'h6f60;
    LUT4 n3_bdd_4_lut (.A(n3_adj_3332), .B(n32105), .C(fsm_state_adj_3443[0]), 
         .D(qspi_data_oe[0]), .Z(qspi_data_in_3__N_1[3])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;
    defparam n3_bdd_4_lut.init = 16'h3500;
    LUT4 i6037_2_lut_rep_822 (.A(addr[3]), .B(addr[2]), .Z(n32027)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6037_2_lut_rep_822.init = 16'h8888;
    LUT4 i1_2_lut_rep_718_3_lut_4_lut (.A(addr[3]), .B(addr[2]), .C(n32035), 
         .D(addr[5]), .Z(n31923)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_718_3_lut_4_lut.init = 16'hf7ff;
    LUT4 i25_4_lut (.A(ui_in_sync[3]), .B(n31962), .C(n31935), .D(n31064), 
         .Z(n24)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    defparam i25_4_lut.init = 16'h3a0a;
    LUT4 i1_2_lut_adj_619 (.A(addr[4]), .B(addr[5]), .Z(n28686)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_619.init = 16'h8888;
    CCU2C time_count_3561_add_4_9 (.A0(time_count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23670), .S0(n38));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561_add_4_9.INIT0 = 16'haaa0;
    defparam time_count_3561_add_4_9.INIT1 = 16'h0000;
    defparam time_count_3561_add_4_9.INJECT1_0 = "NO";
    defparam time_count_3561_add_4_9.INJECT1_1 = "NO";
    L6MUX21 i28229 (.D0(n31063), .D1(n31060), .SD(addr[4]), .Z(n31064));
    FD1S3AX ui_in_sync_i0 (.D(ui_in_sync0[0]), .CK(clk_c), .Q(ui_in_sync[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(103[12] 106[8])
    defparam ui_in_sync_i0.GSR = "DISABLED";
    LUT4 i26581_3_lut (.A(data_stall), .B(data_stall_N_2158), .C(continue_txn_N_2131), 
         .Z(n29198)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam i26581_3_lut.init = 16'hcece;
    PFUMX i28227 (.BLUT(n31062), .ALUT(n31061), .C0(addr[3]), .Z(n31063));
    PFUMX i28224 (.BLUT(n31059), .ALUT(n29633), .C0(addr[3]), .Z(n31060));
    CCU2C time_count_3561_add_4_7 (.A0(time_count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23669), .COUT(n23670), .S0(n40), .S1(n39));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561_add_4_7.INIT0 = 16'haaa0;
    defparam time_count_3561_add_4_7.INIT1 = 16'haaa0;
    defparam time_count_3561_add_4_7.INJECT1_0 = "NO";
    defparam time_count_3561_add_4_7.INJECT1_1 = "NO";
    CCU2C time_count_3561_add_4_5 (.A0(time_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23668), .COUT(n23669), .S0(n42_adj_3278), 
          .S1(n41));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561_add_4_5.INIT0 = 16'haaa0;
    defparam time_count_3561_add_4_5.INIT1 = 16'haaa0;
    defparam time_count_3561_add_4_5.INJECT1_0 = "NO";
    defparam time_count_3561_add_4_5.INJECT1_1 = "NO";
    CCU2C time_count_3561_add_4_3 (.A0(time_count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(time_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23667), .COUT(n23668), .S0(n44), .S1(n43));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561_add_4_3.INIT0 = 16'haaa0;
    defparam time_count_3561_add_4_3.INIT1 = 16'haaa0;
    defparam time_count_3561_add_4_3.INJECT1_0 = "NO";
    defparam time_count_3561_add_4_3.INJECT1_1 = "NO";
    CCU2C time_count_3561_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(time_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n23667), .S1(n45_adj_3282));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(244[32:46])
    defparam time_count_3561_add_4_1.INIT0 = 16'h0000;
    defparam time_count_3561_add_4_1.INIT1 = 16'h555f;
    defparam time_count_3561_add_4_1.INJECT1_0 = "NO";
    defparam time_count_3561_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_5113_add_4_24 (.A0(imm[23]), .B0(pc[23]), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23666), .S0(early_branch_addr[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_24.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_24.INIT1 = 16'h0000;
    defparam _add_1_5113_add_4_24.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_24.INJECT1_1 = "NO";
    CCU2C _add_1_5113_add_4_22 (.A0(imm[21]), .B0(pc[21]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[22]), .B1(pc[22]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23665), .COUT(n23666), .S0(early_branch_addr[21]), .S1(early_branch_addr[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_22.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_22.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_22.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_22.INJECT1_1 = "NO";
    LUT4 instr_1__bdd_3_lut_28478 (.A(n31742), .B(n31853), .C(rd[0]), 
         .Z(n31162)) /* synthesis lut_function=(!(A (C)+!A !(B))) */ ;
    defparam instr_1__bdd_3_lut_28478.init = 16'h4e4e;
    CCU2C _add_1_5113_add_4_20 (.A0(imm[19]), .B0(pc[19]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[20]), .B1(pc[20]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23664), .COUT(n23665), .S0(early_branch_addr[19]), .S1(early_branch_addr[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_20.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_20.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_5113_add_4_18 (.A0(imm[17]), .B0(pc[17]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[18]), .B1(pc[18]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23663), .COUT(n23664), .S0(early_branch_addr[17]), .S1(early_branch_addr[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_18.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_18.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_18.INJECT1_1 = "NO";
    CCU2C _add_1_5122_add_4_13 (.A0(cycle_counter_adj_3465[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3465[12]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n23732), .S0(n33), 
          .S1(n30));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5122_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_5122_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_5122_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5122_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_5113_add_4_16 (.A0(imm[15]), .B0(pc[15]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[16]), .B1(pc[16]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23662), .COUT(n23663), .S0(early_branch_addr[15]), .S1(early_branch_addr[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_16.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_620 (.A(n31880), .B(n31879), .C(addr[2]), .D(n28538), 
         .Z(debug_uart_tx_start)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_620.init = 16'h0200;
    LUT4 i1_2_lut_adj_621 (.A(addr[3]), .B(addr[4]), .Z(n28538)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_621.init = 16'h8888;
    CCU2C _add_1_5113_add_4_14 (.A0(imm[13]), .B0(pc[13]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[14]), .B1(pc[14]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23661), .COUT(n23662), .S0(early_branch_addr[13]), .S1(early_branch_addr[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_5122_add_4_11 (.A0(cycle_counter_adj_3465[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3465[10]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n23731), .COUT(n23732), 
          .S0(n39_adj_3283), .S1(n36_adj_3327));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5122_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_5122_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_5122_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5122_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_5122_add_4_9 (.A0(cycle_counter_adj_3465[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3465[8]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n23730), .COUT(n23731), 
          .S0(n45), .S1(n42_adj_3279));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5122_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_5122_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_5122_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5122_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_5113_add_4_12 (.A0(imm[11]), .B0(pc[11]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[12]), .B1(pc[12]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23660), .COUT(n23661), .S0(early_branch_addr[11]), .S1(early_branch_addr[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_5122_add_4_7 (.A0(cycle_counter_adj_3465[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3465[6]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n23729), .COUT(n23730), 
          .S0(n51), .S1(n48));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5122_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_5122_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_5122_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5122_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_5113_add_4_10 (.A0(imm[9]), .B0(pc[9]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[10]), .B1(pc[10]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23659), .COUT(n23660), .S0(early_branch_addr[9]), .S1(early_branch_addr[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_10.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_10.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_10.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_10.INJECT1_1 = "NO";
    CCU2C _add_1_5122_add_4_5 (.A0(cycle_counter_adj_3465[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3465[4]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n23728), .COUT(n23729), 
          .S0(n57_adj_3280), .S1(n54_adj_3281));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5122_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_5122_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_5122_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5122_add_4_5.INJECT1_1 = "NO";
    LUT4 i13073_3_lut (.A(n15604), .B(\registers[5] [7]), .C(rs1[0]), 
         .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(117[15:18])
    defparam i13073_3_lut.init = 16'hcaca;
    CCU2C _add_1_5113_add_4_8 (.A0(imm[7]), .B0(pc[7]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[8]), .B1(pc[8]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23658), .COUT(n23659), .S0(early_branch_addr[7]), .S1(early_branch_addr[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_8.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_8.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_8.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_8.INJECT1_1 = "NO";
    CCU2C _add_1_5113_add_4_6 (.A0(imm[5]), .B0(pc[5]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[6]), .B1(pc[6]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23657), .COUT(n23658), .S0(early_branch_addr[5]), .S1(early_branch_addr[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_6.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_6.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_6.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_6.INJECT1_1 = "NO";
    CCU2C _add_1_5122_add_4_3 (.A0(cycle_counter_adj_3465[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter_adj_3465[2]), 
          .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n23727), .COUT(n23728), 
          .S0(n63_adj_3286), .S1(n60));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5122_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_5122_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_5122_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5122_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5113_add_4_4 (.A0(imm[3]), .B0(pc[3]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[4]), .B1(pc[4]), .C1(GND_net), .D1(VCC_net), 
          .CIN(n23656), .COUT(n23657), .S0(early_branch_addr[3]), .S1(early_branch_addr[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_4.INIT0 = 16'h666a;
    defparam _add_1_5113_add_4_4.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_4.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_4.INJECT1_1 = "NO";
    CCU2C _add_1_5122_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycle_counter_adj_3465[0]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .COUT(n23727), .S1(n66));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5122_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5122_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_5122_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5122_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_5113_add_4_2 (.A0(imm[1]), .B0(pc[1]), .C0(GND_net), 
          .D0(VCC_net), .A1(imm[2]), .B1(pc[2]), .C1(GND_net), .D1(VCC_net), 
          .COUT(n23656), .S1(early_branch_addr[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(383[37:57])
    defparam _add_1_5113_add_4_2.INIT0 = 16'h0008;
    defparam _add_1_5113_add_4_2.INIT1 = 16'h666a;
    defparam _add_1_5113_add_4_2.INJECT1_0 = "NO";
    defparam _add_1_5113_add_4_2.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_13 (.A0(cycle_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23725), .S0(n33_adj_3276), .S1(n30_adj_3289));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5107_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_5107_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_5107_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_11 (.A0(cycle_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23724), .COUT(n23725), .S0(n39_adj_3277), 
          .S1(n36));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5107_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_5107_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_5107_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_20 (.A0(d_3__N_1868[18]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_3__N_1868[19]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23653), .S0(next_accum[18]), .S1(next_accum[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_20.INIT0 = 16'haaa0;
    defparam _add_1_add_4_add_4_20.INIT1 = 16'haaa0;
    defparam _add_1_add_4_add_4_20.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_20.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_9 (.A0(cycle_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23723), .COUT(n23724), .S0(n45_adj_3291), 
          .S1(n42));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5107_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_5107_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_5107_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_7 (.A0(cycle_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23722), .COUT(n23723), .S0(n51_adj_3275), 
          .S1(n48_adj_3288));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5107_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_5107_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_5107_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_5 (.A0(cycle_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23721), .COUT(n23722), .S0(n57), .S1(n54));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5107_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_5107_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_5107_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_3 (.A0(cycle_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23720), .COUT(n23721), .S0(n63), .S1(n60_adj_3284));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5107_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_5107_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_5107_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_5107_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycle_counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n23720), .S1(n66_adj_3285));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(105[26:46])
    defparam _add_1_5107_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_5107_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_5107_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_5107_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_18 (.A0(d_3__N_1868[16]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(d_3__N_1868[17]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23652), .COUT(n23653), .S0(next_accum[16]), 
          .S1(next_accum[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_18.INIT0 = 16'haaa0;
    defparam _add_1_add_4_add_4_18.INIT1 = 16'haaa0;
    defparam _add_1_add_4_add_4_18.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_18.INJECT1_1 = "NO";
    LUT4 i44_3_lut (.A(debug_rd_3__N_405[31]), .B(n84), .C(alu_b_in_3__N_1504), 
         .Z(alu_b_in[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(118[15:18])
    defparam i44_3_lut.init = 16'hcaca;
    CCU2C _add_1_add_4_add_4_16 (.A0(accum[14]), .B0(d_3__N_1868[14]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[15]), .B1(d_3__N_1868[15]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23651), .COUT(n23652), .S0(next_accum[14]), 
          .S1(next_accum[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_16.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_16.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_16.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_16.INJECT1_1 = "NO";
    CCU2C _add_1_5116_add_4_23 (.A0(early_branch_addr[23]), .B0(was_early_branch), 
          .C0(pc[23]), .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n23719), .S0(instr_addr_23__N_318[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_23.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_23.INIT1 = 16'h0000;
    defparam _add_1_5116_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_23.INJECT1_1 = "NO";
    CCU2C _add_1_5116_add_4_21 (.A0(early_branch_addr[21]), .B0(was_early_branch), 
          .C0(pc[21]), .D0(VCC_net), .A1(early_branch_addr[22]), .B1(was_early_branch), 
          .C1(pc[22]), .D1(VCC_net), .CIN(n23718), .COUT(n23719), .S0(instr_addr_23__N_318[20]), 
          .S1(instr_addr_23__N_318[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_21.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_21.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_14 (.A0(accum[12]), .B0(d_3__N_1868[12]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[13]), .B1(d_3__N_1868[13]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23650), .COUT(n23651), .S0(next_accum[12]), 
          .S1(next_accum[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_14.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_14.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_14.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_14.INJECT1_1 = "NO";
    CCU2C _add_1_5116_add_4_19 (.A0(early_branch_addr[19]), .B0(was_early_branch), 
          .C0(pc[19]), .D0(VCC_net), .A1(early_branch_addr[20]), .B1(was_early_branch), 
          .C1(pc[20]), .D1(VCC_net), .CIN(n23717), .COUT(n23718), .S0(instr_addr_23__N_318[18]), 
          .S1(instr_addr_23__N_318[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_19.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_19.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_add_4_add_4_12 (.A0(accum[10]), .B0(d_3__N_1868[10]), .C0(GND_net), 
          .D0(VCC_net), .A1(accum[11]), .B1(d_3__N_1868[11]), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23649), .COUT(n23650), .S0(next_accum[10]), 
          .S1(next_accum[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[36:83])
    defparam _add_1_add_4_add_4_12.INIT0 = 16'h666a;
    defparam _add_1_add_4_add_4_12.INIT1 = 16'h666a;
    defparam _add_1_add_4_add_4_12.INJECT1_0 = "NO";
    defparam _add_1_add_4_add_4_12.INJECT1_1 = "NO";
    CCU2C _add_1_5116_add_4_17 (.A0(early_branch_addr[17]), .B0(was_early_branch), 
          .C0(pc[17]), .D0(VCC_net), .A1(early_branch_addr[18]), .B1(was_early_branch), 
          .C1(pc[18]), .D1(VCC_net), .CIN(n23716), .COUT(n23717), .S0(instr_addr_23__N_318[16]), 
          .S1(instr_addr_23__N_318[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_17.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_17.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_17.INJECT1_1 = "NO";
    LUT4 i7_3_lut_rep_659 (.A(n2514), .B(n9_adj_3328), .C(n31944), .Z(n31864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i7_3_lut_rep_659.init = 16'hcaca;
    CCU2C _add_1_5116_add_4_15 (.A0(early_branch_addr[15]), .B0(was_early_branch), 
          .C0(pc[15]), .D0(VCC_net), .A1(early_branch_addr[16]), .B1(was_early_branch), 
          .C1(pc[16]), .D1(VCC_net), .CIN(n23715), .COUT(n23716), .S0(instr_addr_23__N_318[14]), 
          .S1(instr_addr_23__N_318[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_15.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_15.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(n2514), .B(n9_adj_3328), .C(n31944), .D(n31735), 
         .Z(n1724)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hffca;
    CCU2C _add_1_5116_add_4_13 (.A0(early_branch_addr[13]), .B0(was_early_branch), 
          .C0(pc[13]), .D0(VCC_net), .A1(early_branch_addr[14]), .B1(was_early_branch), 
          .C1(pc[14]), .D1(VCC_net), .CIN(n23714), .COUT(n23715), .S0(instr_addr_23__N_318[12]), 
          .S1(instr_addr_23__N_318[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_13.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_13.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_5116_add_4_11 (.A0(early_branch_addr[11]), .B0(was_early_branch), 
          .C0(pc[11]), .D0(VCC_net), .A1(early_branch_addr[12]), .B1(was_early_branch), 
          .C1(pc[12]), .D1(VCC_net), .CIN(n23713), .COUT(n23714), .S0(instr_addr_23__N_318[10]), 
          .S1(instr_addr_23__N_318[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_11.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_11.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_5116_add_4_9 (.A0(early_branch_addr[9]), .B0(was_early_branch), 
          .C0(pc[9]), .D0(VCC_net), .A1(early_branch_addr[10]), .B1(was_early_branch), 
          .C1(pc[10]), .D1(VCC_net), .CIN(n23712), .COUT(n23713), .S0(instr_addr_23__N_318[8]), 
          .S1(instr_addr_23__N_318[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_9.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_9.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_5116_add_4_7 (.A0(early_branch_addr[7]), .B0(was_early_branch), 
          .C0(pc[7]), .D0(VCC_net), .A1(early_branch_addr[8]), .B1(was_early_branch), 
          .C1(pc[8]), .D1(VCC_net), .CIN(n23711), .COUT(n23712), .S0(instr_addr_23__N_318[6]), 
          .S1(instr_addr_23__N_318[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[64:119])
    defparam _add_1_5116_add_4_7.INIT0 = 16'hb8b8;
    defparam _add_1_5116_add_4_7.INIT1 = 16'hb8b8;
    defparam _add_1_5116_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_5116_add_4_7.INJECT1_1 = "NO";
    LUT4 i26582_4_lut (.A(is_writing), .B(is_writing_N_2331), .C(n31716), 
         .D(n8135), .Z(n29199)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i26582_4_lut.init = 16'hcaaa;
    LUT4 i15186_2_lut (.A(qspi_data_in[0]), .B(rst_reg_n), .Z(qspi_data_out_3__N_5[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(127[22:56])
    defparam i15186_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_622 (.A(data_out_3__N_1385), .B(n84), .Z(data_out_slice[3])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(118[15:18])
    defparam i1_2_lut_adj_622.init = 16'h4444;
    LUT4 i3862_4_lut (.A(n32077), .B(n31717), .C(n6232), .D(n1084), 
         .Z(clk_c_enable_452)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C))) */ ;
    defparam i3862_4_lut.init = 16'hfcdc;
    PFUMX i28130 (.BLUT(n30905), .ALUT(n30904), .C0(rs2[1]), .Z(n30906));
    LUT4 i15127_3_lut (.A(\instr_data[1] [7]), .B(\instr_data[2] [7]), .C(n2504), 
         .Z(n2152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15127_3_lut.init = 16'hcaca;
    LUT4 mux_34_i2_3_lut (.A(ui_in_c_0), .B(data_to_write[7]), .C(n31844), 
         .Z(gpio_out_sel_7__N_13[1])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(209[13:93])
    defparam mux_34_i2_3_lut.init = 16'hc5c5;
    LUT4 i23_3_lut (.A(n27421), .B(debug_rd_r[3]), .C(debug_register_data), 
         .Z(uo_out_c_5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(157[24:73])
    defparam i23_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(\gpio_out_func_sel[5] [4]), .B(n10), .C(\gpio_out_func_sel[5] [3]), 
         .D(\gpio_out_func_sel[5] [2]), .Z(n27421)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0004;
    LUT4 i24_4_lut (.A(\gpio_out_func_sel[5] [1]), .B(\uo_out_from_user_peri[1] [5]), 
         .C(\gpio_out_func_sel[5] [0]), .D(\uo_out_from_user_peri[2] [7]), 
         .Z(n10)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(157[24:73])
    defparam i24_4_lut.init = 16'h4a40;
    LUT4 debug_uart_txd_I_0_3_lut (.A(debug_uart_txd), .B(peri_out[6]), 
         .C(gpio_out_sel[6]), .Z(uo_out_c_6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(158[24:70])
    defparam debug_uart_txd_I_0_3_lut.init = 16'hcaca;
    LUT4 i15493_2_lut (.A(qspi_data_in[2]), .B(rst_reg_n), .Z(qspi_data_out_3__N_5[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(127[22:56])
    defparam i15493_2_lut.init = 16'h8888;
    LUT4 gnd_bdd_2_lut_28428 (.A(n31388), .B(rst_reg_n_adj_3274), .Z(n31389)) /* synthesis lut_function=(A (B)) */ ;
    defparam gnd_bdd_2_lut_28428.init = 16'h8888;
    LUT4 rst_reg_n_bdd_4_lut (.A(cycle[0]), .B(n18086), .C(clk_c_enable_36), 
         .D(instr_complete_N_1647), .Z(n31388)) /* synthesis lut_function=(!(A (B (C))+!A (((D)+!C)+!B))) */ ;
    defparam rst_reg_n_bdd_4_lut.init = 16'h2a6a;
    LUT4 i26584_4_lut (.A(led_out), .B(data_to_write[0]), .C(n31964), 
         .D(n28840), .Z(n29201)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam i26584_4_lut.init = 16'hacaa;
    LUT4 i3865_4_lut (.A(n27183), .B(n31717), .C(n31713), .D(n31977), 
         .Z(clk_c_enable_324)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;
    defparam i3865_4_lut.init = 16'heefc;
    LUT4 user_interrupt_0__N_2800_I_0_2_lut_rep_650_3_lut_4_lut (.A(n32003), 
         .B(n31967), .C(n31905), .D(n32033), .Z(n31855)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(253[38:70])
    defparam user_interrupt_0__N_2800_I_0_2_lut_rep_650_3_lut_4_lut.init = 16'h0080;
    PFUMX i27136 (.BLUT(n29751), .ALUT(n29752), .C0(rs2[3]), .Z(n84));
    LUT4 i4_4_lut (.A(n28968), .B(\gpio_out_func_sel[7] [3]), .C(gpio_out_sel[7]), 
         .D(n3), .Z(uo_out_c_7)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i4_4_lut.init = 16'h1000;
    tqvp_uart_tx_U1 i_debug_uart_tx (.cycle_counter({cycle_counter}), .clk_c(clk_c), 
            .clk_c_enable_376(clk_c_enable_376), .n6210(n6210), .n72({n30_adj_3289, 
            n33_adj_3276, n36, n39_adj_3277, n42, n45_adj_3291, n48_adj_3288, 
            n51_adj_3275, n54, n57, n60_adj_3284, n63, n66_adj_3285}), 
            .debug_uart_txd(debug_uart_txd), .clk_c_enable_445(clk_c_enable_445), 
            .fsm_state({Open_35, Open_36, Open_37, fsm_state[0]}), .n32013(n32013), 
            .debug_uart_tx_start(debug_uart_tx_start), .n31828(n31828), 
            .n26116(n26116), .rst_reg_n(rst_reg_n), .\data_to_write[7] (data_to_write[7]), 
            .next_bit(next_bit), .clk_c_enable_534(clk_c_enable_534), .n31961(n31961), 
            .\data_to_write[1] (data_to_write[1]), .\data_to_write[2] (data_to_write[2]), 
            .\data_to_write[3] (data_to_write[3]), .\data_to_write[0] (data_to_write[0]), 
            .\data_to_write[4] (data_to_write[4]), .\data_to_write[5] (data_to_write[5]), 
            .\data_to_write[6] (data_to_write[6]), .uart_txd_N_2974(uart_txd_N_2974)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(228[4] 236[3])
    LUT4 i26410_2_lut (.A(\gpio_out_func_sel[7] [4]), .B(\gpio_out_func_sel[7] [2]), 
         .Z(n28968)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26410_2_lut.init = 16'heeee;
    LUT4 i26822_2_lut_rep_556_4_lut (.A(pc[2]), .B(n31978), .C(debug_instr_valid), 
         .D(n4263), .Z(n31761)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(40[23:40])
    defparam i26822_2_lut_rep_556_4_lut.init = 16'h0035;
    sim_qspi_pmod i_qspi (.\addr[2] (addr_adj_3335[2]), .qspi_clk_N_56(qspi_clk_N_56), 
            .qspi_data_in({qspi_data_in}), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), .\addr[1] (addr_adj_3335[1]), 
            .VCC_net(VCC_net), .\addr[14] (addr_adj_3335[14]), .\addr_24__N_228[14] (addr_24__N_228[14]), 
            .\addr[13] (addr_adj_3335[13]), .\addr[12] (addr_adj_3335[12]), 
            .\addr[11] (addr_adj_3335[11]), .\addr[10] (addr_adj_3335[10]), 
            .\addr[9] (addr_adj_3335[9]), .\addr[8] (addr_adj_3335[8]), 
            .\addr[7] (addr_adj_3335[7]), .\addr[6] (addr_adj_3335[6]), 
            .\addr[5] (addr_adj_3335[5]), .\addr[4] (addr_adj_3335[4]), 
            .\addr[3] (addr_adj_3335[3]), .qspi_ram_a_select(qspi_ram_a_select), 
            .qspi_ram_b_select(qspi_ram_b_select), .\addr[0] (addr_adj_3335[0]), 
            .\addr_24__N_228[0] (addr_24__N_228[0]), .\writing_N_164[3] (writing_N_164[3]), 
            .GND_net(GND_net), .\addr_24__N_228[9] (addr_24__N_228[9]), 
            .\addr_24__N_228[7] (addr_24__N_228[7]), .\addr_24__N_228[8] (addr_24__N_228[8]), 
            .\addr_24__N_228[6] (addr_24__N_228[6]), .\addr_24__N_228[5] (addr_24__N_228[5]), 
            .\addr_24__N_228[4] (addr_24__N_228[4]), .\addr_24__N_228[3] (addr_24__N_228[3]), 
            .\addr_24__N_228[2] (addr_24__N_228[2]), .\addr_24__N_228[10] (addr_24__N_228[10]), 
            .\addr_24__N_228[11] (addr_24__N_228[11]), .\addr_24__N_228[12] (addr_24__N_228[12]), 
            .\addr_24__N_228[13] (addr_24__N_228[13]), .\addr_24__N_228[1] (addr_24__N_228[1]), 
            .n32031(n32031)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(42[19] 50[6])
    LUT4 i1_2_lut_adj_623 (.A(rst_reg_n), .B(next_fsm_state_3__N_3015[3]), 
         .Z(clk_c_enable_542)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(31[12:46])
    defparam i1_2_lut_adj_623.init = 16'h2222;
    LUT4 i5316_3_lut (.A(ui_in_c_1), .B(data_to_write[0]), .C(rst_reg_n), 
         .Z(n7884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(250[12] 255[8])
    defparam i5316_3_lut.init = 16'hcaca;
    PFUMX i28638 (.BLUT(n32103), .ALUT(n32104), .C0(is_writing), .Z(n32105));
    PFUMX i28636 (.BLUT(n32100), .ALUT(n32101), .C0(n1160), .Z(clk_c_enable_234));
    PFUMX i27132 (.BLUT(n8), .ALUT(n9), .C0(rs2[1]), .Z(n29749));
    PFUMX i27133 (.BLUT(n11), .ALUT(n12), .C0(rs2[1]), .Z(n29750));
    
endmodule
//
// Verilog Description of module \peripherals_min(CLOCK_MHZ=14) 
//

module \peripherals_min(CLOCK_MHZ=14)  (\peri_data_out[4] , clk_c, clk_c_enable_387, 
            \peri_data_out[3] , \peri_data_out[0] , \peri_data_out[2] , 
            \peri_data_out[1] , \gpio_out_func_sel[5] , clk_c_enable_445, 
            \data_to_write[2] , clk_c_enable_349, \data_to_write[4] , 
            data_out_hold, n31883, clk_c_enable_360, \data_to_write[3] , 
            \gpio_out_func_sel[3] , clk_c_enable_357, clk_c_enable_259, 
            \data_to_write[1] , clk_c_enable_273, \gpio_out_func_sel[7][3] , 
            n32035, n26282, \addr[6] , \addr[9] , n31934, n32034, 
            ui_in_sync, n32019, \gpio_out_func_sel[1][3] , \data_to_write[0] , 
            \addr[2] , \addr[3] , \gpio_out_func_sel[4][3] , \gpio_out_func_sel[7][4] , 
            \gpio_out_func_sel[7][2] , baud_divider, n31922, \gpio_out_func_sel[2][3] , 
            \uo_out_from_user_peri[1][5] , n32003, n26205, \gpio_out_func_sel[6][3] , 
            \gpio_out_func_sel[0][3] , data_ready_r, rst_reg_n, data_ready_r_N_2792, 
            \peri_data_out[12] , \peri_data_out[11] , \peri_data_out[10] , 
            \peri_data_out[9] , \peri_data_out[8] , \peri_data_out[7] , 
            \peri_data_out[6] , \peri_data_out[5] , led_out, \addr[10] , 
            \addr[4] , \addr[8] , n4, n28840, \uo_out_from_user_peri[1][3] , 
            \data_to_write[5] , \data_to_write[6] , \data_to_write[7] , 
            \addr[7] , n31967, n32017, n8819, n31962, n31935, n18241, 
            n31936, \debug_rd_r[0] , debug_register_data, uo_out_c_2, 
            \debug_rd_r[1] , uo_out_c_3, \uo_out_from_user_peri[2][7] , 
            n26266, clk_c_enable_268, n31901, n80, n31900, n1, \debug_rd_r[2] , 
            uo_out_c_4, \peri_out[6] , n3, uo_out_c_0, uo_out_c_1, 
            clk_c_enable_542, clk_c_enable_390, clk_c_enable_395, \data_to_write[8] , 
            \data_to_write[9] , \data_to_write[10] , \data_to_write[11] , 
            \data_to_write[12] , \next_fsm_state_3__N_3015[3] , n27347, 
            n31932, n26116, n26216, n31905, n32033, n31929, \imm[6] , 
            \csr_read_3__N_1447[2] , n29162, cycle_counter, n72, fsm_state, 
            n31855, next_bit, n31963, fsm_state_adj_72, next_bit_adj_56, 
            cycle_counter_adj_73, n28760, GND_net, VCC_net, n31902, 
            n31925, n31923, next_bit_adj_70, n31828, uart_txd_N_2974, 
            clk_c_enable_534, debug_stop_txn, instr_active_N_2106, n32013, 
            \fsm_state[0]_adj_71 , clk_c_enable_376, n28686, n31880, 
            clk_c_enable_355, n1084, stop_txn_reg, stop_txn_now_N_2363, 
            clk_c_enable_239, n31971, n33479, \qspi_data_in[1] , n31593, 
            n31927, n27620, n31906, n27081, n6210, n31819, n28800, 
            n32027, clk_c_enable_531, n31950, n31977, n8135, n10499, 
            n10500, clk_c_enable_186, n32021, n31997, \addr[27] , 
            n31930, n32022, n31958, n26036, instr_complete_N_1647, 
            n28276, n31717, n29201) /* synthesis syn_module_defined=1 */ ;
    output \peri_data_out[4] ;
    input clk_c;
    input clk_c_enable_387;
    output \peri_data_out[3] ;
    output \peri_data_out[0] ;
    output \peri_data_out[2] ;
    output \peri_data_out[1] ;
    output [4:0]\gpio_out_func_sel[5] ;
    output clk_c_enable_445;
    input \data_to_write[2] ;
    input clk_c_enable_349;
    input \data_to_write[4] ;
    output data_out_hold;
    input n31883;
    input clk_c_enable_360;
    input \data_to_write[3] ;
    output [4:0]\gpio_out_func_sel[3] ;
    input clk_c_enable_357;
    input clk_c_enable_259;
    input \data_to_write[1] ;
    input clk_c_enable_273;
    output \gpio_out_func_sel[7][3] ;
    input n32035;
    output n26282;
    input \addr[6] ;
    input \addr[9] ;
    output n31934;
    input n32034;
    input [7:0]ui_in_sync;
    input n32019;
    output \gpio_out_func_sel[1][3] ;
    input \data_to_write[0] ;
    input \addr[2] ;
    input \addr[3] ;
    output \gpio_out_func_sel[4][3] ;
    output \gpio_out_func_sel[7][4] ;
    output \gpio_out_func_sel[7][2] ;
    output [12:0]baud_divider;
    output n31922;
    output \gpio_out_func_sel[2][3] ;
    output \uo_out_from_user_peri[1][5] ;
    output n32003;
    input n26205;
    output \gpio_out_func_sel[6][3] ;
    output \gpio_out_func_sel[0][3] ;
    output data_ready_r;
    input rst_reg_n;
    input data_ready_r_N_2792;
    output \peri_data_out[12] ;
    output \peri_data_out[11] ;
    output \peri_data_out[10] ;
    output \peri_data_out[9] ;
    output \peri_data_out[8] ;
    output \peri_data_out[7] ;
    output \peri_data_out[6] ;
    output \peri_data_out[5] ;
    output led_out;
    input \addr[10] ;
    input \addr[4] ;
    input \addr[8] ;
    output n4;
    output n28840;
    output \uo_out_from_user_peri[1][3] ;
    input \data_to_write[5] ;
    input \data_to_write[6] ;
    input \data_to_write[7] ;
    input \addr[7] ;
    input n31967;
    output n32017;
    output n8819;
    input n31962;
    input n31935;
    output n18241;
    input n31936;
    input \debug_rd_r[0] ;
    input debug_register_data;
    output uo_out_c_2;
    input \debug_rd_r[1] ;
    output uo_out_c_3;
    output \uo_out_from_user_peri[2][7] ;
    input n26266;
    input clk_c_enable_268;
    input n31901;
    input n80;
    input n31900;
    input n1;
    input \debug_rd_r[2] ;
    output uo_out_c_4;
    output \peri_out[6] ;
    output n3;
    output uo_out_c_0;
    output uo_out_c_1;
    input clk_c_enable_542;
    input clk_c_enable_390;
    input clk_c_enable_395;
    input \data_to_write[8] ;
    input \data_to_write[9] ;
    input \data_to_write[10] ;
    input \data_to_write[11] ;
    input \data_to_write[12] ;
    output \next_fsm_state_3__N_3015[3] ;
    input n27347;
    input n31932;
    input n26116;
    input n26216;
    output n31905;
    input n32033;
    input n31929;
    input \imm[6] ;
    input \csr_read_3__N_1447[2] ;
    output n29162;
    output [12:0]cycle_counter;
    input [12:0]n72;
    output [3:0]fsm_state;
    input n31855;
    input next_bit;
    input n31963;
    output [3:0]fsm_state_adj_72;
    input next_bit_adj_56;
    output [12:0]cycle_counter_adj_73;
    input n28760;
    input GND_net;
    input VCC_net;
    input n31902;
    input n31925;
    input n31923;
    input next_bit_adj_70;
    input n31828;
    input uart_txd_N_2974;
    output clk_c_enable_534;
    input debug_stop_txn;
    output instr_active_N_2106;
    input n32013;
    input \fsm_state[0]_adj_71 ;
    output clk_c_enable_376;
    input n28686;
    input n31880;
    output clk_c_enable_355;
    input n1084;
    input stop_txn_reg;
    input stop_txn_now_N_2363;
    output clk_c_enable_239;
    input n31971;
    input n33479;
    input \qspi_data_in[1] ;
    output n31593;
    input n31927;
    input n27620;
    input n31906;
    output n27081;
    output n6210;
    input n31819;
    input n28800;
    input n32027;
    output clk_c_enable_531;
    output n31950;
    input n31977;
    output n8135;
    input n10499;
    output n10500;
    output clk_c_enable_186;
    input n32021;
    input n31997;
    input \addr[27] ;
    output n31930;
    input n32022;
    input n31958;
    output n26036;
    input instr_complete_N_1647;
    input n28276;
    output n31717;
    input n29201;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n6052;
    wire [31:0]data_from_peri_31__N_2415;
    wire [4:0]\gpio_out_func_sel[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    
    wire clk_c_enable_10, n8695, clk_c_enable_352, clk_c_enable_356;
    wire [4:0]\gpio_out_func_sel[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    
    wire clk_c_enable_359;
    wire [4:0]\gpio_out_func_sel[6] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    
    wire clk_c_enable_115;
    wire [4:0]\gpio_out_func_sel[0] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    wire [4:0]\gpio_out_func_sel[4] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    wire [4:0]\gpio_out_func_sel[7] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    
    wire clk_c_enable_223, n8005;
    wire [31:0]data_from_user_peri_1__31__N_2455;
    
    wire n10;
    wire [7:0]\uo_out_from_user_peri[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(59[17:38])
    
    wire clk_c_enable_469, n3_c, n18493;
    wire [4:0]\gpio_out_func_sel[3]_c ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(119[15:32])
    
    wire clk_c_enable_275;
    wire [7:0]uart_rx_buf_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(98[15:31])
    
    wire n2, n1_c, n2_adj_3221, n1_adj_3222, n2_adj_3223, n1_adj_3224, 
        n29626, n29625, n2_adj_3225, n29624, n29623, n1_adj_3226, 
        n2_adj_3227, n2_adj_3228, n1_adj_3229, n1_adj_3230, clk_c_enable_334, 
        clk_c_enable_344, n31, n29, n28742, n27316, n29619, n29618, 
        n29617, n29616, clk_c_enable_377, clk_c_enable_378, clk_c_enable_386, 
        n30982;
    wire [7:0]\uo_out_from_user_peri[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(59[17:38])
    
    wire n30981, n29145, n29144, n29142, n29141, n29778, n29777, 
        n29779, n29780, n29781, n29776, n29775, n29146, n29143;
    wire [4:0]n1371;
    
    wire n25, n27413, n29170, n29620, n29621, n29622, n29627, 
        n29628, n29629, n31476, n27366, n3_adj_3231, n3_adj_3232, 
        n3_adj_3233, n3_adj_3234, n3_adj_3235, n3_adj_3236, n3_adj_3237, 
        clk_c_enable_185, clk_c_enable_35, n30983, n27437, n12, n27432, 
        n10_adj_3238, n27057, n28782, n27401, n9, n3_adj_3240, n3_adj_3242;
    
    FD1P3IX data_out_r__i4 (.D(data_from_peri_31__N_2415[4]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i4.GSR = "DISABLED";
    FD1P3IX data_out_r__i3 (.D(data_from_peri_31__N_2415[3]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i3.GSR = "DISABLED";
    FD1P3IX data_out_r__i0 (.D(data_from_peri_31__N_2415[0]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i0.GSR = "DISABLED";
    FD1P3IX data_out_r__i2 (.D(data_from_peri_31__N_2415[2]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i2.GSR = "DISABLED";
    FD1P3IX data_out_r__i1 (.D(data_from_peri_31__N_2415[1]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[1] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i1.GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_1[[1__362  (.D(n8695), .SP(clk_c_enable_10), 
            .CK(clk_c), .Q(\gpio_out_func_sel[1] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_1[[1__362 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_5[[2__381  (.D(\data_to_write[2] ), .SP(clk_c_enable_352), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[5] [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_5[[2__381 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_1[[2__361  (.D(\data_to_write[2] ), .SP(clk_c_enable_356), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[1] [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_1[[2__361 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_2[[2__366  (.D(\data_to_write[2] ), .SP(clk_c_enable_359), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[2] [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_2[[2__366 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_6[[4__384  (.D(\data_to_write[4] ), .SP(clk_c_enable_349), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[6] [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_6[[4__384 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_2[[4__364  (.D(\data_to_write[4] ), .SP(clk_c_enable_359), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[2] [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_2[[4__364 .GSR = "DISABLED";
    FD1P3IX data_out_hold_350 (.D(n31883), .SP(clk_c_enable_115), .CD(clk_c_enable_445), 
            .CK(clk_c), .Q(data_out_hold)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_hold_350.GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_0[[2__356  (.D(\data_to_write[2] ), .SP(clk_c_enable_360), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[0] [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_0[[2__356 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_5[[3__380  (.D(\data_to_write[3] ), .SP(clk_c_enable_352), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[5] [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_5[[3__380 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_3[[3__370  (.D(\data_to_write[3] ), .SP(clk_c_enable_357), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[3] [3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_3[[3__370 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_4[[1__377  (.D(\data_to_write[1] ), .SP(clk_c_enable_259), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[4] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_4[[1__377 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_0[[4__354  (.D(\data_to_write[4] ), .SP(clk_c_enable_360), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[0] [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_0[[4__354 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_7[[1__392  (.D(\data_to_write[1] ), .SP(clk_c_enable_273), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[7] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_7[[1__392 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_7[[3__390  (.D(\data_to_write[3] ), .SP(clk_c_enable_273), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[7][3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_7[[3__390 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_4[[2__376  (.D(\data_to_write[2] ), .SP(clk_c_enable_259), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[4] [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_4[[2__376 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_5[[1__382  (.D(\data_to_write[1] ), .SP(clk_c_enable_352), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[5] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_5[[1__382 .GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_4[[0__378  (.D(n8005), .SP(clk_c_enable_223), 
            .CK(clk_c), .Q(\gpio_out_func_sel[4] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_4[[0__378 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_4[[4__374  (.D(\data_to_write[4] ), .SP(clk_c_enable_259), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[4] [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_4[[4__374 .GSR = "DISABLED";
    LUT4 i1_2_lut_rep_729_4_lut (.A(n32035), .B(n26282), .C(\addr[6] ), 
         .D(\addr[9] ), .Z(n31934)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(133[45:67])
    defparam i1_2_lut_rep_729_4_lut.init = 16'hfffe;
    LUT4 i15550_2_lut_3_lut_4_lut (.A(n32035), .B(n32034), .C(ui_in_sync[7]), 
         .D(n32019), .Z(data_from_user_peri_1__31__N_2455[7])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15550_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n32035), .B(n32034), .C(ui_in_sync[5]), 
         .D(n32019), .Z(n10)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    FD1P3IX \gpio_out_func_sel_1[[3__360  (.D(\data_to_write[3] ), .SP(clk_c_enable_356), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[1][3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_1[[3__360 .GSR = "DISABLED";
    FD1P3IX gpio_out__i0 (.D(\data_to_write[0] ), .SP(clk_c_enable_469), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\uo_out_from_user_peri[1] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(122[12] 130[8])
    defparam gpio_out__i0.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_589 (.A(n32035), .B(n32034), .C(\addr[2] ), 
         .D(\addr[3] ), .Z(n3_c)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i1_2_lut_3_lut_4_lut_adj_589.init = 16'h1000;
    LUT4 i15551_2_lut_3_lut_4_lut (.A(n32035), .B(n32034), .C(ui_in_sync[6]), 
         .D(n32019), .Z(data_from_user_peri_1__31__N_2455[6])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15551_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i27865_3_lut_4_lut (.A(n32035), .B(n32034), .C(\addr[6] ), .D(\addr[2] ), 
         .Z(n18493)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i27865_3_lut_4_lut.init = 16'h0001;
    FD1P3IX \gpio_out_func_sel_3[[2__371  (.D(\data_to_write[2] ), .SP(clk_c_enable_357), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[3]_c [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_3[[2__371 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_6[[1__387  (.D(\data_to_write[1] ), .SP(clk_c_enable_349), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[6] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_6[[1__387 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_4[[3__375  (.D(\data_to_write[3] ), .SP(clk_c_enable_259), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[4][3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_4[[3__375 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_1[[4__359  (.D(\data_to_write[4] ), .SP(clk_c_enable_356), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[1] [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_1[[4__359 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_7[[4__389  (.D(\data_to_write[4] ), .SP(clk_c_enable_273), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[7][4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_7[[4__389 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_7[[2__391  (.D(\data_to_write[2] ), .SP(clk_c_enable_273), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[7][2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_7[[2__391 .GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_3[[0__373  (.D(n8005), .SP(clk_c_enable_275), 
            .CK(clk_c), .Q(\gpio_out_func_sel[3]_c [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_3[[0__373 .GSR = "DISABLED";
    LUT4 i15926_4_lut (.A(uart_rx_buf_data[7]), .B(n18493), .C(baud_divider[7]), 
         .D(\addr[3] ), .Z(n2)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15926_4_lut.init = 16'hc088;
    LUT4 i15441_4_lut (.A(\uo_out_from_user_peri[1] [7]), .B(\addr[6] ), 
         .C(data_from_user_peri_1__31__N_2455[7]), .D(n31922), .Z(n1_c)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15441_4_lut.init = 16'hc088;
    FD1P3IX \gpio_out_func_sel_6[[2__386  (.D(\data_to_write[2] ), .SP(clk_c_enable_349), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[6] [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_6[[2__386 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_0[[0__358  (.D(\data_to_write[0] ), .SP(clk_c_enable_360), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[0] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_0[[0__358 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_2[[3__365  (.D(\data_to_write[3] ), .SP(clk_c_enable_359), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[2][3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_2[[3__365 .GSR = "DISABLED";
    LUT4 i15927_4_lut (.A(uart_rx_buf_data[6]), .B(n18493), .C(baud_divider[6]), 
         .D(\addr[3] ), .Z(n2_adj_3221)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15927_4_lut.init = 16'hc088;
    LUT4 i15444_4_lut (.A(\uo_out_from_user_peri[1] [6]), .B(\addr[6] ), 
         .C(data_from_user_peri_1__31__N_2455[6]), .D(n31922), .Z(n1_adj_3222)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15444_4_lut.init = 16'hc088;
    LUT4 i15928_4_lut (.A(uart_rx_buf_data[5]), .B(n18493), .C(baud_divider[5]), 
         .D(\addr[3] ), .Z(n2_adj_3223)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15928_4_lut.init = 16'hc088;
    LUT4 i15445_4_lut (.A(\uo_out_from_user_peri[1][5] ), .B(\addr[6] ), 
         .C(n10), .D(n31922), .Z(n1_adj_3224)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15445_4_lut.init = 16'hc088;
    LUT4 i27009_3_lut (.A(\gpio_out_func_sel[6] [1]), .B(\gpio_out_func_sel[7] [1]), 
         .C(\addr[2] ), .Z(n29626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27009_3_lut.init = 16'hcaca;
    LUT4 i27008_3_lut (.A(\gpio_out_func_sel[4] [1]), .B(\gpio_out_func_sel[5] [1]), 
         .C(\addr[2] ), .Z(n29625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27008_3_lut.init = 16'hcaca;
    LUT4 i15929_4_lut (.A(uart_rx_buf_data[4]), .B(n18493), .C(baud_divider[4]), 
         .D(\addr[3] ), .Z(n2_adj_3225)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15929_4_lut.init = 16'hc088;
    LUT4 i27007_3_lut (.A(\gpio_out_func_sel[2] [1]), .B(\gpio_out_func_sel[3]_c [1]), 
         .C(\addr[2] ), .Z(n29624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27007_3_lut.init = 16'hcaca;
    LUT4 i27006_3_lut (.A(\gpio_out_func_sel[0] [1]), .B(\gpio_out_func_sel[1] [1]), 
         .C(\addr[2] ), .Z(n29623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27006_3_lut.init = 16'hcaca;
    LUT4 i15446_4_lut (.A(\uo_out_from_user_peri[1] [4]), .B(\addr[6] ), 
         .C(data_from_user_peri_1__31__N_2455[4]), .D(n31922), .Z(n1_adj_3226)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15446_4_lut.init = 16'hc088;
    LUT4 i15930_4_lut (.A(uart_rx_buf_data[3]), .B(n18493), .C(baud_divider[3]), 
         .D(\addr[3] ), .Z(n2_adj_3227)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15930_4_lut.init = 16'hc088;
    LUT4 i15931_4_lut (.A(uart_rx_buf_data[2]), .B(n18493), .C(baud_divider[2]), 
         .D(\addr[3] ), .Z(n2_adj_3228)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15931_4_lut.init = 16'hc088;
    LUT4 i15447_4_lut (.A(\uo_out_from_user_peri[1] [2]), .B(\addr[6] ), 
         .C(data_from_user_peri_1__31__N_2455[2]), .D(n31922), .Z(n1_adj_3229)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15447_4_lut.init = 16'hc088;
    LUT4 i15448_4_lut (.A(\uo_out_from_user_peri[1] [1]), .B(\addr[6] ), 
         .C(data_from_user_peri_1__31__N_2455[1]), .D(n31922), .Z(n1_adj_3230)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15448_4_lut.init = 16'hc088;
    FD1P3AX \gpio_out_func_sel_5[[0__383  (.D(n8005), .SP(clk_c_enable_334), 
            .CK(clk_c), .Q(\gpio_out_func_sel[5] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_5[[0__383 .GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_7[[0__393  (.D(n8005), .SP(clk_c_enable_344), 
            .CK(clk_c), .Q(\gpio_out_func_sel[7] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_7[[0__393 .GSR = "DISABLED";
    LUT4 i1_4_lut (.A(\addr[9] ), .B(\uo_out_from_user_peri[1] [0]), .C(n31), 
         .D(n31922), .Z(n29)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i1_4_lut.init = 16'h5044;
    LUT4 i1_4_lut_adj_590 (.A(n32003), .B(n26205), .C(n32035), .D(n28742), 
         .Z(n27316)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_590.init = 16'h0800;
    FD1P3IX \gpio_out_func_sel_6[[3__385  (.D(\data_to_write[3] ), .SP(clk_c_enable_349), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[6][3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_6[[3__385 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_3[[1__372  (.D(\data_to_write[1] ), .SP(clk_c_enable_357), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[3]_c [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_3[[1__372 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_5[[4__379  (.D(\data_to_write[4] ), .SP(clk_c_enable_352), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[5] [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_5[[4__379 .GSR = "DISABLED";
    LUT4 i27002_3_lut (.A(\gpio_out_func_sel[6] [4]), .B(\gpio_out_func_sel[7][4] ), 
         .C(\addr[2] ), .Z(n29619)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27002_3_lut.init = 16'hcaca;
    LUT4 i27001_3_lut (.A(\gpio_out_func_sel[4] [4]), .B(\gpio_out_func_sel[5] [4]), 
         .C(\addr[2] ), .Z(n29618)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27001_3_lut.init = 16'hcaca;
    LUT4 i27000_3_lut (.A(\gpio_out_func_sel[2] [4]), .B(\gpio_out_func_sel[3]_c [4]), 
         .C(\addr[2] ), .Z(n29617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27000_3_lut.init = 16'hcaca;
    LUT4 i26999_3_lut (.A(\gpio_out_func_sel[0] [4]), .B(\gpio_out_func_sel[1] [4]), 
         .C(\addr[2] ), .Z(n29616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26999_3_lut.init = 16'hcaca;
    FD1P3IX \gpio_out_func_sel_1[[0__363  (.D(\data_to_write[0] ), .SP(clk_c_enable_356), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[1] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_1[[0__363 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_3[[4__369  (.D(\data_to_write[4] ), .SP(clk_c_enable_357), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[3]_c [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_3[[4__369 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_2[[1__367  (.D(\data_to_write[1] ), .SP(clk_c_enable_359), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[2] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_2[[1__367 .GSR = "DISABLED";
    FD1P3IX \gpio_out_func_sel_0[[3__355  (.D(\data_to_write[3] ), .SP(clk_c_enable_360), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\gpio_out_func_sel[0][3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_0[[3__355 .GSR = "DISABLED";
    FD1P3AX data_ready_r_352 (.D(data_ready_r_N_2792), .SP(rst_reg_n), .CK(clk_c), 
            .Q(data_ready_r)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_ready_r_352.GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_0[[1__357  (.D(n8695), .SP(clk_c_enable_377), 
            .CK(clk_c), .Q(\gpio_out_func_sel[0] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_0[[1__357 .GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_2[[0__368  (.D(n8005), .SP(clk_c_enable_378), 
            .CK(clk_c), .Q(\gpio_out_func_sel[2] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_2[[0__368 .GSR = "DISABLED";
    FD1P3IX data_out_r__i12 (.D(data_from_peri_31__N_2415[12]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[12] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i12.GSR = "DISABLED";
    FD1P3IX data_out_r__i11 (.D(data_from_peri_31__N_2415[11]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[11] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i11.GSR = "DISABLED";
    FD1P3IX data_out_r__i10 (.D(data_from_peri_31__N_2415[10]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i10.GSR = "DISABLED";
    FD1P3IX data_out_r__i9 (.D(data_from_peri_31__N_2415[9]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[9] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i9.GSR = "DISABLED";
    FD1P3IX data_out_r__i8 (.D(data_from_peri_31__N_2415[8]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[8] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i8.GSR = "DISABLED";
    FD1P3IX data_out_r__i7 (.D(data_from_peri_31__N_2415[7]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[7] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i7.GSR = "DISABLED";
    FD1P3IX data_out_r__i6 (.D(data_from_peri_31__N_2415[6]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i6.GSR = "DISABLED";
    FD1P3AX \gpio_out_func_sel_6[[0__388  (.D(n8005), .SP(clk_c_enable_386), 
            .CK(clk_c), .Q(\gpio_out_func_sel[6] [0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam \gpio_out_func_sel_6[[0__388 .GSR = "DISABLED";
    FD1P3IX data_out_r__i5 (.D(data_from_peri_31__N_2415[5]), .SP(clk_c_enable_387), 
            .CD(n6052), .CK(clk_c), .Q(\peri_data_out[5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(68[12] 82[8])
    defparam data_out_r__i5.GSR = "DISABLED";
    LUT4 \uo_out_from_user_peri_2[[6__bdd_4_lut_28734  (.A(led_out), .B(\uo_out_from_user_peri[1] [0]), 
         .C(\gpio_out_func_sel[0] [0]), .D(\gpio_out_func_sel[0][3] ), .Z(n30982)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam \uo_out_from_user_peri_2[[6__bdd_4_lut_28734 .init = 16'h05c0;
    LUT4 \uo_out_from_user_peri_2[[6__bdd_3_lut  (.A(\uo_out_from_user_peri[2] [6]), 
         .B(\gpio_out_func_sel[0] [0]), .C(\gpio_out_func_sel[0][3] ), .Z(n30981)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam \uo_out_from_user_peri_2[[6__bdd_3_lut .init = 16'h0202;
    LUT4 i26528_3_lut (.A(\gpio_out_func_sel[1] [2]), .B(\gpio_out_func_sel[3]_c [2]), 
         .C(\addr[3] ), .Z(n29145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26528_3_lut.init = 16'hcaca;
    LUT4 i26527_3_lut (.A(\gpio_out_func_sel[0] [2]), .B(\gpio_out_func_sel[2] [2]), 
         .C(\addr[3] ), .Z(n29144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26527_3_lut.init = 16'hcaca;
    LUT4 i26525_3_lut (.A(\gpio_out_func_sel[6] [2]), .B(\gpio_out_func_sel[7][2] ), 
         .C(\addr[2] ), .Z(n29142)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26525_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_591 (.A(rst_reg_n), .B(n26205), .C(data_out_hold), 
         .D(\addr[10] ), .Z(n6052)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(71[18] 81[12])
    defparam i1_4_lut_adj_591.init = 16'h0800;
    LUT4 i26524_3_lut (.A(\gpio_out_func_sel[4] [2]), .B(\gpio_out_func_sel[5] [2]), 
         .C(\addr[2] ), .Z(n29141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26524_3_lut.init = 16'hcaca;
    LUT4 i27161_3_lut (.A(\gpio_out_func_sel[6] [0]), .B(\gpio_out_func_sel[7] [0]), 
         .C(\addr[2] ), .Z(n29778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27161_3_lut.init = 16'hcaca;
    LUT4 i27160_3_lut (.A(\gpio_out_func_sel[4] [0]), .B(\gpio_out_func_sel[5] [0]), 
         .C(\addr[2] ), .Z(n29777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27160_3_lut.init = 16'hcaca;
    L6MUX21 i27164 (.D0(n29779), .D1(n29780), .SD(\addr[4] ), .Z(n29781));
    LUT4 i27159_3_lut (.A(\gpio_out_func_sel[2] [0]), .B(\gpio_out_func_sel[3]_c [0]), 
         .C(\addr[2] ), .Z(n29776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27159_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(\addr[8] ), .B(\addr[6] ), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(106[13:36])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i27158_3_lut (.A(\gpio_out_func_sel[0] [0]), .B(\gpio_out_func_sel[1] [0]), 
         .C(\addr[2] ), .Z(n29775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27158_3_lut.init = 16'hcaca;
    LUT4 i27909_2_lut_rep_798 (.A(\addr[2] ), .B(\addr[3] ), .Z(n32003)) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i27909_2_lut_rep_798.init = 16'h1111;
    LUT4 i1_2_lut_rep_717_3_lut_4_lut (.A(\addr[2] ), .B(\addr[3] ), .C(n32034), 
         .D(n32035), .Z(n31922)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i1_2_lut_rep_717_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut (.A(\addr[2] ), .B(\addr[3] ), .C(\addr[9] ), 
         .Z(n28840)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i1_2_lut_3_lut.init = 16'h1010;
    FD1P3IX gpio_out__i1 (.D(\data_to_write[1] ), .SP(clk_c_enable_469), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\uo_out_from_user_peri[1] [1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(122[12] 130[8])
    defparam gpio_out__i1.GSR = "DISABLED";
    FD1P3IX gpio_out__i2 (.D(\data_to_write[2] ), .SP(clk_c_enable_469), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\uo_out_from_user_peri[1] [2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(122[12] 130[8])
    defparam gpio_out__i2.GSR = "DISABLED";
    FD1P3IX gpio_out__i3 (.D(\data_to_write[3] ), .SP(clk_c_enable_469), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\uo_out_from_user_peri[1][3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(122[12] 130[8])
    defparam gpio_out__i3.GSR = "DISABLED";
    FD1P3IX gpio_out__i4 (.D(\data_to_write[4] ), .SP(clk_c_enable_469), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\uo_out_from_user_peri[1] [4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(122[12] 130[8])
    defparam gpio_out__i4.GSR = "DISABLED";
    FD1P3IX gpio_out__i5 (.D(\data_to_write[5] ), .SP(clk_c_enable_469), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\uo_out_from_user_peri[1][5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(122[12] 130[8])
    defparam gpio_out__i5.GSR = "DISABLED";
    FD1P3IX gpio_out__i6 (.D(\data_to_write[6] ), .SP(clk_c_enable_469), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\uo_out_from_user_peri[1] [6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(122[12] 130[8])
    defparam gpio_out__i6.GSR = "DISABLED";
    FD1P3IX gpio_out__i7 (.D(\data_to_write[7] ), .SP(clk_c_enable_469), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(\uo_out_from_user_peri[1] [7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(122[12] 130[8])
    defparam gpio_out__i7.GSR = "DISABLED";
    L6MUX21 mux_74_Mux_2_i7 (.D0(n29146), .D1(n29143), .SD(\addr[4] ), 
            .Z(n1371[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    LUT4 i15220_4_lut (.A(n25), .B(\addr[8] ), .C(n27413), .D(\addr[7] ), 
         .Z(data_from_peri_31__N_2415[0])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15220_4_lut.init = 16'h3022;
    LUT4 i1_4_lut_adj_592 (.A(n29170), .B(n31967), .C(\addr[6] ), .D(\addr[9] ), 
         .Z(n27413)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_592.init = 16'h0008;
    L6MUX21 i27005 (.D0(n29620), .D1(n29621), .SD(\addr[4] ), .Z(n29622));
    L6MUX21 i27012 (.D0(n29627), .D1(n29628), .SD(\addr[4] ), .Z(n29629));
    LUT4 i15562_2_lut_rep_812 (.A(\addr[6] ), .B(\addr[7] ), .Z(n32017)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(108[62:74])
    defparam i15562_2_lut_rep_812.init = 16'heeee;
    LUT4 i7117_2_lut_3_lut (.A(\addr[6] ), .B(\addr[7] ), .C(\addr[9] ), 
         .Z(n8819)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(108[62:74])
    defparam i7117_2_lut_3_lut.init = 16'h1e1e;
    LUT4 i1_3_lut_4_lut_4_lut (.A(\addr[6] ), .B(n31476), .C(n32034), 
         .D(n32035), .Z(n27366)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(106[13:36])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h0004;
    LUT4 i1_4_lut_adj_593 (.A(\addr[8] ), .B(\addr[10] ), .C(\addr[9] ), 
         .D(led_out), .Z(n28742)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_593.init = 16'h1000;
    LUT4 i49_4_lut (.A(ui_in_sync[0]), .B(n31962), .C(n31935), .D(n29781), 
         .Z(n31)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i49_4_lut.init = 16'h3a0a;
    LUT4 mux_3064_i2_4_lut (.A(ui_in_sync[1]), .B(n29629), .C(n31935), 
         .D(n31962), .Z(data_from_user_peri_1__31__N_2455[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(133[45] 135[50])
    defparam mux_3064_i2_4_lut.init = 16'h0aca;
    LUT4 mux_3064_i3_4_lut (.A(ui_in_sync[2]), .B(n1371[2]), .C(n31935), 
         .D(n31962), .Z(data_from_user_peri_1__31__N_2455[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(133[45] 135[50])
    defparam mux_3064_i3_4_lut.init = 16'h0aca;
    LUT4 mux_3064_i5_4_lut (.A(ui_in_sync[4]), .B(n29622), .C(n31935), 
         .D(n31962), .Z(data_from_user_peri_1__31__N_2455[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(133[45] 135[50])
    defparam mux_3064_i5_4_lut.init = 16'h0aca;
    LUT4 i15874_2_lut_3_lut (.A(\addr[8] ), .B(\addr[9] ), .C(n3_adj_3231), 
         .Z(data_from_peri_31__N_2415[7])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15874_2_lut_3_lut.init = 16'h1010;
    LUT4 i15885_2_lut_3_lut (.A(\addr[8] ), .B(\addr[9] ), .C(n3_adj_3232), 
         .Z(data_from_peri_31__N_2415[1])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15885_2_lut_3_lut.init = 16'h1010;
    LUT4 i15881_2_lut_3_lut (.A(\addr[8] ), .B(\addr[9] ), .C(n3_adj_3233), 
         .Z(data_from_peri_31__N_2415[2])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15881_2_lut_3_lut.init = 16'h1010;
    LUT4 i15877_2_lut_3_lut (.A(\addr[8] ), .B(\addr[9] ), .C(n3_adj_3234), 
         .Z(data_from_peri_31__N_2415[4])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15877_2_lut_3_lut.init = 16'h1010;
    LUT4 i15880_2_lut_3_lut (.A(\addr[8] ), .B(\addr[9] ), .C(n3_adj_3235), 
         .Z(data_from_peri_31__N_2415[3])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15880_2_lut_3_lut.init = 16'h1010;
    LUT4 i15875_2_lut_3_lut (.A(\addr[8] ), .B(\addr[9] ), .C(n3_adj_3236), 
         .Z(data_from_peri_31__N_2415[6])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15875_2_lut_3_lut.init = 16'h1010;
    LUT4 i15876_2_lut_3_lut (.A(\addr[8] ), .B(\addr[9] ), .C(n3_adj_3237), 
         .Z(data_from_peri_31__N_2415[5])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15876_2_lut_3_lut.init = 16'h1010;
    PFUMX i27162 (.BLUT(n29775), .ALUT(n29776), .C0(\addr[3] ), .Z(n29779));
    PFUMX i27163 (.BLUT(n29777), .ALUT(n29778), .C0(\addr[3] ), .Z(n29780));
    LUT4 i1_3_lut (.A(n26282), .B(\addr[6] ), .C(\addr[9] ), .Z(n18241)) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam i1_3_lut.init = 16'hfbfb;
    LUT4 i1_3_lut_adj_594 (.A(\addr[10] ), .B(\addr[7] ), .C(\addr[8] ), 
         .Z(n26282)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(106[13:36])
    defparam i1_3_lut_adj_594.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut (.A(n31936), .B(clk_c_enable_185), .C(\addr[2] ), 
         .D(rst_reg_n), .Z(clk_c_enable_35)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h04ff;
    PFUMX i26526 (.BLUT(n29141), .ALUT(n29142), .C0(\addr[3] ), .Z(n29143));
    PFUMX i26529 (.BLUT(n29144), .ALUT(n29145), .C0(\addr[2] ), .Z(n29146));
    PFUMX i28182 (.BLUT(n30982), .ALUT(n30981), .C0(\gpio_out_func_sel[0] [1]), 
          .Z(n30983));
    LUT4 i25_3_lut (.A(n27437), .B(\debug_rd_r[0] ), .C(debug_register_data), 
         .Z(uo_out_c_2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(84[9:28])
    defparam i25_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(\gpio_out_func_sel[2][3] ), .B(\gpio_out_func_sel[2] [4]), 
         .C(n12), .D(\gpio_out_func_sel[2] [2]), .Z(n27437)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    LUT4 i26_4_lut (.A(\uo_out_from_user_peri[2] [6]), .B(\gpio_out_func_sel[2] [0]), 
         .C(\gpio_out_func_sel[2] [1]), .D(\uo_out_from_user_peri[1] [2]), 
         .Z(n12)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(84[9:28])
    defparam i26_4_lut.init = 16'h2c20;
    PFUMX i27003 (.BLUT(n29616), .ALUT(n29617), .C0(\addr[3] ), .Z(n29620));
    LUT4 i23_3_lut (.A(n27432), .B(\debug_rd_r[1] ), .C(debug_register_data), 
         .Z(uo_out_c_3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(84[9:28])
    defparam i23_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut_adj_595 (.A(\gpio_out_func_sel[3] [3]), .B(n10_adj_3238), 
         .C(\gpio_out_func_sel[3]_c [2]), .D(\gpio_out_func_sel[3]_c [4]), 
         .Z(n27432)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i3_4_lut_adj_595.init = 16'h0004;
    LUT4 i24_4_lut (.A(\uo_out_from_user_peri[1][3] ), .B(\uo_out_from_user_peri[2][7] ), 
         .C(\gpio_out_func_sel[3]_c [1]), .D(\gpio_out_func_sel[3]_c [0]), 
         .Z(n10_adj_3238)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(84[9:28])
    defparam i24_4_lut.init = 16'h0ac0;
    PFUMX i27004 (.BLUT(n29618), .ALUT(n29619), .C0(\addr[3] ), .Z(n29621));
    PFUMX i27010 (.BLUT(n29623), .ALUT(n29624), .C0(\addr[3] ), .Z(n29627));
    LUT4 i15946_2_lut (.A(baud_divider[12]), .B(n27057), .Z(data_from_peri_31__N_2415[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15946_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_596 (.A(n31967), .B(n26266), .C(n28782), .D(n4), 
         .Z(n27057)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_596.init = 16'hfffd;
    LUT4 i1_2_lut_adj_597 (.A(\addr[7] ), .B(\addr[9] ), .Z(n28782)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut_adj_597.init = 16'hdddd;
    LUT4 i15592_2_lut (.A(baud_divider[11]), .B(n27057), .Z(data_from_peri_31__N_2415[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15592_2_lut.init = 16'h2222;
    PFUMX i48 (.BLUT(n27316), .ALUT(n29), .C0(\addr[6] ), .Z(n25));
    LUT4 i15920_2_lut (.A(baud_divider[10]), .B(n27057), .Z(data_from_peri_31__N_2415[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15920_2_lut.init = 16'h2222;
    LUT4 i15923_2_lut (.A(baud_divider[9]), .B(n27057), .Z(data_from_peri_31__N_2415[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15923_2_lut.init = 16'h2222;
    LUT4 i15924_2_lut (.A(baud_divider[8]), .B(n27057), .Z(data_from_peri_31__N_2415[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(107[50:62])
    defparam i15924_2_lut.init = 16'h2222;
    PFUMX addr_in_9__I_0_542_Mux_1_i3 (.BLUT(n1_adj_3230), .ALUT(n27366), 
          .C0(\addr[7] ), .Z(n3_adj_3232)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    PFUMX addr_in_9__I_0_542_Mux_2_i3 (.BLUT(n1_adj_3229), .ALUT(n2_adj_3228), 
          .C0(\addr[7] ), .Z(n3_adj_3233)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    LUT4 i1_2_lut_4_lut_adj_598 (.A(clk_c_enable_268), .B(rst_reg_n), .C(n18241), 
         .D(n31901), .Z(clk_c_enable_359)) /* synthesis lut_function=(!((B (C+(D))+!B (D))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam i1_2_lut_4_lut_adj_598.init = 16'h002a;
    LUT4 i1_2_lut_4_lut_adj_599 (.A(clk_c_enable_268), .B(rst_reg_n), .C(n18241), 
         .D(n80), .Z(clk_c_enable_356)) /* synthesis lut_function=(!((B (C+(D))+!B (D))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam i1_2_lut_4_lut_adj_599.init = 16'h002a;
    LUT4 i1_2_lut_4_lut_adj_600 (.A(clk_c_enable_268), .B(rst_reg_n), .C(n18241), 
         .D(n31900), .Z(clk_c_enable_352)) /* synthesis lut_function=(!((B (C+(D))+!B (D))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(142[20] 150[16])
    defparam i1_2_lut_4_lut_adj_600.init = 16'h002a;
    PFUMX addr_in_9__I_0_542_Mux_3_i3 (.BLUT(n1), .ALUT(n2_adj_3227), .C0(\addr[7] ), 
          .Z(n3_adj_3235)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    LUT4 i22_3_lut (.A(n27401), .B(\debug_rd_r[2] ), .C(debug_register_data), 
         .Z(uo_out_c_4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(84[9:28])
    defparam i22_3_lut.init = 16'hcaca;
    PFUMX addr_in_9__I_0_542_Mux_4_i3 (.BLUT(n1_adj_3226), .ALUT(n2_adj_3225), 
          .C0(\addr[7] ), .Z(n3_adj_3234)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    LUT4 i3_4_lut_adj_601 (.A(\gpio_out_func_sel[4][3] ), .B(\gpio_out_func_sel[4] [4]), 
         .C(n9), .D(\gpio_out_func_sel[4] [2]), .Z(n27401)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_601.init = 16'h0010;
    LUT4 i23_4_lut (.A(\uo_out_from_user_peri[1] [4]), .B(\uo_out_from_user_peri[2] [6]), 
         .C(\gpio_out_func_sel[4] [1]), .D(\gpio_out_func_sel[4] [0]), .Z(n9)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(84[9:28])
    defparam i23_4_lut.init = 16'h0ac0;
    PFUMX i27011 (.BLUT(n29625), .ALUT(n29626), .C0(\addr[3] ), .Z(n29628));
    PFUMX addr_in_9__I_0_542_Mux_5_i3 (.BLUT(n1_adj_3224), .ALUT(n2_adj_3223), 
          .C0(\addr[7] ), .Z(n3_adj_3237)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    PFUMX addr_in_9__I_0_542_Mux_6_i3 (.BLUT(n1_adj_3222), .ALUT(n2_adj_3221), 
          .C0(\addr[7] ), .Z(n3_adj_3236)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    PFUMX addr_in_9__I_0_542_Mux_7_i3 (.BLUT(n1_c), .ALUT(n2), .C0(\addr[7] ), 
          .Z(n3_adj_3231)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=46, LSE_RCOL=6, LSE_LLINE=161, LSE_RLINE=180 */ ;
    LUT4 i3_4_lut_adj_602 (.A(n3_adj_3240), .B(\gpio_out_func_sel[6] [4]), 
         .C(\gpio_out_func_sel[6] [2]), .D(\gpio_out_func_sel[6][3] ), .Z(\peri_out[6] )) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut_adj_602.init = 16'h0002;
    LUT4 mux_239_Mux_0_i3_4_lut (.A(\uo_out_from_user_peri[1] [6]), .B(\uo_out_from_user_peri[2] [6]), 
         .C(\gpio_out_func_sel[6] [1]), .D(\gpio_out_func_sel[6] [0]), .Z(n3_adj_3240)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(156[62:87])
    defparam mux_239_Mux_0_i3_4_lut.init = 16'h0ac0;
    LUT4 mux_240_Mux_0_i3_4_lut (.A(\gpio_out_func_sel[7] [0]), .B(\uo_out_from_user_peri[2][7] ), 
         .C(\gpio_out_func_sel[7] [1]), .D(\uo_out_from_user_peri[1] [7]), 
         .Z(n3)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(156[62:87])
    defparam mux_240_Mux_0_i3_4_lut.init = 16'h4a40;
    LUT4 i2_3_lut (.A(\gpio_out_func_sel[0] [4]), .B(n30983), .C(\gpio_out_func_sel[0] [2]), 
         .Z(uo_out_c_0)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut.init = 16'h0404;
    LUT4 i3_4_lut_adj_603 (.A(n3_adj_3242), .B(\gpio_out_func_sel[1] [4]), 
         .C(\gpio_out_func_sel[1][3] ), .D(\gpio_out_func_sel[1] [2]), .Z(uo_out_c_1)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut_adj_603.init = 16'h0002;
    LUT4 mux_234_Mux_0_i3_4_lut (.A(\uo_out_from_user_peri[1] [1]), .B(\uo_out_from_user_peri[2][7] ), 
         .C(\gpio_out_func_sel[1] [1]), .D(\gpio_out_func_sel[1] [0]), .Z(n3_adj_3242)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(156[62:87])
    defparam mux_234_Mux_0_i3_4_lut.init = 16'h0ac0;
    \tqvp_uart_wrapper(CLOCK_MHZ=14)  i_uart (.baud_divider({baud_divider}), 
            .clk_c(clk_c), .clk_c_enable_35(clk_c_enable_35), .clk_c_enable_445(clk_c_enable_445), 
            .\data_to_write[6] (\data_to_write[6] ), .\data_to_write[5] (\data_to_write[5] ), 
            .\data_to_write[4] (\data_to_write[4] ), .\data_to_write[3] (\data_to_write[3] ), 
            .\data_to_write[0] (\data_to_write[0] ), .\addr[3] (\addr[3] ), 
            .n31476(n31476), .clk_c_enable_185(clk_c_enable_185), .\addr[2] (\addr[2] ), 
            .clk_c_enable_542(clk_c_enable_542), .clk_c_enable_390(clk_c_enable_390), 
            .\data_to_write[1] (\data_to_write[1] ), .\data_to_write[2] (\data_to_write[2] ), 
            .\data_to_write[7] (\data_to_write[7] ), .clk_c_enable_395(clk_c_enable_395), 
            .\data_to_write[8] (\data_to_write[8] ), .\data_to_write[9] (\data_to_write[9] ), 
            .\data_to_write[10] (\data_to_write[10] ), .\data_to_write[11] (\data_to_write[11] ), 
            .\data_to_write[12] (\data_to_write[12] ), .\ui_in_sync[7] (ui_in_sync[7]), 
            .\ui_in_sync[3] (ui_in_sync[3]), .\next_fsm_state_3__N_3015[3] (\next_fsm_state_3__N_3015[3] ), 
            .n27347(n27347), .\uart_rx_buf_data[2] (uart_rx_buf_data[2]), 
            .\uart_rx_buf_data[3] (uart_rx_buf_data[3]), .\uart_rx_buf_data[4] (uart_rx_buf_data[4]), 
            .\uart_rx_buf_data[5] (uart_rx_buf_data[5]), .\uart_rx_buf_data[6] (uart_rx_buf_data[6]), 
            .\uart_rx_buf_data[7] (uart_rx_buf_data[7]), .n31922(n31922), 
            .rst_reg_n(rst_reg_n), .n31932(n31932), .n26116(n26116), .\addr[9] (\addr[9] ), 
            .n26216(n26216), .\addr[10] (\addr[10] ), .n31905(n31905), 
            .n32033(n32033), .n31929(n31929), .\imm[6] (\imm[6] ), .\csr_read_3__N_1447[2] (\csr_read_3__N_1447[2] ), 
            .n29162(n29162), .n29170(n29170), .cycle_counter({cycle_counter}), 
            .n72({n72}), .fsm_state({fsm_state}), .\uo_out_from_user_peri[2][6] (\uo_out_from_user_peri[2] [6]), 
            .n31855(n31855), .next_bit(next_bit), .n31963(n31963), .fsm_state_adj_50({fsm_state_adj_72}), 
            .next_bit_adj_34(next_bit_adj_56), .cycle_counter_adj_51({cycle_counter_adj_73}), 
            .\uo_out_from_user_peri[2][7] (\uo_out_from_user_peri[2][7] ), 
            .n28760(n28760), .GND_net(GND_net), .VCC_net(VCC_net), .n31902(n31902), 
            .n31925(n31925), .n32003(n32003), .clk_c_enable_223(clk_c_enable_223), 
            .n31923(n31923), .\addr[4] (\addr[4] ), .clk_c_enable_275(clk_c_enable_275), 
            .next_bit_adj_48(next_bit_adj_70), .n31828(n31828), .uart_txd_N_2974(uart_txd_N_2974), 
            .clk_c_enable_534(clk_c_enable_534), .debug_stop_txn(debug_stop_txn), 
            .instr_active_N_2106(instr_active_N_2106), .clk_c_enable_344(clk_c_enable_344), 
            .n3(n3_c), .n32013(n32013), .\fsm_state[0]_adj_49 (\fsm_state[0]_adj_71 ), 
            .clk_c_enable_376(clk_c_enable_376), .n28686(n28686), .n31880(n31880), 
            .clk_c_enable_355(clk_c_enable_355), .n8005(n8005), .n1084(n1084), 
            .stop_txn_reg(stop_txn_reg), .stop_txn_now_N_2363(stop_txn_now_N_2363), 
            .clk_c_enable_239(clk_c_enable_239), .n31971(n31971), .n33479(n33479), 
            .\qspi_data_in[1] (\qspi_data_in[1] ), .n31593(n31593), .n26266(n26266), 
            .n31927(n31927), .clk_c_enable_378(clk_c_enable_378), .n27620(n27620), 
            .n31906(n31906), .n27081(n27081), .clk_c_enable_377(clk_c_enable_377), 
            .n6210(n6210), .n31819(n31819), .n28800(n28800), .n32027(n32027), 
            .n32034(n32034), .clk_c_enable_531(clk_c_enable_531), .n31950(n31950), 
            .n18241(n18241), .clk_c_enable_268(clk_c_enable_268), .clk_c_enable_469(clk_c_enable_469), 
            .clk_c_enable_386(clk_c_enable_386), .n8695(n8695), .n31977(n31977), 
            .n8135(n8135), .n10499(n10499), .n10500(n10500), .clk_c_enable_186(clk_c_enable_186), 
            .n32021(n32021), .n31997(n31997), .\addr[27] (\addr[27] ), 
            .n31930(n31930), .n32022(n32022), .n31958(n31958), .n26036(n26036), 
            .instr_complete_N_1647(instr_complete_N_1647), .n28276(n28276), 
            .n31883(n31883), .clk_c_enable_115(clk_c_enable_115), .n32019(n32019), 
            .clk_c_enable_334(clk_c_enable_334), .n31717(n31717), .n80(n80), 
            .clk_c_enable_10(clk_c_enable_10)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(190[45] 202[3])
    led i_led (.led_out(led_out), .clk_c(clk_c), .clk_c_enable_268(clk_c_enable_268), 
        .clk_c_enable_445(clk_c_enable_445), .n29201(n29201)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peripherals_min.v(217[6] 229[3])
    
endmodule
//
// Verilog Description of module \tqvp_uart_wrapper(CLOCK_MHZ=14) 
//

module \tqvp_uart_wrapper(CLOCK_MHZ=14)  (baud_divider, clk_c, clk_c_enable_35, 
            clk_c_enable_445, \data_to_write[6] , \data_to_write[5] , 
            \data_to_write[4] , \data_to_write[3] , \data_to_write[0] , 
            \addr[3] , n31476, clk_c_enable_185, \addr[2] , clk_c_enable_542, 
            clk_c_enable_390, \data_to_write[1] , \data_to_write[2] , 
            \data_to_write[7] , clk_c_enable_395, \data_to_write[8] , 
            \data_to_write[9] , \data_to_write[10] , \data_to_write[11] , 
            \data_to_write[12] , \ui_in_sync[7] , \ui_in_sync[3] , \next_fsm_state_3__N_3015[3] , 
            n27347, \uart_rx_buf_data[2] , \uart_rx_buf_data[3] , \uart_rx_buf_data[4] , 
            \uart_rx_buf_data[5] , \uart_rx_buf_data[6] , \uart_rx_buf_data[7] , 
            n31922, rst_reg_n, n31932, n26116, \addr[9] , n26216, 
            \addr[10] , n31905, n32033, n31929, \imm[6] , \csr_read_3__N_1447[2] , 
            n29162, n29170, cycle_counter, n72, fsm_state, \uo_out_from_user_peri[2][6] , 
            n31855, next_bit, n31963, fsm_state_adj_50, next_bit_adj_34, 
            cycle_counter_adj_51, \uo_out_from_user_peri[2][7] , n28760, 
            GND_net, VCC_net, n31902, n31925, n32003, clk_c_enable_223, 
            n31923, \addr[4] , clk_c_enable_275, next_bit_adj_48, n31828, 
            uart_txd_N_2974, clk_c_enable_534, debug_stop_txn, instr_active_N_2106, 
            clk_c_enable_344, n3, n32013, \fsm_state[0]_adj_49 , clk_c_enable_376, 
            n28686, n31880, clk_c_enable_355, n8005, n1084, stop_txn_reg, 
            stop_txn_now_N_2363, clk_c_enable_239, n31971, n33479, \qspi_data_in[1] , 
            n31593, n26266, n31927, clk_c_enable_378, n27620, n31906, 
            n27081, clk_c_enable_377, n6210, n31819, n28800, n32027, 
            n32034, clk_c_enable_531, n31950, n18241, clk_c_enable_268, 
            clk_c_enable_469, clk_c_enable_386, n8695, n31977, n8135, 
            n10499, n10500, clk_c_enable_186, n32021, n31997, \addr[27] , 
            n31930, n32022, n31958, n26036, instr_complete_N_1647, 
            n28276, n31883, clk_c_enable_115, n32019, clk_c_enable_334, 
            n31717, n80, clk_c_enable_10) /* synthesis syn_module_defined=1 */ ;
    output [12:0]baud_divider;
    input clk_c;
    input clk_c_enable_35;
    output clk_c_enable_445;
    input \data_to_write[6] ;
    input \data_to_write[5] ;
    input \data_to_write[4] ;
    input \data_to_write[3] ;
    input \data_to_write[0] ;
    input \addr[3] ;
    output n31476;
    output clk_c_enable_185;
    input \addr[2] ;
    input clk_c_enable_542;
    input clk_c_enable_390;
    input \data_to_write[1] ;
    input \data_to_write[2] ;
    input \data_to_write[7] ;
    input clk_c_enable_395;
    input \data_to_write[8] ;
    input \data_to_write[9] ;
    input \data_to_write[10] ;
    input \data_to_write[11] ;
    input \data_to_write[12] ;
    input \ui_in_sync[7] ;
    input \ui_in_sync[3] ;
    output \next_fsm_state_3__N_3015[3] ;
    input n27347;
    output \uart_rx_buf_data[2] ;
    output \uart_rx_buf_data[3] ;
    output \uart_rx_buf_data[4] ;
    output \uart_rx_buf_data[5] ;
    output \uart_rx_buf_data[6] ;
    output \uart_rx_buf_data[7] ;
    input n31922;
    input rst_reg_n;
    input n31932;
    input n26116;
    input \addr[9] ;
    input n26216;
    input \addr[10] ;
    output n31905;
    input n32033;
    input n31929;
    input \imm[6] ;
    input \csr_read_3__N_1447[2] ;
    output n29162;
    output n29170;
    output [12:0]cycle_counter;
    input [12:0]n72;
    output [3:0]fsm_state;
    output \uo_out_from_user_peri[2][6] ;
    input n31855;
    input next_bit;
    input n31963;
    output [3:0]fsm_state_adj_50;
    input next_bit_adj_34;
    output [12:0]cycle_counter_adj_51;
    output \uo_out_from_user_peri[2][7] ;
    input n28760;
    input GND_net;
    input VCC_net;
    input n31902;
    input n31925;
    input n32003;
    output clk_c_enable_223;
    input n31923;
    input \addr[4] ;
    output clk_c_enable_275;
    input next_bit_adj_48;
    input n31828;
    input uart_txd_N_2974;
    output clk_c_enable_534;
    input debug_stop_txn;
    output instr_active_N_2106;
    output clk_c_enable_344;
    input n3;
    input n32013;
    input \fsm_state[0]_adj_49 ;
    output clk_c_enable_376;
    input n28686;
    input n31880;
    output clk_c_enable_355;
    output n8005;
    input n1084;
    input stop_txn_reg;
    input stop_txn_now_N_2363;
    output clk_c_enable_239;
    input n31971;
    input n33479;
    input \qspi_data_in[1] ;
    output n31593;
    input n26266;
    input n31927;
    output clk_c_enable_378;
    input n27620;
    input n31906;
    output n27081;
    output clk_c_enable_377;
    output n6210;
    input n31819;
    input n28800;
    input n32027;
    input n32034;
    output clk_c_enable_531;
    output n31950;
    input n18241;
    input clk_c_enable_268;
    output clk_c_enable_469;
    output clk_c_enable_386;
    output n8695;
    input n31977;
    output n8135;
    input n10499;
    output n10500;
    output clk_c_enable_186;
    input n32021;
    input n31997;
    input \addr[27] ;
    output n31930;
    input n32022;
    input n31958;
    output n26036;
    input instr_complete_N_1647;
    input n28276;
    input n31883;
    output clk_c_enable_115;
    input n32019;
    output clk_c_enable_334;
    output n31717;
    input n80;
    output clk_c_enable_10;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n31475, n31474, rxd_select, n29200, n29169;
    wire [7:0]uart_rx_buf_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(98[15:31])
    wire [7:0]uart_rx_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(81[16:28])
    
    wire n32000, mid_bit;
    wire [3:0]next_fsm_state_3__N_3011;
    
    wire clk_c_enable_535, n31811, n9493, n26118, n29168, clk_c_enable_152, 
        n6158, clk_c_enable_525, n18596;
    
    FD1P3JX baud_divider_i6 (.D(\data_to_write[6] ), .SP(clk_c_enable_35), 
            .PD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[6])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i6.GSR = "DISABLED";
    FD1P3JX baud_divider_i5 (.D(\data_to_write[5] ), .SP(clk_c_enable_35), 
            .PD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[5])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i5.GSR = "DISABLED";
    FD1P3JX baud_divider_i4 (.D(\data_to_write[4] ), .SP(clk_c_enable_35), 
            .PD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[4])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i4.GSR = "DISABLED";
    FD1P3JX baud_divider_i3 (.D(\data_to_write[3] ), .SP(clk_c_enable_35), 
            .PD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[3])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i3.GSR = "DISABLED";
    FD1P3JX baud_divider_i0 (.D(\data_to_write[0] ), .SP(clk_c_enable_35), 
            .PD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[0])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i0.GSR = "DISABLED";
    PFUMX i28476 (.BLUT(n31475), .ALUT(n31474), .C0(\addr[3] ), .Z(n31476));
    FD1P3IX rxd_select_58 (.D(n29200), .SP(clk_c_enable_185), .CD(clk_c_enable_445), 
            .CK(clk_c), .Q(rxd_select)) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(50[12] 58[8])
    defparam rxd_select_58.GSR = "DISABLED";
    LUT4 i26552_3_lut (.A(baud_divider[0]), .B(rxd_select), .C(\addr[2] ), 
         .Z(n29169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26552_3_lut.init = 16'hcaca;
    FD1P3AX uart_rx_buf_data_i0_i0 (.D(uart_rx_data[0]), .SP(clk_c_enable_542), 
            .CK(clk_c), .Q(uart_rx_buf_data[0])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i0.GSR = "DISABLED";
    FD1P3IX baud_divider_i1 (.D(\data_to_write[1] ), .SP(clk_c_enable_390), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[1])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i1.GSR = "DISABLED";
    FD1P3IX baud_divider_i2 (.D(\data_to_write[2] ), .SP(clk_c_enable_390), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[2])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i2.GSR = "DISABLED";
    FD1P3IX baud_divider_i7 (.D(\data_to_write[7] ), .SP(clk_c_enable_390), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[7])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i7.GSR = "DISABLED";
    FD1P3IX baud_divider_i8 (.D(\data_to_write[8] ), .SP(clk_c_enable_395), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[8])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i8.GSR = "DISABLED";
    FD1P3IX baud_divider_i9 (.D(\data_to_write[9] ), .SP(clk_c_enable_395), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[9])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i9.GSR = "DISABLED";
    FD1P3IX baud_divider_i10 (.D(\data_to_write[10] ), .SP(clk_c_enable_395), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[10])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i10.GSR = "DISABLED";
    FD1P3IX baud_divider_i11 (.D(\data_to_write[11] ), .SP(clk_c_enable_395), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[11])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i11.GSR = "DISABLED";
    FD1P3IX baud_divider_i12 (.D(\data_to_write[12] ), .SP(clk_c_enable_395), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(baud_divider[12])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(37[12] 46[8])
    defparam baud_divider_i12.GSR = "DISABLED";
    LUT4 ui_in_7__I_0_3_lut_rep_795 (.A(\ui_in_sync[7] ), .B(\ui_in_sync[3] ), 
         .C(rxd_select), .Z(n32000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(82[21:53])
    defparam ui_in_7__I_0_3_lut_rep_795.init = 16'hcaca;
    LUT4 i15791_2_lut_4_lut (.A(\ui_in_sync[7] ), .B(\ui_in_sync[3] ), .C(rxd_select), 
         .D(mid_bit), .Z(next_fsm_state_3__N_3011[1])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(82[21:53])
    defparam i15791_2_lut_4_lut.init = 16'hcaff;
    FD1P3AX uart_rx_buf_data_i0_i1 (.D(uart_rx_data[1]), .SP(clk_c_enable_542), 
            .CK(clk_c), .Q(uart_rx_buf_data[1])) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i1.GSR = "DISABLED";
    FD1P3AX uart_rx_buffered_59 (.D(n27347), .SP(clk_c_enable_535), .CK(clk_c), 
            .Q(\next_fsm_state_3__N_3015[3] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buffered_59.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i2 (.D(uart_rx_data[2]), .SP(clk_c_enable_542), 
            .CK(clk_c), .Q(\uart_rx_buf_data[2] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i2.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i3 (.D(uart_rx_data[3]), .SP(clk_c_enable_542), 
            .CK(clk_c), .Q(\uart_rx_buf_data[3] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i3.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i4 (.D(uart_rx_data[4]), .SP(clk_c_enable_542), 
            .CK(clk_c), .Q(\uart_rx_buf_data[4] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i4.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i5 (.D(uart_rx_data[5]), .SP(clk_c_enable_542), 
            .CK(clk_c), .Q(\uart_rx_buf_data[5] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i5.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i6 (.D(uart_rx_data[6]), .SP(clk_c_enable_542), 
            .CK(clk_c), .Q(\uart_rx_buf_data[6] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i6.GSR = "DISABLED";
    FD1P3AX uart_rx_buf_data_i0_i7 (.D(uart_rx_data[7]), .SP(clk_c_enable_542), 
            .CK(clk_c), .Q(\uart_rx_buf_data[7] )) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=45, LSE_RCOL=3, LSE_LLINE=190, LSE_RLINE=202 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam uart_rx_buf_data_i0_i7.GSR = "DISABLED";
    LUT4 i27718_3_lut_rep_606_4_lut (.A(n31922), .B(clk_c_enable_185), .C(rst_reg_n), 
         .D(n31932), .Z(n31811)) /* synthesis lut_function=(!(A (C (D))+!A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(69[21:63])
    defparam i27718_3_lut_rep_606_4_lut.init = 16'h0fbf;
    LUT4 i1_2_lut_4_lut_2_lut_2_lut (.A(rst_reg_n), .B(n31932), .Z(n9493)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(69[21:63])
    defparam i1_2_lut_4_lut_2_lut_2_lut.init = 16'h7777;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n31922), .B(clk_c_enable_185), .C(n26116), 
         .D(n31932), .Z(n26118)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(69[21:63])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_3_lut_rep_700 (.A(\addr[9] ), .B(n26216), .C(\addr[10] ), 
         .Z(n31905)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_3_lut_rep_700.init = 16'h0404;
    LUT4 i1_2_lut_rep_681_4_lut (.A(\addr[9] ), .B(n26216), .C(\addr[10] ), 
         .D(n32033), .Z(clk_c_enable_185)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_681_4_lut.init = 16'h0004;
    LUT4 i27360_3_lut_4_lut (.A(\next_fsm_state_3__N_3015[3] ), .B(n31929), 
         .C(\imm[6] ), .D(\csr_read_3__N_1447[2] ), .Z(n29162)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(100[12] 113[8])
    defparam i27360_3_lut_4_lut.init = 16'h8f80;
    LUT4 uart_rx_buf_data_1__bdd_2_lut (.A(baud_divider[1]), .B(\addr[2] ), 
         .Z(n31474)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam uart_rx_buf_data_1__bdd_2_lut.init = 16'h2222;
    LUT4 uart_rx_buf_data_1__bdd_3_lut (.A(uart_rx_buf_data[1]), .B(\next_fsm_state_3__N_3015[3] ), 
         .C(\addr[2] ), .Z(n31475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam uart_rx_buf_data_1__bdd_3_lut.init = 16'hcaca;
    PFUMX i26553 (.BLUT(n29168), .ALUT(n29169), .C0(\addr[3] ), .Z(n29170));
    tqvp_uart_tx i_uart_tx (.cycle_counter({cycle_counter}), .clk_c(clk_c), 
            .clk_c_enable_152(clk_c_enable_152), .n6158(n6158), .n72({n72}), 
            .clk_c_enable_525(clk_c_enable_525), .clk_c_enable_445(clk_c_enable_445), 
            .fsm_state({fsm_state}), .n31811(n31811), .\uo_out_from_user_peri[2][6] (\uo_out_from_user_peri[2][6] ), 
            .n31932(n31932), .n31855(n31855), .\data_to_write[0] (\data_to_write[0] ), 
            .next_bit(next_bit), .\data_to_write[4] (\data_to_write[4] ), 
            .\data_to_write[6] (\data_to_write[6] ), .\data_to_write[5] (\data_to_write[5] ), 
            .\data_to_write[3] (\data_to_write[3] ), .\data_to_write[2] (\data_to_write[2] ), 
            .\data_to_write[1] (\data_to_write[1] ), .n9493(n9493), .n26118(n26118), 
            .n18596(n18596), .n31963(n31963), .\addr[2] (\addr[2] ), .\uart_rx_buf_data[0] (uart_rx_buf_data[0]), 
            .n29168(n29168)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(65[18] 73[6])
    tqvp_uart_rx i_uart_rx (.uart_rx_data({uart_rx_data}), .clk_c(clk_c), 
            .fsm_state({fsm_state_adj_50}), .next_bit(next_bit_adj_34), 
            .cycle_counter({cycle_counter_adj_51}), .clk_c_enable_445(clk_c_enable_445), 
            .\uo_out_from_user_peri[2][7] (\uo_out_from_user_peri[2][7] ), 
            .\next_fsm_state_3__N_3011[1] (next_fsm_state_3__N_3011[1]), .\next_fsm_state_3__N_3015[3] (\next_fsm_state_3__N_3015[3] ), 
            .n32000(n32000), .mid_bit(mid_bit), .rst_reg_n(rst_reg_n), 
            .n28760(n28760), .n31922(n31922), .clk_c_enable_535(clk_c_enable_535), 
            .\baud_divider[4] (baud_divider[4]), .\baud_divider[3] (baud_divider[3]), 
            .\baud_divider[2] (baud_divider[2]), .\baud_divider[1] (baud_divider[1]), 
            .GND_net(GND_net), .VCC_net(VCC_net), .\baud_divider[8] (baud_divider[8]), 
            .\baud_divider[7] (baud_divider[7]), .\baud_divider[6] (baud_divider[6]), 
            .\baud_divider[5] (baud_divider[5]), .\baud_divider[12] (baud_divider[12]), 
            .\baud_divider[11] (baud_divider[11]), .\baud_divider[10] (baud_divider[10]), 
            .\baud_divider[9] (baud_divider[9]), .n31902(n31902), .n31925(n31925), 
            .n32003(n32003), .clk_c_enable_223(clk_c_enable_223), .n31923(n31923), 
            .\addr[4] (\addr[4] ), .clk_c_enable_275(clk_c_enable_275), 
            .next_bit_adj_26(next_bit_adj_48), .n31828(n31828), .uart_txd_N_2974(uart_txd_N_2974), 
            .clk_c_enable_534(clk_c_enable_534), .debug_stop_txn(debug_stop_txn), 
            .instr_active_N_2106(instr_active_N_2106), .clk_c_enable_344(clk_c_enable_344), 
            .n3(n3), .\data_to_write[0] (\data_to_write[0] ), .rxd_select(rxd_select), 
            .n29200(n29200), .n32013(n32013), .\fsm_state[0]_adj_27 (\fsm_state[0]_adj_49 ), 
            .clk_c_enable_376(clk_c_enable_376), .n28686(n28686), .n31880(n31880), 
            .clk_c_enable_355(clk_c_enable_355), .n8005(n8005), .n1084(n1084), 
            .stop_txn_reg(stop_txn_reg), .stop_txn_now_N_2363(stop_txn_now_N_2363), 
            .clk_c_enable_239(clk_c_enable_239), .n31971(n31971), .n33479(n33479), 
            .\qspi_data_in[1] (\qspi_data_in[1] ), .n31593(n31593), .n26266(n26266), 
            .n31927(n31927), .clk_c_enable_378(clk_c_enable_378), .n27620(n27620), 
            .n31906(n31906), .n27081(n27081), .clk_c_enable_377(clk_c_enable_377), 
            .n6210(n6210), .n18596(n18596), .n31819(n31819), .n28800(n28800), 
            .clk_c_enable_525(clk_c_enable_525), .n32027(n32027), .n32034(n32034), 
            .clk_c_enable_531(clk_c_enable_531), .next_bit_adj_28(next_bit), 
            .n6158(n6158), .n31963(n31963), .\fsm_state[0]_adj_29 (fsm_state[0]), 
            .clk_c_enable_152(clk_c_enable_152), .n31950(n31950), .n18241(n18241), 
            .clk_c_enable_268(clk_c_enable_268), .clk_c_enable_469(clk_c_enable_469), 
            .clk_c_enable_386(clk_c_enable_386), .\data_to_write[1] (\data_to_write[1] ), 
            .n8695(n8695), .n31977(n31977), .n8135(n8135), .n10499(n10499), 
            .n10500(n10500), .clk_c_enable_186(clk_c_enable_186), .n32021(n32021), 
            .n31997(n31997), .\addr[27] (\addr[27] ), .n31930(n31930), 
            .n32022(n32022), .n31958(n31958), .n26036(n26036), .instr_complete_N_1647(instr_complete_N_1647), 
            .n28276(n28276), .n31883(n31883), .clk_c_enable_115(clk_c_enable_115), 
            .n32019(n32019), .clk_c_enable_334(clk_c_enable_334), .n31717(n31717), 
            .n80(n80), .clk_c_enable_10(clk_c_enable_10)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/peri_uart.v(85[18] 94[6])
    
endmodule
//
// Verilog Description of module tqvp_uart_tx
//

module tqvp_uart_tx (cycle_counter, clk_c, clk_c_enable_152, n6158, 
            n72, clk_c_enable_525, clk_c_enable_445, fsm_state, n31811, 
            \uo_out_from_user_peri[2][6] , n31932, n31855, \data_to_write[0] , 
            next_bit, \data_to_write[4] , \data_to_write[6] , \data_to_write[5] , 
            \data_to_write[3] , \data_to_write[2] , \data_to_write[1] , 
            n9493, n26118, n18596, n31963, \addr[2] , \uart_rx_buf_data[0] , 
            n29168) /* synthesis syn_module_defined=1 */ ;
    output [12:0]cycle_counter;
    input clk_c;
    input clk_c_enable_152;
    input n6158;
    input [12:0]n72;
    input clk_c_enable_525;
    input clk_c_enable_445;
    output [3:0]fsm_state;
    input n31811;
    output \uo_out_from_user_peri[2][6] ;
    input n31932;
    input n31855;
    input \data_to_write[0] ;
    input next_bit;
    input \data_to_write[4] ;
    input \data_to_write[6] ;
    input \data_to_write[5] ;
    input \data_to_write[3] ;
    input \data_to_write[2] ;
    input \data_to_write[1] ;
    input n9493;
    input n26118;
    output n18596;
    input n31963;
    input \addr[2] ;
    input \uart_rx_buf_data[0] ;
    output n29168;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [7:0]data_to_send;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(39[24:36])
    wire [7:0]data_to_send_7__N_2944;
    
    wire clk_c_enable_244, n32060, uart_txd_N_2972;
    wire [3:0]n162;
    
    wire n31552, n31551;
    
    FD1P3IX cycle_counter__i0 (.D(n72[0]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i0.GSR = "DISABLED";
    FD1P3IX data_to_send__i0 (.D(data_to_send_7__N_2944[0]), .SP(clk_c_enable_525), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i0.GSR = "DISABLED";
    FD1P3IX cycle_counter__i12 (.D(n72[12]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[12])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i12.GSR = "DISABLED";
    FD1P3IX cycle_counter__i11 (.D(n72[11]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[11])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i11.GSR = "DISABLED";
    FD1P3IX cycle_counter__i10 (.D(n72[10]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[10])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i10.GSR = "DISABLED";
    FD1P3IX cycle_counter__i9 (.D(n72[9]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[9])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i9.GSR = "DISABLED";
    FD1P3IX cycle_counter__i8 (.D(n72[8]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[8])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i8.GSR = "DISABLED";
    FD1P3IX cycle_counter__i7 (.D(n72[7]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[7])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i7.GSR = "DISABLED";
    FD1P3IX cycle_counter__i6 (.D(n72[6]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[6])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i6.GSR = "DISABLED";
    FD1P3IX cycle_counter__i5 (.D(n72[5]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[5])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i5.GSR = "DISABLED";
    FD1P3IX cycle_counter__i4 (.D(n72[4]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[4])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i4.GSR = "DISABLED";
    FD1P3IX cycle_counter__i3 (.D(n72[3]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i3.GSR = "DISABLED";
    FD1P3IX cycle_counter__i2 (.D(n72[2]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i2.GSR = "DISABLED";
    FD1P3IX cycle_counter__i1 (.D(n72[1]), .SP(clk_c_enable_152), .CD(n6158), 
            .CK(clk_c), .Q(cycle_counter[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i1.GSR = "DISABLED";
    FD1P3IX fsm_state__i0 (.D(n32060), .SP(clk_c_enable_244), .CD(n31811), 
            .CK(clk_c), .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i0.GSR = "DISABLED";
    FD1S3JX txd_reg_46 (.D(uart_txd_N_2972), .CK(clk_c), .PD(clk_c_enable_445), 
            .Q(\uo_out_from_user_peri[2][6] )) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(123[8] 133[4])
    defparam txd_reg_46.GSR = "DISABLED";
    LUT4 mux_13_i1_3_lut_4_lut (.A(n31932), .B(n31855), .C(\data_to_write[0] ), 
         .D(data_to_send[1]), .Z(data_to_send_7__N_2944[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut (.A(n31932), .B(n31855), .C(next_bit), .D(n31811), 
         .Z(clk_c_enable_244)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam i1_3_lut_4_lut.init = 16'hfff4;
    LUT4 mux_13_i5_3_lut_4_lut (.A(n31932), .B(n31855), .C(\data_to_write[4] ), 
         .D(data_to_send[5]), .Z(data_to_send_7__N_2944[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i7_3_lut_4_lut (.A(n31932), .B(n31855), .C(\data_to_write[6] ), 
         .D(data_to_send[7]), .Z(data_to_send_7__N_2944[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i6_3_lut_4_lut (.A(n31932), .B(n31855), .C(\data_to_write[5] ), 
         .D(data_to_send[6]), .Z(data_to_send_7__N_2944[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i4_3_lut_4_lut (.A(n31932), .B(n31855), .C(\data_to_write[3] ), 
         .D(data_to_send[4]), .Z(data_to_send_7__N_2944[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i3_3_lut_4_lut (.A(n31932), .B(n31855), .C(\data_to_write[2] ), 
         .D(data_to_send[3]), .Z(data_to_send_7__N_2944[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i2_3_lut_4_lut (.A(n31932), .B(n31855), .C(\data_to_write[1] ), 
         .D(data_to_send[2]), .Z(data_to_send_7__N_2944[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 fsm_state_0__bdd_4_lut (.A(fsm_state[0]), .B(fsm_state[2]), .C(fsm_state[1]), 
         .D(fsm_state[3]), .Z(n32060)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;
    defparam fsm_state_0__bdd_4_lut.init = 16'h4555;
    LUT4 i1_3_lut_3_lut_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(fsm_state[0]), .Z(n162[1])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(D)))) */ ;
    defparam i1_3_lut_3_lut_4_lut.init = 16'h33c4;
    FD1P3IX data_to_send__i6 (.D(data_to_send_7__N_2944[6]), .SP(clk_c_enable_525), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[6])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i6.GSR = "DISABLED";
    FD1P3IX data_to_send__i5 (.D(data_to_send_7__N_2944[5]), .SP(clk_c_enable_525), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[5])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i5.GSR = "DISABLED";
    FD1P3IX data_to_send__i4 (.D(data_to_send_7__N_2944[4]), .SP(clk_c_enable_525), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[4])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i4.GSR = "DISABLED";
    FD1P3IX data_to_send__i3 (.D(data_to_send_7__N_2944[3]), .SP(clk_c_enable_525), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i3.GSR = "DISABLED";
    FD1P3IX data_to_send__i2 (.D(data_to_send_7__N_2944[2]), .SP(clk_c_enable_525), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i2.GSR = "DISABLED";
    FD1P3IX data_to_send__i1 (.D(data_to_send_7__N_2944[1]), .SP(clk_c_enable_525), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i1.GSR = "DISABLED";
    FD1P3IX fsm_state__i1 (.D(n162[1]), .SP(next_bit), .CD(n9493), .CK(clk_c), 
            .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i1.GSR = "DISABLED";
    FD1P3IX fsm_state__i2 (.D(n31552), .SP(next_bit), .CD(n9493), .CK(clk_c), 
            .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1P3IX fsm_state__i3 (.D(n31551), .SP(next_bit), .CD(n9493), .CK(clk_c), 
            .Q(fsm_state[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i3.GSR = "DISABLED";
    FD1P3AX data_to_send__i7 (.D(n26118), .SP(clk_c_enable_525), .CK(clk_c), 
            .Q(data_to_send[7])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=65, LSE_RLINE=73 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i7.GSR = "DISABLED";
    LUT4 i16023_3_lut (.A(fsm_state[1]), .B(fsm_state[3]), .C(fsm_state[2]), 
         .Z(n18596)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i16023_3_lut.init = 16'hc8c8;
    LUT4 i20106_4_lut (.A(fsm_state[0]), .B(n18596), .C(n31963), .D(data_to_send[0]), 
         .Z(uart_txd_N_2972)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(21[25:33])
    defparam i20106_4_lut.init = 16'hf5c5;
    LUT4 i26551_3_lut_4_lut (.A(fsm_state[0]), .B(n31963), .C(\addr[2] ), 
         .D(\uart_rx_buf_data[0] ), .Z(n29168)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i26551_3_lut_4_lut.init = 16'hefe0;
    LUT4 fsm_state_1__bdd_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[0]), 
         .Z(n31552)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;
    defparam fsm_state_1__bdd_3_lut.init = 16'h6c6c;
    LUT4 fsm_state_1__bdd_4_lut (.A(fsm_state[1]), .B(fsm_state[3]), .C(fsm_state[2]), 
         .D(fsm_state[0]), .Z(n31551)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)))+!A !(B))) */ ;
    defparam fsm_state_1__bdd_4_lut.init = 16'h6cc4;
    
endmodule
//
// Verilog Description of module tqvp_uart_rx
//

module tqvp_uart_rx (uart_rx_data, clk_c, fsm_state, next_bit, cycle_counter, 
            clk_c_enable_445, \uo_out_from_user_peri[2][7] , \next_fsm_state_3__N_3011[1] , 
            \next_fsm_state_3__N_3015[3] , n32000, mid_bit, rst_reg_n, 
            n28760, n31922, clk_c_enable_535, \baud_divider[4] , \baud_divider[3] , 
            \baud_divider[2] , \baud_divider[1] , GND_net, VCC_net, 
            \baud_divider[8] , \baud_divider[7] , \baud_divider[6] , \baud_divider[5] , 
            \baud_divider[12] , \baud_divider[11] , \baud_divider[10] , 
            \baud_divider[9] , n31902, n31925, n32003, clk_c_enable_223, 
            n31923, \addr[4] , clk_c_enable_275, next_bit_adj_26, n31828, 
            uart_txd_N_2974, clk_c_enable_534, debug_stop_txn, instr_active_N_2106, 
            clk_c_enable_344, n3, \data_to_write[0] , rxd_select, n29200, 
            n32013, \fsm_state[0]_adj_27 , clk_c_enable_376, n28686, 
            n31880, clk_c_enable_355, n8005, n1084, stop_txn_reg, 
            stop_txn_now_N_2363, clk_c_enable_239, n31971, n33479, \qspi_data_in[1] , 
            n31593, n26266, n31927, clk_c_enable_378, n27620, n31906, 
            n27081, clk_c_enable_377, n6210, n18596, n31819, n28800, 
            clk_c_enable_525, n32027, n32034, clk_c_enable_531, next_bit_adj_28, 
            n6158, n31963, \fsm_state[0]_adj_29 , clk_c_enable_152, 
            n31950, n18241, clk_c_enable_268, clk_c_enable_469, clk_c_enable_386, 
            \data_to_write[1] , n8695, n31977, n8135, n10499, n10500, 
            clk_c_enable_186, n32021, n31997, \addr[27] , n31930, 
            n32022, n31958, n26036, instr_complete_N_1647, n28276, 
            n31883, clk_c_enable_115, n32019, clk_c_enable_334, n31717, 
            n80, clk_c_enable_10) /* synthesis syn_module_defined=1 */ ;
    output [7:0]uart_rx_data;
    input clk_c;
    output [3:0]fsm_state;
    input next_bit;
    output [12:0]cycle_counter;
    output clk_c_enable_445;
    output \uo_out_from_user_peri[2][7] ;
    input \next_fsm_state_3__N_3011[1] ;
    input \next_fsm_state_3__N_3015[3] ;
    input n32000;
    output mid_bit;
    input rst_reg_n;
    input n28760;
    input n31922;
    output clk_c_enable_535;
    input \baud_divider[4] ;
    input \baud_divider[3] ;
    input \baud_divider[2] ;
    input \baud_divider[1] ;
    input GND_net;
    input VCC_net;
    input \baud_divider[8] ;
    input \baud_divider[7] ;
    input \baud_divider[6] ;
    input \baud_divider[5] ;
    input \baud_divider[12] ;
    input \baud_divider[11] ;
    input \baud_divider[10] ;
    input \baud_divider[9] ;
    input n31902;
    input n31925;
    input n32003;
    output clk_c_enable_223;
    input n31923;
    input \addr[4] ;
    output clk_c_enable_275;
    input next_bit_adj_26;
    input n31828;
    input uart_txd_N_2974;
    output clk_c_enable_534;
    input debug_stop_txn;
    output instr_active_N_2106;
    output clk_c_enable_344;
    input n3;
    input \data_to_write[0] ;
    input rxd_select;
    output n29200;
    input n32013;
    input \fsm_state[0]_adj_27 ;
    output clk_c_enable_376;
    input n28686;
    input n31880;
    output clk_c_enable_355;
    output n8005;
    input n1084;
    input stop_txn_reg;
    input stop_txn_now_N_2363;
    output clk_c_enable_239;
    input n31971;
    input n33479;
    input \qspi_data_in[1] ;
    output n31593;
    input n26266;
    input n31927;
    output clk_c_enable_378;
    input n27620;
    input n31906;
    output n27081;
    output clk_c_enable_377;
    output n6210;
    input n18596;
    input n31819;
    input n28800;
    output clk_c_enable_525;
    input n32027;
    input n32034;
    output clk_c_enable_531;
    input next_bit_adj_28;
    output n6158;
    input n31963;
    input \fsm_state[0]_adj_29 ;
    output clk_c_enable_152;
    output n31950;
    input n18241;
    input clk_c_enable_268;
    output clk_c_enable_469;
    output clk_c_enable_386;
    input \data_to_write[1] ;
    output n8695;
    input n31977;
    output n8135;
    input n10499;
    output n10500;
    output clk_c_enable_186;
    input n32021;
    input n31997;
    input \addr[27] ;
    output n31930;
    input n32022;
    input n31958;
    output n26036;
    input instr_complete_N_1647;
    input n28276;
    input n31883;
    output clk_c_enable_115;
    input n32019;
    output clk_c_enable_334;
    output n31717;
    input n80;
    output clk_c_enable_10;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire uart_rx_data_7__N_3059, n32091;
    wire [2:0]n5272;
    
    wire n32090, n1117;
    wire [12:0]n57;
    wire [3:0]next_fsm_state;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(71[11:25])
    
    wire uart_rts_N_3079, n32051, n31775, bit_sample, clk_c_enable_361;
    wire [2:0]n5252;
    
    wire n23550, n23551, n23679, n23678, n9, n23677, n23676, n23675, 
        n9470;
    wire [31:0]next_fsm_state_3__N_3027;
    
    wire n23548, n23549, n23674, n29255;
    
    FD1P3AX recieved_data_i0_i0 (.D(uart_rx_data[1]), .SP(uart_rx_data_7__N_3059), 
            .CK(clk_c), .Q(uart_rx_data[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i0.GSR = "DISABLED";
    LUT4 mux_3032_i4_4_lut_then_4_lut (.A(fsm_state[3]), .B(fsm_state[1]), 
         .C(next_bit), .D(fsm_state[0]), .Z(n32091)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3032_i4_4_lut_then_4_lut.init = 16'h6aaa;
    LUT4 mux_3032_i4_4_lut_else_4_lut (.A(fsm_state[3]), .B(n5272[1]), .C(fsm_state[1]), 
         .D(fsm_state[0]), .Z(n32090)) /* synthesis lut_function=(A (B+!(C))+!A !((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3032_i4_4_lut_else_4_lut.init = 16'h8a8e;
    FD1S3IX cycle_counter_3565__i0 (.D(n57[0]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i0.GSR = "DISABLED";
    FD1S3IX fsm_state__i0 (.D(next_fsm_state[0]), .CK(clk_c), .CD(clk_c_enable_445), 
            .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(136[8] 142[4])
    defparam fsm_state__i0.GSR = "DISABLED";
    FD1S3JX uart_rts_50 (.D(uart_rts_N_3079), .CK(clk_c), .PD(clk_c_enable_445), 
            .Q(\uo_out_from_user_peri[2][7] )) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(145[8] 152[4])
    defparam uart_rts_50.GSR = "DISABLED";
    LUT4 mux_3032_i2_4_lut (.A(fsm_state[1]), .B(n5272[1]), .C(n32051), 
         .D(n31775), .Z(next_fsm_state[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3032_i2_4_lut.init = 16'hc5ca;
    LUT4 mux_3173_i2_4_lut (.A(\next_fsm_state_3__N_3011[1] ), .B(\next_fsm_state_3__N_3015[3] ), 
         .C(fsm_state[0]), .D(fsm_state[1]), .Z(n5272[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3173_i2_4_lut.init = 16'hcac0;
    FD1P3IX bit_sample_47 (.D(n32000), .SP(clk_c_enable_361), .CD(clk_c_enable_445), 
            .CK(clk_c), .Q(bit_sample)) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(112[8] 118[4])
    defparam bit_sample_47.GSR = "DISABLED";
    LUT4 mux_3173_i1_4_lut (.A(\next_fsm_state_3__N_3015[3] ), .B(fsm_state[0]), 
         .C(n32051), .D(next_bit), .Z(n5272[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A !(B (C+(D))+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3173_i1_4_lut.init = 16'ha3ac;
    LUT4 mux_3169_i1_3_lut (.A(n32000), .B(mid_bit), .C(fsm_state[1]), 
         .Z(n5252[0])) /* synthesis lut_function=(A (B (C))+!A !(C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(73[3] 95[10])
    defparam mux_3169_i1_3_lut.init = 16'h8585;
    FD1P3AX recieved_data_i0_i1 (.D(uart_rx_data[2]), .SP(uart_rx_data_7__N_3059), 
            .CK(clk_c), .Q(uart_rx_data[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i1.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i2 (.D(uart_rx_data[3]), .SP(uart_rx_data_7__N_3059), 
            .CK(clk_c), .Q(uart_rx_data[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i2.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i3 (.D(uart_rx_data[4]), .SP(uart_rx_data_7__N_3059), 
            .CK(clk_c), .Q(uart_rx_data[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i3.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i4 (.D(uart_rx_data[5]), .SP(uart_rx_data_7__N_3059), 
            .CK(clk_c), .Q(uart_rx_data[4])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i4.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i5 (.D(uart_rx_data[6]), .SP(uart_rx_data_7__N_3059), 
            .CK(clk_c), .Q(uart_rx_data[5])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i5.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i6 (.D(uart_rx_data[7]), .SP(uart_rx_data_7__N_3059), 
            .CK(clk_c), .Q(uart_rx_data[6])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i6.GSR = "DISABLED";
    FD1P3AX recieved_data_i0_i7 (.D(bit_sample), .SP(uart_rx_data_7__N_3059), 
            .CK(clk_c), .Q(uart_rx_data[7])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(104[8] 108[4])
    defparam recieved_data_i0_i7.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(rst_reg_n), .B(n28760), .C(\next_fsm_state_3__N_3015[3] ), 
         .D(n31922), .Z(clk_c_enable_535)) /* synthesis lut_function=(!(A (B (C (D))+!B (C)))) */ ;
    defparam i1_4_lut.init = 16'h5fdf;
    CCU2C cycle_counter_12__I_0_13_21152 (.A0(\baud_divider[4] ), .B0(cycle_counter[3]), 
          .C0(\baud_divider[3] ), .D0(cycle_counter[2]), .A1(\baud_divider[2] ), 
          .B1(cycle_counter[1]), .C1(\baud_divider[1] ), .D1(cycle_counter[0]), 
          .CIN(n23550), .COUT(n23551));
    defparam cycle_counter_12__I_0_13_21152.INIT0 = 16'h9009;
    defparam cycle_counter_12__I_0_13_21152.INIT1 = 16'h9009;
    defparam cycle_counter_12__I_0_13_21152.INJECT1_0 = "YES";
    defparam cycle_counter_12__I_0_13_21152.INJECT1_1 = "YES";
    CCU2C cycle_counter_3565_add_4_13 (.A0(cycle_counter[11]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[12]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23679), .S0(n57[11]), .S1(n57[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565_add_4_13.INIT0 = 16'haaa0;
    defparam cycle_counter_3565_add_4_13.INIT1 = 16'haaa0;
    defparam cycle_counter_3565_add_4_13.INJECT1_0 = "NO";
    defparam cycle_counter_3565_add_4_13.INJECT1_1 = "NO";
    CCU2C cycle_counter_3565_add_4_11 (.A0(cycle_counter[9]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[10]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23678), .COUT(n23679), .S0(n57[9]), 
          .S1(n57[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565_add_4_11.INIT0 = 16'haaa0;
    defparam cycle_counter_3565_add_4_11.INIT1 = 16'haaa0;
    defparam cycle_counter_3565_add_4_11.INJECT1_0 = "NO";
    defparam cycle_counter_3565_add_4_11.INJECT1_1 = "NO";
    FD1S3IX cycle_counter_3565__i1 (.D(n57[1]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i1.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i2 (.D(n57[2]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i2.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i3 (.D(n57[3]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i3.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i4 (.D(n57[4]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i4.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i5 (.D(n57[5]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i5.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i6 (.D(n57[6]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i6.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i7 (.D(n57[7]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i7.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i8 (.D(n57[8]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i8.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i9 (.D(n57[9]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i9.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i10 (.D(n57[10]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i10.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i11 (.D(n57[11]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i11.GSR = "DISABLED";
    FD1S3IX cycle_counter_3565__i12 (.D(n57[12]), .CK(clk_c), .CD(n1117), 
            .Q(cycle_counter[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565__i12.GSR = "DISABLED";
    LUT4 uart_rts_I_258_2_lut_3_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[3]), 
         .C(\next_fsm_state_3__N_3015[3] ), .D(fsm_state[2]), .Z(uart_rts_N_3079)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam uart_rts_I_258_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i22_4_lut_3_lut (.A(fsm_state[1]), .B(fsm_state[3]), .C(fsm_state[0]), 
         .Z(n9)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;
    defparam i22_4_lut_3_lut.init = 16'h8181;
    CCU2C cycle_counter_3565_add_4_9 (.A0(cycle_counter[7]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[8]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23677), .COUT(n23678), .S0(n57[7]), 
          .S1(n57[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565_add_4_9.INIT0 = 16'haaa0;
    defparam cycle_counter_3565_add_4_9.INIT1 = 16'haaa0;
    defparam cycle_counter_3565_add_4_9.INJECT1_0 = "NO";
    defparam cycle_counter_3565_add_4_9.INJECT1_1 = "NO";
    FD1S3IX fsm_state__i1 (.D(next_fsm_state[1]), .CK(clk_c), .CD(clk_c_enable_445), 
            .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(136[8] 142[4])
    defparam fsm_state__i1.GSR = "DISABLED";
    CCU2C cycle_counter_3565_add_4_7 (.A0(cycle_counter[5]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[6]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23676), .COUT(n23677), .S0(n57[5]), 
          .S1(n57[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565_add_4_7.INIT0 = 16'haaa0;
    defparam cycle_counter_3565_add_4_7.INIT1 = 16'haaa0;
    defparam cycle_counter_3565_add_4_7.INJECT1_0 = "NO";
    defparam cycle_counter_3565_add_4_7.INJECT1_1 = "NO";
    CCU2C cycle_counter_3565_add_4_5 (.A0(cycle_counter[3]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[4]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23675), .COUT(n23676), .S0(n57[3]), 
          .S1(n57[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565_add_4_5.INIT0 = 16'haaa0;
    defparam cycle_counter_3565_add_4_5.INIT1 = 16'haaa0;
    defparam cycle_counter_3565_add_4_5.INJECT1_0 = "NO";
    defparam cycle_counter_3565_add_4_5.INJECT1_1 = "NO";
    FD1S3IX fsm_state__i2 (.D(next_fsm_state_3__N_3027[2]), .CK(clk_c), 
            .CD(n9470), .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(136[8] 142[4])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1S3IX fsm_state__i3 (.D(next_fsm_state[3]), .CK(clk_c), .CD(clk_c_enable_445), 
            .Q(fsm_state[3])) /* synthesis LSE_LINE_FILE_ID=22, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=85, LSE_RLINE=94 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(136[8] 142[4])
    defparam fsm_state__i3.GSR = "DISABLED";
    CCU2C cycle_counter_12__I_0_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cycle_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n23548));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(67[21:55])
    defparam cycle_counter_12__I_0_0.INIT0 = 16'h000F;
    defparam cycle_counter_12__I_0_0.INIT1 = 16'h5555;
    defparam cycle_counter_12__I_0_0.INJECT1_0 = "NO";
    defparam cycle_counter_12__I_0_0.INJECT1_1 = "YES";
    CCU2C cycle_counter_12__I_0_11 (.A0(\baud_divider[8] ), .B0(cycle_counter[7]), 
          .C0(\baud_divider[7] ), .D0(cycle_counter[6]), .A1(\baud_divider[6] ), 
          .B1(cycle_counter[5]), .C1(\baud_divider[5] ), .D1(cycle_counter[4]), 
          .CIN(n23549), .COUT(n23550));
    defparam cycle_counter_12__I_0_11.INIT0 = 16'h9009;
    defparam cycle_counter_12__I_0_11.INIT1 = 16'h9009;
    defparam cycle_counter_12__I_0_11.INJECT1_0 = "YES";
    defparam cycle_counter_12__I_0_11.INJECT1_1 = "YES";
    CCU2C cycle_counter_3565_add_4_3 (.A0(cycle_counter[1]), .B0(GND_net), 
          .C0(GND_net), .D0(VCC_net), .A1(cycle_counter[2]), .B1(GND_net), 
          .C1(GND_net), .D1(VCC_net), .CIN(n23674), .COUT(n23675), .S0(n57[1]), 
          .S1(n57[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565_add_4_3.INIT0 = 16'haaa0;
    defparam cycle_counter_3565_add_4_3.INIT1 = 16'haaa0;
    defparam cycle_counter_3565_add_4_3.INJECT1_0 = "NO";
    defparam cycle_counter_3565_add_4_3.INJECT1_1 = "NO";
    CCU2C cycle_counter_3565_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycle_counter[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n23674), .S1(n57[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(129[26:46])
    defparam cycle_counter_3565_add_4_1.INIT0 = 16'h0000;
    defparam cycle_counter_3565_add_4_1.INIT1 = 16'h555f;
    defparam cycle_counter_3565_add_4_1.INJECT1_0 = "NO";
    defparam cycle_counter_3565_add_4_1.INJECT1_1 = "NO";
    CCU2C cycle_counter_12__I_0_9 (.A0(\baud_divider[12] ), .B0(cycle_counter[11]), 
          .C0(\baud_divider[11] ), .D0(cycle_counter[10]), .A1(\baud_divider[10] ), 
          .B1(cycle_counter[9]), .C1(\baud_divider[9] ), .D1(cycle_counter[8]), 
          .CIN(n23548), .COUT(n23549));
    defparam cycle_counter_12__I_0_9.INIT0 = 16'h9009;
    defparam cycle_counter_12__I_0_9.INIT1 = 16'h9009;
    defparam cycle_counter_12__I_0_9.INJECT1_0 = "YES";
    defparam cycle_counter_12__I_0_9.INJECT1_1 = "YES";
    LUT4 i4678_2_lut_rep_570 (.A(fsm_state[0]), .B(next_bit), .Z(n31775)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(93[33:48])
    defparam i4678_2_lut_rep_570.init = 16'h8888;
    LUT4 rst_reg_n_I_0_1_lut_rep_832 (.A(rst_reg_n), .Z(clk_c_enable_445)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam rst_reg_n_I_0_1_lut_rep_832.init = 16'h5555;
    LUT4 i1_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(n31902), .C(n31925), 
         .D(n32003), .Z(clk_c_enable_223)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h5d55;
    LUT4 i1_3_lut_4_lut_4_lut_adj_570 (.A(rst_reg_n), .B(n31902), .C(n31923), 
         .D(\addr[4] ), .Z(clk_c_enable_275)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_570.init = 16'h555d;
    LUT4 i1_4_lut_4_lut (.A(rst_reg_n), .B(next_bit_adj_26), .C(n31828), 
         .D(uart_txd_N_2974), .Z(clk_c_enable_534)) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut.init = 16'hfdf5;
    LUT4 rstn_N_2029_I_0_2_lut_2_lut (.A(rst_reg_n), .B(debug_stop_txn), 
         .Z(instr_active_N_2106)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam rstn_N_2029_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_571 (.A(rst_reg_n), .B(n31902), .C(n31923), 
         .D(\addr[4] ), .Z(clk_c_enable_344)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_571.init = 16'h5d55;
    LUT4 i26583_4_lut_4_lut (.A(rst_reg_n), .B(n3), .C(\data_to_write[0] ), 
         .D(rxd_select), .Z(n29200)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i26583_4_lut_4_lut.init = 16'hf2d0;
    LUT4 i1_3_lut_4_lut_4_lut_adj_572 (.A(rst_reg_n), .B(next_bit_adj_26), 
         .C(n32013), .D(\fsm_state[0]_adj_27 ), .Z(clk_c_enable_376)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_572.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_573 (.A(rst_reg_n), .B(n28686), .C(n31880), 
         .D(n32003), .Z(clk_c_enable_355)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_573.init = 16'hd555;
    LUT4 i15383_2_lut_2_lut (.A(rst_reg_n), .B(\data_to_write[0] ), .Z(n8005)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i15383_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n1084), .C(stop_txn_reg), 
         .D(stop_txn_now_N_2363), .Z(clk_c_enable_239)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_2_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 n5570_bdd_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(n31971), .C(n33479), 
         .D(\qspi_data_in[1] ), .Z(n31593)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam n5570_bdd_2_lut_3_lut_4_lut_4_lut.init = 16'h3010;
    LUT4 i1_3_lut_4_lut_4_lut_adj_574 (.A(rst_reg_n), .B(n31902), .C(n26266), 
         .D(n31927), .Z(clk_c_enable_378)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_574.init = 16'h555d;
    LUT4 i1_4_lut_4_lut_adj_575 (.A(rst_reg_n), .B(n27620), .C(stop_txn_now_N_2363), 
         .D(n31906), .Z(n27081)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_575.init = 16'hfffd;
    LUT4 i6870_2_lut_2_lut (.A(rst_reg_n), .B(n32051), .Z(n9470)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i6870_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_576 (.A(rst_reg_n), .B(n31902), .C(n31927), 
         .D(n32003), .Z(clk_c_enable_377)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_576.init = 16'h5d55;
    LUT4 i1_4_lut_4_lut_adj_577 (.A(rst_reg_n), .B(n9), .C(next_bit), 
         .D(fsm_state[2]), .Z(n1117)) /* synthesis lut_function=((B (C+!(D))+!B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_577.init = 16'hf5fd;
    LUT4 i459_2_lut_2_lut (.A(rst_reg_n), .B(next_bit_adj_26), .Z(n6210)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i459_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut_adj_578 (.A(rst_reg_n), .B(n18596), .C(n31819), 
         .D(n28800), .Z(clk_c_enable_525)) /* synthesis lut_function=((B (C)+!B (C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_578.init = 16'hf7f5;
    LUT4 i1_2_lut_4_lut_4_lut_adj_579 (.A(rst_reg_n), .B(n32027), .C(n31880), 
         .D(n32034), .Z(clk_c_enable_531)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_2_lut_4_lut_4_lut_adj_579.init = 16'h55d5;
    LUT4 i1_2_lut_2_lut (.A(rst_reg_n), .B(next_bit_adj_28), .Z(n6158)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_580 (.A(rst_reg_n), .B(next_bit_adj_28), 
         .C(n31963), .D(\fsm_state[0]_adj_29 ), .Z(clk_c_enable_152)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_580.init = 16'hfffd;
    LUT4 i15501_2_lut_rep_745_2_lut (.A(rst_reg_n), .B(\qspi_data_in[1] ), 
         .Z(n31950)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i15501_2_lut_rep_745_2_lut.init = 16'hdddd;
    LUT4 i3606_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(n31922), .C(n18241), 
         .D(clk_c_enable_268), .Z(clk_c_enable_469)) /* synthesis lut_function=(!(A (B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i3606_3_lut_4_lut_4_lut.init = 16'h5755;
    LUT4 i1_3_lut_4_lut_4_lut_adj_581 (.A(rst_reg_n), .B(n31902), .C(n26266), 
         .D(n31925), .Z(clk_c_enable_386)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_581.init = 16'h555d;
    LUT4 i15604_2_lut_2_lut (.A(rst_reg_n), .B(\data_to_write[1] ), .Z(n8695)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i15604_2_lut_2_lut.init = 16'hdddd;
    LUT4 i4691_2_lut_3_lut_4_lut (.A(fsm_state[0]), .B(next_bit), .C(fsm_state[2]), 
         .D(fsm_state[1]), .Z(next_fsm_state_3__N_3027[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_rx.v(93[33:48])
    defparam i4691_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_4_lut_4_lut_adj_582 (.A(rst_reg_n), .B(stop_txn_reg), .C(stop_txn_now_N_2363), 
         .D(n31977), .Z(n8135)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_582.init = 16'hfdff;
    LUT4 i1_2_lut_2_lut_adj_583 (.A(rst_reg_n), .B(n10499), .Z(n10500)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_2_lut_2_lut_adj_583.init = 16'hdddd;
    LUT4 i3882_2_lut_2_lut (.A(rst_reg_n), .B(mid_bit), .Z(clk_c_enable_361)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i3882_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut_adj_584 (.A(rst_reg_n), .B(stop_txn_reg), .C(n31977), 
         .D(stop_txn_now_N_2363), .Z(clk_c_enable_186)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_584.init = 16'hfffd;
    LUT4 i1_3_lut_rep_725_4_lut_4_lut (.A(rst_reg_n), .B(n32021), .C(n31997), 
         .D(\addr[27] ), .Z(n31930)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_rep_725_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_4_lut_4_lut_adj_585 (.A(rst_reg_n), .B(n32022), .C(n32021), 
         .D(n31958), .Z(n26036)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_2_lut_4_lut_4_lut_adj_585.init = 16'hfffd;
    LUT4 i1_4_lut_4_lut_adj_586 (.A(rst_reg_n), .B(instr_complete_N_1647), 
         .C(n28276), .D(n31883), .Z(clk_c_enable_115)) /* synthesis lut_function=((B (C+(D))+!B (D))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_4_lut_4_lut_adj_586.init = 16'hffd5;
    LUT4 i1_3_lut_4_lut_4_lut_adj_587 (.A(rst_reg_n), .B(n31902), .C(n31925), 
         .D(n32019), .Z(clk_c_enable_334)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_587.init = 16'h555d;
    LUT4 i1_3_lut_rep_512_3_lut (.A(rst_reg_n), .B(stop_txn_reg), .C(stop_txn_now_N_2363), 
         .Z(n31717)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_rep_512_3_lut.init = 16'hfdfd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_588 (.A(rst_reg_n), .B(n80), .C(n18241), 
         .D(clk_c_enable_268), .Z(clk_c_enable_10)) /* synthesis lut_function=(!(A (B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(205[13:23])
    defparam i1_3_lut_4_lut_4_lut_adj_588.init = 16'h5755;
    CCU2C cycle_counter_12__I_0_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23551), .S0(mid_bit));
    defparam cycle_counter_12__I_0_13.INIT0 = 16'h0000;
    defparam cycle_counter_12__I_0_13.INIT1 = 16'h0000;
    defparam cycle_counter_12__I_0_13.INJECT1_0 = "NO";
    defparam cycle_counter_12__I_0_13.INJECT1_1 = "NO";
    LUT4 i1_4_lut_rep_846 (.A(fsm_state[2]), .B(fsm_state[0]), .C(fsm_state[1]), 
         .D(fsm_state[3]), .Z(n32051)) /* synthesis lut_function=(!(A+!(B (C (D))+!B (C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_rep_846.init = 16'h5001;
    LUT4 i27947_2_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(fsm_state[1]), 
         .D(fsm_state[3]), .Z(n29255)) /* synthesis lut_function=(A+(B+!(C (D)+!C !(D)))) */ ;
    defparam i27947_2_lut_4_lut.init = 16'heffe;
    PFUMX mux_3032_i1 (.BLUT(n5252[0]), .ALUT(n5272[0]), .C0(n29255), 
          .Z(next_fsm_state[0]));
    LUT4 next_bit_bdd_4_lut (.A(next_bit), .B(fsm_state[1]), .C(fsm_state[3]), 
         .D(fsm_state[2]), .Z(uart_rx_data_7__N_3059)) /* synthesis lut_function=(!((B (C)+!B (C (D)+!C !(D)))+!A)) */ ;
    defparam next_bit_bdd_4_lut.init = 16'h0a28;
    PFUMX i28630 (.BLUT(n32090), .ALUT(n32091), .C0(fsm_state[2]), .Z(next_fsm_state[3]));
    
endmodule
//
// Verilog Description of module led
//

module led (led_out, clk_c, clk_c_enable_268, clk_c_enable_445, n29201) /* synthesis syn_module_defined=1 */ ;
    output led_out;
    input clk_c;
    input clk_c_enable_268;
    input clk_c_enable_445;
    input n29201;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    FD1P3BX led_14 (.D(n29201), .SP(clk_c_enable_268), .CK(clk_c), .PD(clk_c_enable_445), 
            .Q(led_out)) /* synthesis LSE_LINE_FILE_ID=11, LSE_LCOL=6, LSE_RCOL=3, LSE_LLINE=217, LSE_RLINE=229 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/led.v(21[7] 22[21])
    defparam led_14.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module tinyQV
//

module tinyQV (rst_reg_n_adj_17, clk_c, rst_reg_n, data_out_hold, data_ready_r_N_2792, 
            n31883, clk_c_enable_387, \addr[10] , n26205, n8819, \addr[8] , 
            clk_c_enable_36, n31958, n28276, n26216, n31936, clk_c_enable_395, 
            \addr[2] , \addr[9] , n32033, n10467, n31934, n31880, 
            data_ready_r, n18241, n31977, n26036, data_stall, n29198, 
            n31930, clk_c_enable_445, is_writing, stop_txn_now_N_2363, 
            n31713, \instr_addr_23__N_318[7] , \instr_addr_23__N_318[11] , 
            instr_active_N_2106, \instr_addr_23__N_318[9] , \instr_addr_23__N_318[12] , 
            n10500, \instr_addr_23__N_318[13] , \instr_addr_23__N_318[3] , 
            \addr[4] , \instr_addr_23__N_318[22] , \instr_addr_23__N_318[10] , 
            \instr_addr_23__N_318[4] , \addr[5] , \instr_data[15] , \instr_data[13] , 
            \instr_addr_23__N_318[8] , \instr_addr_23__N_318[6] , \addr[7] , 
            \instr_addr_23__N_318[5] , \addr[6] , \instr_addr_23__N_318[14] , 
            \instr_addr_23__N_318[15] , \instr_addr_23__N_318[16] , \instr_addr_23__N_318[17] , 
            \instr_addr_23__N_318[18] , \instr_addr_23__N_318[19] , \instr_addr_23__N_318[20] , 
            \instr_addr_23__N_318[21] , \instr_addr_23__N_318[2] , \addr[3] , 
            \instr_addr[1] , data_stall_N_2158, continue_txn_N_2131, n10499, 
            data_to_write, \data_to_write[12] , \data_to_write[11] , \data_to_write[10] , 
            \data_to_write[9] , \data_to_write[8] , \data_to_write[7] , 
            \data_to_write[6] , \data_to_write[5] , \data_to_write[4] , 
            \data_to_write[3] , \data_to_write[2] , \data_to_write[1] , 
            n31716, is_writing_N_2331, n33479, fsm_state, clk_c_enable_231, 
            n31717, clk_c_enable_186, qspi_ram_b_select, clk_c_enable_239, 
            qspi_ram_a_select, n29199, \qspi_data_out_3__N_5[0] , \nibbles_remaining[0] , 
            n32077, clk_c_enable_452, n31906, n6228, n1084, \writing_N_164[3] , 
            n31971, n27464, clk_N_45, \qspi_data_out_3__N_5[2] , n27081, 
            \qspi_data_oe[0] , clk_c_enable_324, stop_txn_reg, n8135, 
            debug_stop_txn, n31950, \qspi_data_in[0] , \qspi_data_out_3__N_5[3] , 
            \qspi_data_in_3__N_1[0] , \addr[21] , spi_clk_pos_derived_59, 
            qspi_clk_N_56, n31712, n27030, n8, n3, n6232, n27620, 
            n27183, \qspi_data_in[2] , \qspi_data_in[3] , \instr_addr_23__N_318[0] , 
            n31593, \data_from_read[2] , counter_hi, was_early_branch, 
            \rd[0] , \rs1[0] , \addr[27] , \instr_write_offset[3] , 
            n31860, rs2, \instr_len[2] , n31869, debug_instr_valid, 
            \pc[1] , \pc[2] , n2565, n2208, n31742, \data_out_slice[3] , 
            n31879, n19, n31885, \peri_data_out[9] , n4, n31865, 
            n31944, n2524, n2504, VCC_net, n31997, n31902, \pc[5] , 
            \pc[13] , n28964, \peri_data_out[6] , n31867, n4_adj_18, 
            n4263, \pc[9] , \imm[23] , \imm[22] , \imm[21] , \imm[20] , 
            \imm[19] , \imm[18] , \imm[17] , \imm[16] , \imm[15] , 
            \imm[14] , \imm[13] , \imm[12] , \imm[11] , \imm[10] , 
            \imm[9] , \imm[8] , \imm[7] , \imm[6] , \imm[5] , \imm[4] , 
            \imm[3] , \imm[2] , \imm[1] , n32035, n32019, n31900, 
            n26266, n31901, n80, n31868, n31978, n31847, instr_complete_N_1647, 
            n2152, \early_branch_addr[2] , n31863, \instr_data[1][7] , 
            \instr_data[2][7] , n31853, n31849, \instr_data[3][7] , 
            n32055, \debug_rd_3__N_405[31] , \next_pc_for_core[6] , n2136, 
            n2514, \next_pc_for_core[4] , \next_pc_for_core[9] , \next_pc_for_core[13] , 
            \next_pc_for_core[10] , \next_pc_for_core[14] , \peri_data_out[10] , 
            n31761, \cycle[0] , data_out_3__N_1385, is_ret_de, n32027, 
            clk_c_enable_268, \next_pc_for_core[8] , \next_pc_for_core[12] , 
            n31905, n28760, \next_pc_for_core[3] , \pc[23] , \pc[22] , 
            \pc[21] , \pc[20] , \pc[19] , \pc[18] , \pc[17] , \pc[16] , 
            \pc[15] , \pc[14] , \pc[12] , \pc[11] , \pc[10] , \pc[8] , 
            \pc[7] , \next_pc_for_core[5] , \pc[6] , \pc[4] , \next_pc_for_core[7] , 
            n84, \next_pc_for_core[11] , \next_pc_for_core[15] , \pc[3] , 
            \early_branch_addr[5] , n32016, \next_pc_for_core[16] , \early_branch_addr[6] , 
            \next_pc_for_core[17] , \next_pc_for_core[18] , \next_pc_for_core[19] , 
            \next_pc_for_core[20] , \early_branch_addr[4] , \early_branch_addr[3] , 
            \early_branch_addr[7] , \early_branch_addr[8] , \early_branch_addr[9] , 
            \early_branch_addr[10] , \next_pc_for_core[21] , \early_branch_addr[11] , 
            \early_branch_addr[12] , \early_branch_addr[13] , \early_branch_addr[14] , 
            \early_branch_addr[15] , \next_pc_for_core[22] , \early_branch_addr[16] , 
            \early_branch_addr[17] , \next_pc_for_core[23] , n32034, \gpio_out_sel_7__N_13[0] , 
            \early_branch_addr[18] , \early_branch_addr[19] , \early_branch_addr[20] , 
            \early_branch_addr[21] , \early_branch_addr[22] , \early_branch_addr[23] , 
            n31864, n1724, n31935, n32021, n32022, n31962, n31925, 
            n31927, n26282, n31964, n31967, n31735, n31164, n32017, 
            n31163, clk_c_enable_390, \data_from_read[7] , \data_from_read[3] , 
            \data_from_read[0] , \data_from_read[4] , \data_from_read[8] , 
            \data_from_read[12] , \data_from_read[1] , \data_from_read[5] , 
            n31932, n31922, n31819, \peri_data_out[11] , gpio_out_sel, 
            n14, n14_adj_19, n31961, n5171, n28686, clk_c_enable_273, 
            clk_c_enable_357, clk_c_enable_349, n32003, clk_c_enable_259, 
            clk_c_enable_360, n31904, n10573, n31841, n15604, n29004, 
            n31798, clk_c_enable_234, \ui_in_sync[0] , n1160, \alu_b_in[3] , 
            debug_rd, \ui_in_sync[1] , \next_fsm_state_3__N_3015[3] , 
            fsm_state_adj_25, accum, d_3__N_1868, n31929, \mul_out[1] , 
            \mul_out[2] , \mul_out[3] , n31963, next_bit, n28800, 
            n31389, alu_b_in_3__N_1504, n29162, n18086, \csr_read_3__N_1447[2] , 
            GND_net, \next_accum[5] , \next_accum[6] , \next_accum[7] , 
            \next_accum[8] , \next_accum[9] , \next_accum[10] , \next_accum[11] , 
            \next_accum[12] , \next_accum[13] , \next_accum[14] , \next_accum[15] , 
            \next_accum[16] , \next_accum[17] , \next_accum[18] , \next_accum[19] , 
            \next_accum[4] , n12, n11, n9, n8_adj_23, \registers[5][7] , 
            \registers[6][7] , \registers[7][7] , n29747, n4_adj_24) /* synthesis syn_module_defined=1 */ ;
    output rst_reg_n_adj_17;
    input clk_c;
    input rst_reg_n;
    input data_out_hold;
    output data_ready_r_N_2792;
    output n31883;
    output clk_c_enable_387;
    output \addr[10] ;
    output n26205;
    input n8819;
    output \addr[8] ;
    output clk_c_enable_36;
    output n31958;
    output n28276;
    output n26216;
    output n31936;
    output clk_c_enable_395;
    output \addr[2] ;
    output \addr[9] ;
    output n32033;
    output n10467;
    input n31934;
    output n31880;
    input data_ready_r;
    input n18241;
    output n31977;
    input n26036;
    output data_stall;
    input n29198;
    input n31930;
    input clk_c_enable_445;
    output is_writing;
    output stop_txn_now_N_2363;
    output n31713;
    input \instr_addr_23__N_318[7] ;
    input \instr_addr_23__N_318[11] ;
    input instr_active_N_2106;
    input \instr_addr_23__N_318[9] ;
    input \instr_addr_23__N_318[12] ;
    input n10500;
    input \instr_addr_23__N_318[13] ;
    input \instr_addr_23__N_318[3] ;
    output \addr[4] ;
    input \instr_addr_23__N_318[22] ;
    input \instr_addr_23__N_318[10] ;
    input \instr_addr_23__N_318[4] ;
    output \addr[5] ;
    output \instr_data[15] ;
    output \instr_data[13] ;
    input \instr_addr_23__N_318[8] ;
    input \instr_addr_23__N_318[6] ;
    output \addr[7] ;
    input \instr_addr_23__N_318[5] ;
    output \addr[6] ;
    input \instr_addr_23__N_318[14] ;
    input \instr_addr_23__N_318[15] ;
    input \instr_addr_23__N_318[16] ;
    input \instr_addr_23__N_318[17] ;
    input \instr_addr_23__N_318[18] ;
    input \instr_addr_23__N_318[19] ;
    input \instr_addr_23__N_318[20] ;
    input \instr_addr_23__N_318[21] ;
    input \instr_addr_23__N_318[2] ;
    output \addr[3] ;
    input \instr_addr[1] ;
    output data_stall_N_2158;
    output continue_txn_N_2131;
    output n10499;
    output [31:0]data_to_write;
    output \data_to_write[12] ;
    output \data_to_write[11] ;
    output \data_to_write[10] ;
    output \data_to_write[9] ;
    output \data_to_write[8] ;
    output \data_to_write[7] ;
    output \data_to_write[6] ;
    output \data_to_write[5] ;
    output \data_to_write[4] ;
    output \data_to_write[3] ;
    output \data_to_write[2] ;
    output \data_to_write[1] ;
    output n31716;
    output is_writing_N_2331;
    output n33479;
    output [2:0]fsm_state;
    input clk_c_enable_231;
    input n31717;
    input clk_c_enable_186;
    output qspi_ram_b_select;
    input clk_c_enable_239;
    output qspi_ram_a_select;
    input n29199;
    input \qspi_data_out_3__N_5[0] ;
    output \nibbles_remaining[0] ;
    output n32077;
    input clk_c_enable_452;
    output n31906;
    output n6228;
    output n1084;
    output \writing_N_164[3] ;
    output n31971;
    output n27464;
    input clk_N_45;
    input \qspi_data_out_3__N_5[2] ;
    input n27081;
    output \qspi_data_oe[0] ;
    input clk_c_enable_324;
    output stop_txn_reg;
    input n8135;
    output debug_stop_txn;
    input n31950;
    input \qspi_data_in[0] ;
    input \qspi_data_out_3__N_5[3] ;
    output \qspi_data_in_3__N_1[0] ;
    output \addr[21] ;
    output spi_clk_pos_derived_59;
    output qspi_clk_N_56;
    output n31712;
    output n27030;
    output n8;
    output n3;
    output n6232;
    output n27620;
    output n27183;
    input \qspi_data_in[2] ;
    input \qspi_data_in[3] ;
    output \instr_addr_23__N_318[0] ;
    input n31593;
    input \data_from_read[2] ;
    output [4:2]counter_hi;
    output was_early_branch;
    output \rd[0] ;
    output \rs1[0] ;
    output \addr[27] ;
    output \instr_write_offset[3] ;
    output n31860;
    output [3:0]rs2;
    output \instr_len[2] ;
    output n31869;
    output debug_instr_valid;
    output \pc[1] ;
    output \pc[2] ;
    output n2565;
    output n2208;
    output n31742;
    input \data_out_slice[3] ;
    output n31879;
    output n19;
    output n31885;
    input \peri_data_out[9] ;
    output n4;
    output n31865;
    output n31944;
    input n2524;
    input n2504;
    input VCC_net;
    output n31997;
    output n31902;
    output \pc[5] ;
    output \pc[13] ;
    input n28964;
    input \peri_data_out[6] ;
    output n31867;
    input n4_adj_18;
    output n4263;
    output \pc[9] ;
    output \imm[23] ;
    output \imm[22] ;
    output \imm[21] ;
    output \imm[20] ;
    output \imm[19] ;
    output \imm[18] ;
    output \imm[17] ;
    output \imm[16] ;
    output \imm[15] ;
    output \imm[14] ;
    output \imm[13] ;
    output \imm[12] ;
    output \imm[11] ;
    output \imm[10] ;
    output \imm[9] ;
    output \imm[8] ;
    output \imm[7] ;
    output \imm[6] ;
    output \imm[5] ;
    output \imm[4] ;
    output \imm[3] ;
    output \imm[2] ;
    output \imm[1] ;
    output n32035;
    output n32019;
    output n31900;
    output n26266;
    output n31901;
    output n80;
    output n31868;
    output n31978;
    output n31847;
    output instr_complete_N_1647;
    input n2152;
    input \early_branch_addr[2] ;
    output n31863;
    output \instr_data[1][7] ;
    output \instr_data[2][7] ;
    output n31853;
    output n31849;
    output \instr_data[3][7] ;
    output n32055;
    output \debug_rd_3__N_405[31] ;
    input \next_pc_for_core[6] ;
    output n2136;
    output n2514;
    input \next_pc_for_core[4] ;
    input \next_pc_for_core[9] ;
    input \next_pc_for_core[13] ;
    input \next_pc_for_core[10] ;
    input \next_pc_for_core[14] ;
    input \peri_data_out[10] ;
    input n31761;
    output \cycle[0] ;
    output data_out_3__N_1385;
    input is_ret_de;
    input n32027;
    output clk_c_enable_268;
    input \next_pc_for_core[8] ;
    input \next_pc_for_core[12] ;
    input n31905;
    output n28760;
    input \next_pc_for_core[3] ;
    output \pc[23] ;
    output \pc[22] ;
    output \pc[21] ;
    output \pc[20] ;
    output \pc[19] ;
    output \pc[18] ;
    output \pc[17] ;
    output \pc[16] ;
    output \pc[15] ;
    output \pc[14] ;
    output \pc[12] ;
    output \pc[11] ;
    output \pc[10] ;
    output \pc[8] ;
    output \pc[7] ;
    input \next_pc_for_core[5] ;
    output \pc[6] ;
    output \pc[4] ;
    input \next_pc_for_core[7] ;
    input n84;
    input \next_pc_for_core[11] ;
    input \next_pc_for_core[15] ;
    output \pc[3] ;
    input \early_branch_addr[5] ;
    input n32016;
    input \next_pc_for_core[16] ;
    input \early_branch_addr[6] ;
    input \next_pc_for_core[17] ;
    input \next_pc_for_core[18] ;
    input \next_pc_for_core[19] ;
    input \next_pc_for_core[20] ;
    input \early_branch_addr[4] ;
    input \early_branch_addr[3] ;
    input \early_branch_addr[7] ;
    input \early_branch_addr[8] ;
    input \early_branch_addr[9] ;
    input \early_branch_addr[10] ;
    input \next_pc_for_core[21] ;
    input \early_branch_addr[11] ;
    input \early_branch_addr[12] ;
    input \early_branch_addr[13] ;
    input \early_branch_addr[14] ;
    input \early_branch_addr[15] ;
    input \next_pc_for_core[22] ;
    input \early_branch_addr[16] ;
    input \early_branch_addr[17] ;
    input \next_pc_for_core[23] ;
    output n32034;
    output \gpio_out_sel_7__N_13[0] ;
    input \early_branch_addr[18] ;
    input \early_branch_addr[19] ;
    input \early_branch_addr[20] ;
    input \early_branch_addr[21] ;
    input \early_branch_addr[22] ;
    input \early_branch_addr[23] ;
    input n31864;
    input n1724;
    output n31935;
    output n32021;
    output n32022;
    output n31962;
    output n31925;
    output n31927;
    input n26282;
    output n31964;
    output n31967;
    output n31735;
    input n31164;
    input n32017;
    output n31163;
    output clk_c_enable_390;
    input \data_from_read[7] ;
    input \data_from_read[3] ;
    input \data_from_read[0] ;
    input \data_from_read[4] ;
    input \data_from_read[8] ;
    input \data_from_read[12] ;
    input \data_from_read[1] ;
    input \data_from_read[5] ;
    output n31932;
    input n31922;
    output n31819;
    input \peri_data_out[11] ;
    input [7:6]gpio_out_sel;
    output n14;
    output n14_adj_19;
    input n31961;
    output n5171;
    input n28686;
    output clk_c_enable_273;
    output clk_c_enable_357;
    output clk_c_enable_349;
    input n32003;
    output clk_c_enable_259;
    output clk_c_enable_360;
    output n31904;
    input n10573;
    output n31841;
    output n15604;
    output n29004;
    output n31798;
    input clk_c_enable_234;
    input \ui_in_sync[0] ;
    output n1160;
    input \alu_b_in[3] ;
    output [3:0]debug_rd;
    input \ui_in_sync[1] ;
    input \next_fsm_state_3__N_3015[3] ;
    input [3:0]fsm_state_adj_25;
    output [15:0]accum;
    output [19:0]d_3__N_1868;
    output n31929;
    input \mul_out[1] ;
    input \mul_out[2] ;
    input \mul_out[3] ;
    output n31963;
    input next_bit;
    output n28800;
    input n31389;
    output alu_b_in_3__N_1504;
    input n29162;
    output n18086;
    output \csr_read_3__N_1447[2] ;
    input GND_net;
    input \next_accum[5] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[4] ;
    output n12;
    output n11;
    output n9;
    output n8_adj_23;
    output \registers[5][7] ;
    output \registers[6][7] ;
    output \registers[7][7] ;
    output n29747;
    input n4_adj_24;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    
    wire n33488, stall_core, is_load, n28928, n28788;
    wire [1:0]qv_data_write_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(64[15:30])
    
    wire n18680, data_ready, n31899, n32006, n31940, n31862, qspi_write_done, 
        n31907, n31908, n31887;
    wire [1:0]data_txn_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(49[15:27])
    wire [15:0]instr_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(61[15:25])
    wire [31:0]mem_data_from_read;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(74[15:33])
    wire [31:0]qspi_data_buf;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(58[16:29])
    
    wire debug_data_continue, instr_active, start_instr, instr_fetch_stopped;
    wire [27:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    
    wire instr_fetch_running_N_945, n31730, mem_data_ready;
    wire [23:1]instr_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(56[15:25])
    
    wire qspi_data_ready;
    wire [1:0]txn_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(56[16:23])
    
    wire debug_stop_txn_N_2147, n58, n18588, n31939, n31941;
    wire [31:0]data_to_write_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(56[17:30])
    
    wire n32052, n31792, n27702, n13146, n31725, n27310, n31741, 
        n8_c, n27762, instr_fetch_running_N_943, n31770, instr_fetch_running, 
        n31942, n31736, n1176, n32020, n27680, n31910, n31994, 
        n27776, n31991, n27772, n31990, n27780;
    
    FD1S3AX rst_reg_n_16 (.D(rst_reg_n), .CK(clk_c), .Q(rst_reg_n_adj_17)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=111, LSE_RLINE=150 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(92[10:43])
    defparam rst_reg_n_16.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_678 (.A(data_out_hold), .B(data_ready_r_N_2792), .Z(n31883)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_rep_678.init = 16'h4444;
    LUT4 i444_2_lut_3_lut (.A(data_out_hold), .B(data_ready_r_N_2792), .C(rst_reg_n), 
         .Z(clk_c_enable_387)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i444_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_4_lut (.A(\addr[10] ), .B(n26205), .C(n8819), .D(\addr[8] ), 
         .Z(data_ready_r_N_2792)) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_4_lut.init = 16'h88c8;
    FD1S3AX rst_reg_n_16_rep_862 (.D(rst_reg_n), .CK(clk_c), .Q(n33488)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=12, LSE_RCOL=6, LSE_LLINE=111, LSE_RLINE=150 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(92[10:43])
    defparam rst_reg_n_16_rep_862.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_568 (.A(stall_core), .B(clk_c_enable_36), .C(n31958), 
         .D(is_load), .Z(n28276)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(86[31:66])
    defparam i1_4_lut_adj_568.init = 16'h8000;
    LUT4 i1_4_lut_adj_569 (.A(n26216), .B(n31936), .C(n28928), .D(n28788), 
         .Z(clk_c_enable_395)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_569.init = 16'h0200;
    LUT4 i26370_2_lut (.A(\addr[2] ), .B(\addr[9] ), .Z(n28928)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26370_2_lut.init = 16'heeee;
    LUT4 i1_3_lut (.A(\addr[10] ), .B(qv_data_write_n[1]), .C(qv_data_write_n[0]), 
         .Z(n28788)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;
    defparam i1_3_lut.init = 16'h1414;
    LUT4 i1_2_lut_rep_675_3_lut_4_lut (.A(n31958), .B(n32033), .C(n10467), 
         .D(n31934), .Z(n31880)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_2_lut_rep_675_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_3_lut_4_lut (.A(n31958), .B(n32033), .C(data_ready_r), .D(n18680), 
         .Z(data_ready)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_3_lut_4_lut.init = 16'hf2ff;
    LUT4 i1_3_lut_rep_694_4_lut (.A(n31958), .B(n32033), .C(n18241), .D(rst_reg_n), 
         .Z(n31899)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(76[17:41])
    defparam i1_3_lut_rep_694_4_lut.init = 16'h0222;
    LUT4 i26386_2_lut_rep_657_3_lut_4_lut_3_lut_4_lut_4_lut (.A(n31958), .B(n32006), 
         .C(n31940), .D(n32033), .Z(n31862)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i26386_2_lut_rep_657_3_lut_4_lut_3_lut_4_lut_4_lut.init = 16'hfefa;
    LUT4 i5555_2_lut_rep_702_3_lut_4_lut (.A(n31958), .B(n32006), .C(qspi_write_done), 
         .D(n31977), .Z(n31907)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;
    defparam i5555_2_lut_rep_702_3_lut_4_lut.init = 16'hfff1;
    LUT4 i15669_2_lut_rep_703_3_lut_4_lut (.A(n31958), .B(n32006), .C(qspi_write_done), 
         .D(n31977), .Z(n31908)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15669_2_lut_rep_703_3_lut_4_lut.init = 16'hfffe;
    LUT4 i15942_2_lut_rep_682_3_lut_4_lut_4_lut (.A(n31958), .B(n32006), 
         .C(n31940), .D(n32033), .Z(n31887)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i15942_2_lut_rep_682_3_lut_4_lut_4_lut.init = 16'hfffb;
    tinyqv_mem_ctrl mem (.clk_c(clk_c), .data_txn_len({data_txn_len}), .n26036(n26036), 
            .qspi_write_done(qspi_write_done), .data_stall(data_stall), 
            .rst_reg_n(rst_reg_n), .n29198(n29198), .instr_data({\instr_data[15] , 
            instr_data[14], \instr_data[13] , instr_data[12:0]}), .\mem_data_from_read[23] (mem_data_from_read[23]), 
            .\mem_data_from_read[22] (mem_data_from_read[22]), .\mem_data_from_read[21] (mem_data_from_read[21]), 
            .\mem_data_from_read[20] (mem_data_from_read[20]), .\mem_data_from_read[19] (mem_data_from_read[19]), 
            .\mem_data_from_read[18] (mem_data_from_read[18]), .\mem_data_from_read[17] (mem_data_from_read[17]), 
            .\mem_data_from_read[16] (mem_data_from_read[16]), .\qspi_data_buf[15] (qspi_data_buf[15]), 
            .\qspi_data_buf[14] (qspi_data_buf[14]), .\qspi_data_buf[13] (qspi_data_buf[13]), 
            .\qspi_data_buf[11] (qspi_data_buf[11]), .\qspi_data_buf[10] (qspi_data_buf[10]), 
            .\qspi_data_buf[9] (qspi_data_buf[9]), .n31930(n31930), .clk_c_enable_445(clk_c_enable_445), 
            .debug_data_continue(debug_data_continue), .instr_active(instr_active), 
            .start_instr(start_instr), .n31940(n31940), .is_writing(is_writing), 
            .stop_txn_now_N_2363(stop_txn_now_N_2363), .n31862(n31862), 
            .n31713(n31713), .instr_fetch_stopped(instr_fetch_stopped), 
            .n31977(n31977), .\instr_addr_23__N_318[7] (\instr_addr_23__N_318[7] ), 
            .\addr[8] (\addr[8] ), .\instr_addr_23__N_318[11] (\instr_addr_23__N_318[11] ), 
            .\addr[12] (addr[12]), .\addr[24] (addr[24]), .instr_active_N_2106(instr_active_N_2106), 
            .\instr_addr_23__N_318[9] (\instr_addr_23__N_318[9] ), .\addr[10] (\addr[10] ), 
            .\instr_addr_23__N_318[12] (\instr_addr_23__N_318[12] ), .\addr[13] (addr[13]), 
            .instr_fetch_running_N_945(instr_fetch_running_N_945), .n10500(n10500), 
            .n31730(n31730), .\instr_addr_23__N_318[13] (\instr_addr_23__N_318[13] ), 
            .\addr[14] (addr[14]), .\instr_addr_23__N_318[3] (\instr_addr_23__N_318[3] ), 
            .\addr[4] (\addr[4] ), .\instr_addr_23__N_318[22] (\instr_addr_23__N_318[22] ), 
            .\addr[23] (addr[23]), .\instr_addr_23__N_318[10] (\instr_addr_23__N_318[10] ), 
            .\addr[11] (addr[11]), .\instr_addr_23__N_318[4] (\instr_addr_23__N_318[4] ), 
            .\addr[5] (\addr[5] ), .mem_data_ready(mem_data_ready), .\mem_data_from_read[31] (mem_data_from_read[31]), 
            .\mem_data_from_read[27] (mem_data_from_read[27]), .\mem_data_from_read[30] (mem_data_from_read[30]), 
            .\mem_data_from_read[26] (mem_data_from_read[26]), .\mem_data_from_read[29] (mem_data_from_read[29]), 
            .\mem_data_from_read[25] (mem_data_from_read[25]), .\mem_data_from_read[28] (mem_data_from_read[28]), 
            .\mem_data_from_read[24] (mem_data_from_read[24]), .\instr_addr_23__N_318[8] (\instr_addr_23__N_318[8] ), 
            .\addr[9] (\addr[9] ), .\instr_addr_23__N_318[6] (\instr_addr_23__N_318[6] ), 
            .\addr[7] (\addr[7] ), .\instr_addr_23__N_318[5] (\instr_addr_23__N_318[5] ), 
            .\addr[6] (\addr[6] ), .\instr_addr_23__N_318[14] (\instr_addr_23__N_318[14] ), 
            .\addr[15] (addr[15]), .\instr_addr_23__N_318[15] (\instr_addr_23__N_318[15] ), 
            .\addr[16] (addr[16]), .\instr_addr_23__N_318[16] (\instr_addr_23__N_318[16] ), 
            .\addr[17] (addr[17]), .\instr_addr_23__N_318[17] (\instr_addr_23__N_318[17] ), 
            .\addr[18] (addr[18]), .\instr_addr_23__N_318[18] (\instr_addr_23__N_318[18] ), 
            .\addr[19] (addr[19]), .\instr_addr_23__N_318[19] (\instr_addr_23__N_318[19] ), 
            .\addr[20] (addr[20]), .\instr_addr_23__N_318[20] (\instr_addr_23__N_318[20] ), 
            .\addr[21] (addr[21]), .\instr_addr_23__N_318[21] (\instr_addr_23__N_318[21] ), 
            .\addr[22] (addr[22]), .\instr_addr_23__N_318[2] (\instr_addr_23__N_318[2] ), 
            .\addr[3] (\addr[3] ), .\instr_addr[2] (instr_addr[2]), .\addr[2] (\addr[2] ), 
            .\instr_addr[1] (\instr_addr[1] ), .\addr[1] (addr[1]), .qspi_data_ready(qspi_data_ready), 
            .\txn_len[1] (txn_len[1]), .n31958(n31958), .debug_stop_txn_N_2147(debug_stop_txn_N_2147), 
            .n58(n58), .n18588(n18588), .n31939(n31939), .data_stall_N_2158(data_stall_N_2158), 
            .n31941(n31941), .continue_txn_N_2131(continue_txn_N_2131), 
            .n10499(n10499), .n31908(n31908), .n31887(n31887), .data_to_write({data_to_write_c[31:13], 
            \data_to_write[12] , \data_to_write[11] , \data_to_write[10] , 
            \data_to_write[9] , \data_to_write[8] , \data_to_write[7] , 
            \data_to_write[6] , \data_to_write[5] , \data_to_write[4] , 
            \data_to_write[3] , \data_to_write[2] , \data_to_write[1] , 
            data_to_write[0]}), .n32052(n32052), .n31792(n31792), .\mem_data_from_read[5] (mem_data_from_read[5]), 
            .n31716(n31716), .n27702(n27702), .n13146(n13146), .\mem_data_from_read[1] (mem_data_from_read[1]), 
            .\mem_data_from_read[4] (mem_data_from_read[4]), .\mem_data_from_read[0] (mem_data_from_read[0]), 
            .\mem_data_from_read[3] (mem_data_from_read[3]), .\mem_data_from_read[7] (mem_data_from_read[7]), 
            .n31725(n31725), .is_writing_N_2331(is_writing_N_2331), .n33479(n33479), 
            .\mem_data_from_read[12] (mem_data_from_read[12]), .n27310(n27310), 
            .\mem_data_from_read[8] (mem_data_from_read[8]), .n31741(n31741), 
            .n8(n8_c), .n27762(n27762), .instr_fetch_running_N_943(instr_fetch_running_N_943), 
            .n31907(n31907), .\addr[0] (addr[0]), .n31770(n31770), .fsm_state({fsm_state}), 
            .clk_c_enable_231(clk_c_enable_231), .n31717(n31717), .clk_c_enable_186(clk_c_enable_186), 
            .qspi_ram_b_select(qspi_ram_b_select), .clk_c_enable_239(clk_c_enable_239), 
            .qspi_ram_a_select(qspi_ram_a_select), .n29199(n29199), .\qspi_data_out_3__N_5[0] (\qspi_data_out_3__N_5[0] ), 
            .\nibbles_remaining[0] (\nibbles_remaining[0] ), .n32077(n32077), 
            .clk_c_enable_452(clk_c_enable_452), .n31906(n31906), .n6228(n6228), 
            .n1084(n1084), .\writing_N_164[3] (\writing_N_164[3] ), .n31971(n31971), 
            .n27464(n27464), .clk_N_45(clk_N_45), .\qspi_data_out_3__N_5[2] (\qspi_data_out_3__N_5[2] ), 
            .n27081(n27081), .\qspi_data_oe[0] (\qspi_data_oe[0] ), .clk_c_enable_324(clk_c_enable_324), 
            .stop_txn_reg(stop_txn_reg), .n8135(n8135), .instr_fetch_running(instr_fetch_running), 
            .n31942(n31942), .debug_stop_txn(debug_stop_txn), .n31950(n31950), 
            .\qspi_data_in[0] (\qspi_data_in[0] ), .\qspi_data_out_3__N_5[3] (\qspi_data_out_3__N_5[3] ), 
            .\qspi_data_in_3__N_1[0] (\qspi_data_in_3__N_1[0] ), .\addr[21]_adj_15 (\addr[21] ), 
            .n31736(n31736), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .qspi_clk_N_56(qspi_clk_N_56), .n31712(n31712), .n1176(n1176), 
            .n27030(n27030), .n8_adj_16(n8), .n3(n3), .n6232(n6232), 
            .n27620(n27620), .n27183(n27183), .\qspi_data_in[2] (\qspi_data_in[2] ), 
            .\qspi_data_in[3] (\qspi_data_in[3] ), .n32020(n32020), .n27680(n27680), 
            .\instr_addr_23__N_318[0] (\instr_addr_23__N_318[0] ), .n31910(n31910), 
            .n31994(n31994), .n27776(n27776), .n31991(n31991), .n27772(n27772), 
            .n31990(n31990), .n27780(n27780), .n31593(n31593)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(132[19] 164[6])
    tinyqv_cpu cpu (.clk_c(clk_c), .\data_from_read[2] (\data_from_read[2] ), 
            .counter_hi({counter_hi}), .was_early_branch(was_early_branch), 
            .data_to_write({data_to_write_c[31:13], \data_to_write[12] , 
            \data_to_write[11] , \data_to_write[10] , \data_to_write[9] , 
            \data_to_write[8] , \data_to_write[7] , \data_to_write[6] , 
            \data_to_write[5] , \data_to_write[4] , \data_to_write[3] , 
            \data_to_write[2] , \data_to_write[1] , data_to_write[0]}), 
            .qv_data_write_n({qv_data_write_n}), .rd({Open_38, Open_39, 
            Open_40, \rd[0] }), .rs1({Open_41, Open_42, Open_43, \rs1[0] }), 
            .\instr_addr_23__N_318[0] (\instr_addr_23__N_318[0] ), .addr({\addr[27] , 
            Open_44, Open_45, Open_46, Open_47, Open_48, Open_49, 
            Open_50, Open_51, Open_52, Open_53, Open_54, Open_55, 
            Open_56, Open_57, Open_58, Open_59, Open_60, Open_61, 
            Open_62, Open_63, Open_64, Open_65, Open_66, Open_67, 
            Open_68, Open_69, addr[0]}), .\addr[24] (addr[24]), .\addr[23] (addr[23]), 
            .\addr[22] (addr[22]), .\addr[21] (addr[21]), .\addr[20] (addr[20]), 
            .\addr[19] (addr[19]), .\addr[18] (addr[18]), .\addr[17] (addr[17]), 
            .\addr[16] (addr[16]), .\addr[15] (addr[15]), .\addr[14] (addr[14]), 
            .\addr[13] (addr[13]), .\addr[12] (addr[12]), .\addr[11] (addr[11]), 
            .\addr[10] (\addr[10] ), .\addr[9] (\addr[9] ), .\addr[8] (\addr[8] ), 
            .\addr[7] (\addr[7] ), .\addr[6] (\addr[6] ), .\addr[5] (\addr[5] ), 
            .\addr[4] (\addr[4] ), .\addr[3] (\addr[3] ), .\addr[2] (\addr[2] ), 
            .\addr[1] (addr[1]), .\instr_write_offset[3] (\instr_write_offset[3] ), 
            .debug_data_continue(debug_data_continue), .is_load(is_load), 
            .n31860(n31860), .rs2({rs2}), .\instr_len[2] (\instr_len[2] ), 
            .n31869(n31869), .debug_instr_valid(debug_instr_valid), .\pc[1] (\pc[1] ), 
            .\pc[2] (\pc[2] ), .n2565(n2565), .n31770(n31770), .n2208(n2208), 
            .n31742(n31742), .\data_out_slice[3] (\data_out_slice[3] ), 
            .n31879(n31879), .n19(n19), .n31885(n31885), .\peri_data_out[9] (\peri_data_out[9] ), 
            .n4(n4), .\mem_data_from_read[20] (mem_data_from_read[20]), 
            .\mem_data_from_read[16] (mem_data_from_read[16]), .n31865(n31865), 
            .n31944(n31944), .n2524(n2524), .n2504(n2504), .n31958(n31958), 
            .VCC_net(VCC_net), .rst_reg_n(rst_reg_n_adj_17), .n31792(n31792), 
            .data_txn_len({data_txn_len}), .instr_data({\instr_data[15] , 
            instr_data[14], \instr_data[13] , instr_data[12:0]}), .n31997(n31997), 
            .n18241(n18241), .n32033(n32033), .n31902(n31902), .\pc[5] (\pc[5] ), 
            .\pc[13] (\pc[13] ), .n28964(n28964), .n10467(n10467), .\peri_data_out[6] (\peri_data_out[6] ), 
            .n31867(n31867), .n4_adj_11(n4_adj_18), .n26216(n26216), .n4263(n4263), 
            .\pc[9] (\pc[9] ), .\imm[23] (\imm[23] ), .\imm[22] (\imm[22] ), 
            .\imm[21] (\imm[21] ), .\imm[20] (\imm[20] ), .\imm[19] (\imm[19] ), 
            .\imm[18] (\imm[18] ), .\imm[17] (\imm[17] ), .\imm[16] (\imm[16] ), 
            .\imm[15] (\imm[15] ), .\imm[14] (\imm[14] ), .\imm[13] (\imm[13] ), 
            .\imm[12] (\imm[12] ), .\imm[11] (\imm[11] ), .\imm[10] (\imm[10] ), 
            .\imm[9] (\imm[9] ), .\imm[8] (\imm[8] ), .\imm[7] (\imm[7] ), 
            .\imm[6] (\imm[6] ), .\imm[5] (\imm[5] ), .\imm[4] (\imm[4] ), 
            .\imm[3] (\imm[3] ), .\imm[2] (\imm[2] ), .\imm[1] (\imm[1] ), 
            .n33488(n33488), .n10499(n10499), .n31730(n31730), .instr_active(instr_active), 
            .\txn_len[1] (txn_len[1]), .n32035(n32035), .n32019(n32019), 
            .n31900(n31900), .n26266(n26266), .n31901(n31901), .n80(n80), 
            .n31868(n31868), .n31978(n31978), .n31847(n31847), .n27702(n27702), 
            .n13146(n13146), .instr_complete_N_1647(instr_complete_N_1647), 
            .instr_fetch_running(instr_fetch_running), .n2152(n2152), .\early_branch_addr[2] (\early_branch_addr[2] ), 
            .\instr_addr[2] (instr_addr[2]), .n31863(n31863), .\instr_data[1][7] (\instr_data[1][7] ), 
            .\instr_data[2][7] (\instr_data[2][7] ), .n31853(n31853), .debug_stop_txn_N_2147(debug_stop_txn_N_2147), 
            .instr_fetch_running_N_945(instr_fetch_running_N_945), .qspi_data_ready(qspi_data_ready), 
            .n32052(n32052), .n58(n58), .n31849(n31849), .\instr_data[3][7] (\instr_data[3][7] ), 
            .n32055(n32055), .stall_core(stall_core), .start_instr(start_instr), 
            .n31741(n31741), .n8(n8_c), .\debug_rd_3__N_405[31] (\debug_rd_3__N_405[31] ), 
            .\next_pc_for_core[6] (\next_pc_for_core[6] ), .n2136(n2136), 
            .n2514(n2514), .\next_pc_for_core[4] (\next_pc_for_core[4] ), 
            .n31940(n31940), .n32006(n32006), .\next_pc_for_core[9] (\next_pc_for_core[9] ), 
            .\next_pc_for_core[13] (\next_pc_for_core[13] ), .\next_pc_for_core[10] (\next_pc_for_core[10] ), 
            .\next_pc_for_core[14] (\next_pc_for_core[14] ), .\peri_data_out[10] (\peri_data_out[10] ), 
            .n31761(n31761), .\mem_data_from_read[19] (mem_data_from_read[19]), 
            .\mem_data_from_read[23] (mem_data_from_read[23]), .cycle({Open_70, 
            \cycle[0] }), .data_out_3__N_1385(data_out_3__N_1385), .is_ret_de(is_ret_de), 
            .n31990(n31990), .n31991(n31991), .n31994(n31994), .n31939(n31939), 
            .n31934(n31934), .n32027(n32027), .n26205(n26205), .clk_c_enable_268(clk_c_enable_268), 
            .n31941(n31941), .\next_pc_for_core[8] (\next_pc_for_core[8] ), 
            .\next_pc_for_core[12] (\next_pc_for_core[12] ), .data_ready_r(data_ready_r), 
            .n31905(n31905), .n28760(n28760), .\next_pc_for_core[3] (\next_pc_for_core[3] ), 
            .\pc[23] (\pc[23] ), .\pc[22] (\pc[22] ), .\pc[21] (\pc[21] ), 
            .\pc[20] (\pc[20] ), .\pc[19] (\pc[19] ), .\pc[18] (\pc[18] ), 
            .\pc[17] (\pc[17] ), .\pc[16] (\pc[16] ), .\pc[15] (\pc[15] ), 
            .\pc[14] (\pc[14] ), .\pc[12] (\pc[12] ), .\pc[11] (\pc[11] ), 
            .\pc[10] (\pc[10] ), .\pc[8] (\pc[8] ), .\pc[7] (\pc[7] ), 
            .\next_pc_for_core[5] (\next_pc_for_core[5] ), .\pc[6] (\pc[6] ), 
            .\pc[4] (\pc[4] ), .\next_pc_for_core[7] (\next_pc_for_core[7] ), 
            .n84(n84), .\next_pc_for_core[11] (\next_pc_for_core[11] ), 
            .\next_pc_for_core[15] (\next_pc_for_core[15] ), .\pc[3] (\pc[3] ), 
            .\early_branch_addr[5] (\early_branch_addr[5] ), .n32016(n32016), 
            .\next_pc_for_core[16] (\next_pc_for_core[16] ), .\early_branch_addr[6] (\early_branch_addr[6] ), 
            .\next_pc_for_core[17] (\next_pc_for_core[17] ), .\next_pc_for_core[18] (\next_pc_for_core[18] ), 
            .\next_pc_for_core[19] (\next_pc_for_core[19] ), .\next_pc_for_core[20] (\next_pc_for_core[20] ), 
            .\early_branch_addr[4] (\early_branch_addr[4] ), .\early_branch_addr[3] (\early_branch_addr[3] ), 
            .\early_branch_addr[7] (\early_branch_addr[7] ), .\early_branch_addr[8] (\early_branch_addr[8] ), 
            .\early_branch_addr[9] (\early_branch_addr[9] ), .\early_branch_addr[10] (\early_branch_addr[10] ), 
            .\next_pc_for_core[21] (\next_pc_for_core[21] ), .\early_branch_addr[11] (\early_branch_addr[11] ), 
            .\early_branch_addr[12] (\early_branch_addr[12] ), .\early_branch_addr[13] (\early_branch_addr[13] ), 
            .\early_branch_addr[14] (\early_branch_addr[14] ), .\early_branch_addr[15] (\early_branch_addr[15] ), 
            .\next_pc_for_core[22] (\next_pc_for_core[22] ), .\early_branch_addr[16] (\early_branch_addr[16] ), 
            .\early_branch_addr[17] (\early_branch_addr[17] ), .\next_pc_for_core[23] (\next_pc_for_core[23] ), 
            .n32034(n32034), .n31880(n31880), .\gpio_out_sel_7__N_13[0] (\gpio_out_sel_7__N_13[0] ), 
            .n31725(n31725), .\early_branch_addr[18] (\early_branch_addr[18] ), 
            .\early_branch_addr[19] (\early_branch_addr[19] ), .\early_branch_addr[20] (\early_branch_addr[20] ), 
            .\early_branch_addr[21] (\early_branch_addr[21] ), .\early_branch_addr[22] (\early_branch_addr[22] ), 
            .\early_branch_addr[23] (\early_branch_addr[23] ), .n31864(n31864), 
            .n1724(n1724), .n31935(n31935), .n32020(n32020), .n27310(n27310), 
            .n31736(n31736), .n33479(n33479), .n31906(n31906), .n1176(n1176), 
            .n32021(n32021), .n32022(n32022), .n18588(n18588), .clk_c_enable_36(clk_c_enable_36), 
            .mem_data_ready(mem_data_ready), .data_ready(data_ready), .n31936(n31936), 
            .n31962(n31962), .n31925(n31925), .n31927(n31927), .n26282(n26282), 
            .n31964(n31964), .n31967(n31967), .n31735(n31735), .n31164(n31164), 
            .n27680(n27680), .n32017(n32017), .n31163(n31163), .clk_c_enable_390(clk_c_enable_390), 
            .\mem_data_from_read[7] (mem_data_from_read[7]), .\data_from_read[7] (\data_from_read[7] ), 
            .\mem_data_from_read[3] (mem_data_from_read[3]), .\data_from_read[3] (\data_from_read[3] ), 
            .instr_fetch_running_N_943(instr_fetch_running_N_943), .\mem_data_from_read[0] (mem_data_from_read[0]), 
            .\data_from_read[0] (\data_from_read[0] ), .\mem_data_from_read[4] (mem_data_from_read[4]), 
            .\data_from_read[4] (\data_from_read[4] ), .\mem_data_from_read[8] (mem_data_from_read[8]), 
            .\data_from_read[8] (\data_from_read[8] ), .\mem_data_from_read[12] (mem_data_from_read[12]), 
            .\data_from_read[12] (\data_from_read[12] ), .\mem_data_from_read[1] (mem_data_from_read[1]), 
            .\data_from_read[1] (\data_from_read[1] ), .\mem_data_from_read[5] (mem_data_from_read[5]), 
            .\data_from_read[5] (\data_from_read[5] ), .n31932(n31932), 
            .n31922(n31922), .n31819(n31819), .\mem_data_from_read[24] (mem_data_from_read[24]), 
            .\mem_data_from_read[28] (mem_data_from_read[28]), .\mem_data_from_read[25] (mem_data_from_read[25]), 
            .\mem_data_from_read[29] (mem_data_from_read[29]), .\peri_data_out[11] (\peri_data_out[11] ), 
            .\mem_data_from_read[26] (mem_data_from_read[26]), .\mem_data_from_read[30] (mem_data_from_read[30]), 
            .\mem_data_from_read[27] (mem_data_from_read[27]), .\mem_data_from_read[31] (mem_data_from_read[31]), 
            .n31910(n31910), .n31942(n31942), .\mem_data_from_read[18] (mem_data_from_read[18]), 
            .\mem_data_from_read[22] (mem_data_from_read[22]), .gpio_out_sel({gpio_out_sel}), 
            .n14(n14), .n14_adj_12(n14_adj_19), .n31961(n31961), .n5171(n5171), 
            .n28686(n28686), .n18680(n18680), .\qspi_data_buf[9] (qspi_data_buf[9]), 
            .\qspi_data_buf[13] (qspi_data_buf[13]), .n27776(n27776), .n27772(n27772), 
            .n27780(n27780), .\qspi_data_buf[11] (qspi_data_buf[11]), .\qspi_data_buf[15] (qspi_data_buf[15]), 
            .\qspi_data_buf[10] (qspi_data_buf[10]), .\qspi_data_buf[14] (qspi_data_buf[14]), 
            .n31899(n31899), .clk_c_enable_273(clk_c_enable_273), .clk_c_enable_357(clk_c_enable_357), 
            .clk_c_enable_349(clk_c_enable_349), .n32003(n32003), .clk_c_enable_259(clk_c_enable_259), 
            .clk_c_enable_360(clk_c_enable_360), .n31904(n31904), .n10573(n10573), 
            .instr_fetch_stopped(instr_fetch_stopped), .n31841(n31841), 
            .n15604(n15604), .n29004(n29004), .n31798(n31798), .clk_c_enable_234(clk_c_enable_234), 
            .\ui_in_sync[0] (\ui_in_sync[0] ), .n1160(n1160), .\alu_b_in[3] (\alu_b_in[3] ), 
            .debug_rd({debug_rd}), .\ui_in_sync[1] (\ui_in_sync[1] ), .\next_fsm_state_3__N_3015[3] (\next_fsm_state_3__N_3015[3] ), 
            .fsm_state({fsm_state_adj_25}), .accum({accum}), .d_3__N_1868({d_3__N_1868}), 
            .n31929(n31929), .\mul_out[1] (\mul_out[1] ), .\mul_out[2] (\mul_out[2] ), 
            .\mul_out[3] (\mul_out[3] ), .n31963(n31963), .next_bit(next_bit), 
            .n28800(n28800), .n31389(n31389), .alu_b_in_3__N_1504(alu_b_in_3__N_1504), 
            .\mem_data_from_read[17] (mem_data_from_read[17]), .\mem_data_from_read[21] (mem_data_from_read[21]), 
            .n29162(n29162), .n18086(n18086), .\csr_read_3__N_1447[2] (\csr_read_3__N_1447[2] ), 
            .GND_net(GND_net), .\next_accum[5] (\next_accum[5] ), .\next_accum[6] (\next_accum[6] ), 
            .\next_accum[7] (\next_accum[7] ), .\next_accum[8] (\next_accum[8] ), 
            .\next_accum[9] (\next_accum[9] ), .\next_accum[10] (\next_accum[10] ), 
            .\next_accum[11] (\next_accum[11] ), .\next_accum[12] (\next_accum[12] ), 
            .\next_accum[13] (\next_accum[13] ), .\next_accum[14] (\next_accum[14] ), 
            .\next_accum[15] (\next_accum[15] ), .\next_accum[16] (\next_accum[16] ), 
            .\next_accum[17] (\next_accum[17] ), .\next_accum[18] (\next_accum[18] ), 
            .\next_accum[19] (\next_accum[19] ), .\next_accum[4] (\next_accum[4] ), 
            .n12(n12), .n11(n11), .n9(n9), .n8_adj_13(n8_adj_23), .\registers[5][7] (\registers[5][7] ), 
            .\registers[6][7] (\registers[6][7] ), .\registers[7][7] (\registers[7][7] ), 
            .n27762(n27762), .n29747(n29747), .n4_adj_14(n4_adj_24)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(94[14] 130[6])
    
endmodule
//
// Verilog Description of module tinyqv_mem_ctrl
//

module tinyqv_mem_ctrl (clk_c, data_txn_len, n26036, qspi_write_done, 
            data_stall, rst_reg_n, n29198, instr_data, \mem_data_from_read[23] , 
            \mem_data_from_read[22] , \mem_data_from_read[21] , \mem_data_from_read[20] , 
            \mem_data_from_read[19] , \mem_data_from_read[18] , \mem_data_from_read[17] , 
            \mem_data_from_read[16] , \qspi_data_buf[15] , \qspi_data_buf[14] , 
            \qspi_data_buf[13] , \qspi_data_buf[11] , \qspi_data_buf[10] , 
            \qspi_data_buf[9] , n31930, clk_c_enable_445, debug_data_continue, 
            instr_active, start_instr, n31940, is_writing, stop_txn_now_N_2363, 
            n31862, n31713, instr_fetch_stopped, n31977, \instr_addr_23__N_318[7] , 
            \addr[8] , \instr_addr_23__N_318[11] , \addr[12] , \addr[24] , 
            instr_active_N_2106, \instr_addr_23__N_318[9] , \addr[10] , 
            \instr_addr_23__N_318[12] , \addr[13] , instr_fetch_running_N_945, 
            n10500, n31730, \instr_addr_23__N_318[13] , \addr[14] , 
            \instr_addr_23__N_318[3] , \addr[4] , \instr_addr_23__N_318[22] , 
            \addr[23] , \instr_addr_23__N_318[10] , \addr[11] , \instr_addr_23__N_318[4] , 
            \addr[5] , mem_data_ready, \mem_data_from_read[31] , \mem_data_from_read[27] , 
            \mem_data_from_read[30] , \mem_data_from_read[26] , \mem_data_from_read[29] , 
            \mem_data_from_read[25] , \mem_data_from_read[28] , \mem_data_from_read[24] , 
            \instr_addr_23__N_318[8] , \addr[9] , \instr_addr_23__N_318[6] , 
            \addr[7] , \instr_addr_23__N_318[5] , \addr[6] , \instr_addr_23__N_318[14] , 
            \addr[15] , \instr_addr_23__N_318[15] , \addr[16] , \instr_addr_23__N_318[16] , 
            \addr[17] , \instr_addr_23__N_318[17] , \addr[18] , \instr_addr_23__N_318[18] , 
            \addr[19] , \instr_addr_23__N_318[19] , \addr[20] , \instr_addr_23__N_318[20] , 
            \addr[21] , \instr_addr_23__N_318[21] , \addr[22] , \instr_addr_23__N_318[2] , 
            \addr[3] , \instr_addr[2] , \addr[2] , \instr_addr[1] , 
            \addr[1] , qspi_data_ready, \txn_len[1] , n31958, debug_stop_txn_N_2147, 
            n58, n18588, n31939, data_stall_N_2158, n31941, continue_txn_N_2131, 
            n10499, n31908, n31887, data_to_write, n32052, n31792, 
            \mem_data_from_read[5] , n31716, n27702, n13146, \mem_data_from_read[1] , 
            \mem_data_from_read[4] , \mem_data_from_read[0] , \mem_data_from_read[3] , 
            \mem_data_from_read[7] , n31725, is_writing_N_2331, n33479, 
            \mem_data_from_read[12] , n27310, \mem_data_from_read[8] , 
            n31741, n8, n27762, instr_fetch_running_N_943, n31907, 
            \addr[0] , n31770, fsm_state, clk_c_enable_231, n31717, 
            clk_c_enable_186, qspi_ram_b_select, clk_c_enable_239, qspi_ram_a_select, 
            n29199, \qspi_data_out_3__N_5[0] , \nibbles_remaining[0] , 
            n32077, clk_c_enable_452, n31906, n6228, n1084, \writing_N_164[3] , 
            n31971, n27464, clk_N_45, \qspi_data_out_3__N_5[2] , n27081, 
            \qspi_data_oe[0] , clk_c_enable_324, stop_txn_reg, n8135, 
            instr_fetch_running, n31942, debug_stop_txn, n31950, \qspi_data_in[0] , 
            \qspi_data_out_3__N_5[3] , \qspi_data_in_3__N_1[0] , \addr[21]_adj_15 , 
            n31736, spi_clk_pos_derived_59, qspi_clk_N_56, n31712, n1176, 
            n27030, n8_adj_16, n3, n6232, n27620, n27183, \qspi_data_in[2] , 
            \qspi_data_in[3] , n32020, n27680, \instr_addr_23__N_318[0] , 
            n31910, n31994, n27776, n31991, n27772, n31990, n27780, 
            n31593) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output [1:0]data_txn_len;
    input n26036;
    output qspi_write_done;
    output data_stall;
    input rst_reg_n;
    input n29198;
    output [15:0]instr_data;
    output \mem_data_from_read[23] ;
    output \mem_data_from_read[22] ;
    output \mem_data_from_read[21] ;
    output \mem_data_from_read[20] ;
    output \mem_data_from_read[19] ;
    output \mem_data_from_read[18] ;
    output \mem_data_from_read[17] ;
    output \mem_data_from_read[16] ;
    output \qspi_data_buf[15] ;
    output \qspi_data_buf[14] ;
    output \qspi_data_buf[13] ;
    output \qspi_data_buf[11] ;
    output \qspi_data_buf[10] ;
    output \qspi_data_buf[9] ;
    input n31930;
    input clk_c_enable_445;
    input debug_data_continue;
    output instr_active;
    input start_instr;
    output n31940;
    output is_writing;
    output stop_txn_now_N_2363;
    input n31862;
    output n31713;
    output instr_fetch_stopped;
    output n31977;
    input \instr_addr_23__N_318[7] ;
    input \addr[8] ;
    input \instr_addr_23__N_318[11] ;
    input \addr[12] ;
    input \addr[24] ;
    input instr_active_N_2106;
    input \instr_addr_23__N_318[9] ;
    input \addr[10] ;
    input \instr_addr_23__N_318[12] ;
    input \addr[13] ;
    output instr_fetch_running_N_945;
    input n10500;
    input n31730;
    input \instr_addr_23__N_318[13] ;
    input \addr[14] ;
    input \instr_addr_23__N_318[3] ;
    input \addr[4] ;
    input \instr_addr_23__N_318[22] ;
    input \addr[23] ;
    input \instr_addr_23__N_318[10] ;
    input \addr[11] ;
    input \instr_addr_23__N_318[4] ;
    input \addr[5] ;
    output mem_data_ready;
    output \mem_data_from_read[31] ;
    output \mem_data_from_read[27] ;
    output \mem_data_from_read[30] ;
    output \mem_data_from_read[26] ;
    output \mem_data_from_read[29] ;
    output \mem_data_from_read[25] ;
    output \mem_data_from_read[28] ;
    output \mem_data_from_read[24] ;
    input \instr_addr_23__N_318[8] ;
    input \addr[9] ;
    input \instr_addr_23__N_318[6] ;
    input \addr[7] ;
    input \instr_addr_23__N_318[5] ;
    input \addr[6] ;
    input \instr_addr_23__N_318[14] ;
    input \addr[15] ;
    input \instr_addr_23__N_318[15] ;
    input \addr[16] ;
    input \instr_addr_23__N_318[16] ;
    input \addr[17] ;
    input \instr_addr_23__N_318[17] ;
    input \addr[18] ;
    input \instr_addr_23__N_318[18] ;
    input \addr[19] ;
    input \instr_addr_23__N_318[19] ;
    input \addr[20] ;
    input \instr_addr_23__N_318[20] ;
    input \addr[21] ;
    input \instr_addr_23__N_318[21] ;
    input \addr[22] ;
    input \instr_addr_23__N_318[2] ;
    input \addr[3] ;
    input \instr_addr[2] ;
    input \addr[2] ;
    input \instr_addr[1] ;
    input \addr[1] ;
    output qspi_data_ready;
    input \txn_len[1] ;
    input n31958;
    input debug_stop_txn_N_2147;
    input n58;
    input n18588;
    input n31939;
    output data_stall_N_2158;
    input n31941;
    output continue_txn_N_2131;
    input n10499;
    input n31908;
    input n31887;
    input [31:0]data_to_write;
    output n32052;
    output n31792;
    output \mem_data_from_read[5] ;
    output n31716;
    output n27702;
    input n13146;
    output \mem_data_from_read[1] ;
    output \mem_data_from_read[4] ;
    output \mem_data_from_read[0] ;
    output \mem_data_from_read[3] ;
    output \mem_data_from_read[7] ;
    input n31725;
    output is_writing_N_2331;
    output n33479;
    output \mem_data_from_read[12] ;
    output n27310;
    output \mem_data_from_read[8] ;
    input n31741;
    input n8;
    input n27762;
    output instr_fetch_running_N_943;
    input n31907;
    input \addr[0] ;
    output n31770;
    output [2:0]fsm_state;
    input clk_c_enable_231;
    input n31717;
    input clk_c_enable_186;
    output qspi_ram_b_select;
    input clk_c_enable_239;
    output qspi_ram_a_select;
    input n29199;
    input \qspi_data_out_3__N_5[0] ;
    output \nibbles_remaining[0] ;
    output n32077;
    input clk_c_enable_452;
    output n31906;
    output n6228;
    output n1084;
    output \writing_N_164[3] ;
    output n31971;
    output n27464;
    input clk_N_45;
    input \qspi_data_out_3__N_5[2] ;
    input n27081;
    output \qspi_data_oe[0] ;
    input clk_c_enable_324;
    output stop_txn_reg;
    input n8135;
    input instr_fetch_running;
    output n31942;
    output debug_stop_txn;
    input n31950;
    input \qspi_data_in[0] ;
    input \qspi_data_out_3__N_5[3] ;
    output \qspi_data_in_3__N_1[0] ;
    output \addr[21]_adj_15 ;
    output n31736;
    output spi_clk_pos_derived_59;
    output qspi_clk_N_56;
    output n31712;
    input n1176;
    output n27030;
    output n8_adj_16;
    output n3;
    output n6232;
    output n27620;
    output n27183;
    input \qspi_data_in[2] ;
    input \qspi_data_in[3] ;
    input n32020;
    output n27680;
    input \instr_addr_23__N_318[0] ;
    output n31910;
    input n31994;
    output n27776;
    input n31991;
    output n27772;
    input n31990;
    output n27780;
    input n31593;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    wire [1:0]qspi_data_byte_idx;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(59[15:33])
    
    wire clk_c_enable_153, qspi_data_byte_idx_1__N_2025, n9, clk_c_enable_110, 
        n11527, data_ready_N_2109, n6085, clk_c_enable_76;
    wire [31:0]instr_data_7__N_1969;
    wire [31:0]qspi_data_buf;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(58[16:29])
    
    wire clk_c_enable_53, clk_c_enable_61, clk_c_enable_69, continue_txn, 
        clk_c_enable_140;
    wire [1:0]n174;
    
    wire n33476, debug_stop_txn_N_2119, spi_clk_pos, clk_c_enable_118, 
        n23983, n8114, n482, clk_c_enable_495, n11586, n23;
    wire [24:0]addr_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(57[17:24])
    
    wire n31723, n27466, last_ram_b_sel, clk_c_enable_367, n32009, 
        n31881, n32010, debug_stop_txn_N_2120, debug_stop_txn_N_2142, 
        spi_ram_b_select_N_2313, n32018, n1;
    wire [1:0]write_qspi_data_byte_idx_1__N_2021;
    
    wire n31857, n32028, data_ready_N_2113, n29082, n29085, n29088, 
        n29091, n29078, n29075, n29072, n31594, n31583, n31577, 
        n30603, n29069, n29081, n29084, n29087, n29090, data_ready_N_2108, 
        data_ready_N_2112, n27644, spi_ram_a_select_N_2309, n28716, 
        n32038, n31721, n31976;
    wire [1:0]read_cycles_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(105[15:32])
    
    wire data_ready_N_2347, n5, n26722, n31739, n31970;
    wire [2:0]n329;
    
    wire n32041, n31731, n31726, n6738;
    wire [23:0]addr_23__N_2188;
    
    FD1P3IX qspi_data_byte_idx__i0 (.D(n9), .SP(clk_c_enable_153), .CD(qspi_data_byte_idx_1__N_2025), 
            .CK(clk_c), .Q(qspi_data_byte_idx[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam qspi_data_byte_idx__i0.GSR = "DISABLED";
    FD1P3AX data_txn_len_i0_i0 (.D(n26036), .SP(clk_c_enable_110), .CK(clk_c), 
            .Q(data_txn_len[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(177[12] 183[8])
    defparam data_txn_len_i0_i0.GSR = "DISABLED";
    FD1S3IX qspi_write_done_185 (.D(data_ready_N_2109), .CK(clk_c), .CD(n11527), 
            .Q(qspi_write_done)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(173[12] 175[8])
    defparam qspi_write_done_185.GSR = "DISABLED";
    FD1P3IX data_stall_188 (.D(n29198), .SP(rst_reg_n), .CD(n6085), .CK(clk_c), 
            .Q(data_stall)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam data_stall_188.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i1 (.D(instr_data_7__N_1969[0]), .SP(clk_c_enable_76), 
            .CK(clk_c), .Q(instr_data[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i1.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i32 (.D(instr_data_7__N_1969[31]), .SP(clk_c_enable_53), 
            .CK(clk_c), .Q(qspi_data_buf[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i32.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i31 (.D(instr_data_7__N_1969[30]), .SP(clk_c_enable_53), 
            .CK(clk_c), .Q(qspi_data_buf[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i31.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i30 (.D(instr_data_7__N_1969[29]), .SP(clk_c_enable_53), 
            .CK(clk_c), .Q(qspi_data_buf[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i30.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i29 (.D(instr_data_7__N_1969[28]), .SP(clk_c_enable_53), 
            .CK(clk_c), .Q(qspi_data_buf[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i29.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i28 (.D(instr_data_7__N_1969[27]), .SP(clk_c_enable_53), 
            .CK(clk_c), .Q(qspi_data_buf[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i28.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i27 (.D(instr_data_7__N_1969[26]), .SP(clk_c_enable_53), 
            .CK(clk_c), .Q(qspi_data_buf[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i27.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i26 (.D(instr_data_7__N_1969[25]), .SP(clk_c_enable_53), 
            .CK(clk_c), .Q(qspi_data_buf[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i26.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i25 (.D(instr_data_7__N_1969[24]), .SP(clk_c_enable_53), 
            .CK(clk_c), .Q(qspi_data_buf[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i25.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i24 (.D(instr_data_7__N_1969[23]), .SP(clk_c_enable_61), 
            .CK(clk_c), .Q(\mem_data_from_read[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i24.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i23 (.D(instr_data_7__N_1969[22]), .SP(clk_c_enable_61), 
            .CK(clk_c), .Q(\mem_data_from_read[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i23.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i22 (.D(instr_data_7__N_1969[21]), .SP(clk_c_enable_61), 
            .CK(clk_c), .Q(\mem_data_from_read[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i22.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i21 (.D(instr_data_7__N_1969[20]), .SP(clk_c_enable_61), 
            .CK(clk_c), .Q(\mem_data_from_read[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i21.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i20 (.D(instr_data_7__N_1969[19]), .SP(clk_c_enable_61), 
            .CK(clk_c), .Q(\mem_data_from_read[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i20.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i19 (.D(instr_data_7__N_1969[18]), .SP(clk_c_enable_61), 
            .CK(clk_c), .Q(\mem_data_from_read[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i19.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i18 (.D(instr_data_7__N_1969[17]), .SP(clk_c_enable_61), 
            .CK(clk_c), .Q(\mem_data_from_read[17] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i18.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i17 (.D(instr_data_7__N_1969[16]), .SP(clk_c_enable_61), 
            .CK(clk_c), .Q(\mem_data_from_read[16] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i17.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i16 (.D(instr_data_7__N_1969[15]), .SP(clk_c_enable_69), 
            .CK(clk_c), .Q(\qspi_data_buf[15] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i16.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i15 (.D(instr_data_7__N_1969[14]), .SP(clk_c_enable_69), 
            .CK(clk_c), .Q(\qspi_data_buf[14] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i15.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i14 (.D(instr_data_7__N_1969[13]), .SP(clk_c_enable_69), 
            .CK(clk_c), .Q(\qspi_data_buf[13] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i14.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i13 (.D(instr_data_7__N_1969[12]), .SP(clk_c_enable_69), 
            .CK(clk_c), .Q(qspi_data_buf[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i13.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i12 (.D(instr_data_7__N_1969[11]), .SP(clk_c_enable_69), 
            .CK(clk_c), .Q(\qspi_data_buf[11] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i12.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i11 (.D(instr_data_7__N_1969[10]), .SP(clk_c_enable_69), 
            .CK(clk_c), .Q(\qspi_data_buf[10] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i11.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i10 (.D(instr_data_7__N_1969[9]), .SP(clk_c_enable_69), 
            .CK(clk_c), .Q(\qspi_data_buf[9] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i10.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i9 (.D(instr_data_7__N_1969[8]), .SP(clk_c_enable_69), 
            .CK(clk_c), .Q(qspi_data_buf[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i9.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i8 (.D(instr_data_7__N_1969[7]), .SP(clk_c_enable_76), 
            .CK(clk_c), .Q(instr_data[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i8.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i7 (.D(instr_data_7__N_1969[6]), .SP(clk_c_enable_76), 
            .CK(clk_c), .Q(instr_data[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i7.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i6 (.D(instr_data_7__N_1969[5]), .SP(clk_c_enable_76), 
            .CK(clk_c), .Q(instr_data[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i6.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i5 (.D(instr_data_7__N_1969[4]), .SP(clk_c_enable_76), 
            .CK(clk_c), .Q(instr_data[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i5.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i4 (.D(instr_data_7__N_1969[3]), .SP(clk_c_enable_76), 
            .CK(clk_c), .Q(instr_data[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i4.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i3 (.D(instr_data_7__N_1969[2]), .SP(clk_c_enable_76), 
            .CK(clk_c), .Q(instr_data[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i3.GSR = "DISABLED";
    FD1P3AX qspi_data_buf_i2 (.D(instr_data_7__N_1969[1]), .SP(clk_c_enable_76), 
            .CK(clk_c), .Q(instr_data[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(162[12] 168[8])
    defparam qspi_data_buf_i2.GSR = "DISABLED";
    FD1P3AX data_txn_len_i0_i1 (.D(n31930), .SP(clk_c_enable_110), .CK(clk_c), 
            .Q(data_txn_len[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(177[12] 183[8])
    defparam data_txn_len_i0_i1.GSR = "DISABLED";
    FD1P3IX continue_txn_187 (.D(debug_data_continue), .SP(clk_c_enable_140), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(continue_txn)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam continue_txn_187.GSR = "DISABLED";
    FD1P3IX qspi_data_byte_idx__i1 (.D(n174[1]), .SP(clk_c_enable_153), 
            .CD(qspi_data_byte_idx_1__N_2025), .CK(clk_c), .Q(qspi_data_byte_idx[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam qspi_data_byte_idx__i1.GSR = "DISABLED";
    LUT4 instr_active_I_0_2_lut_rep_852 (.A(instr_active), .B(start_instr), 
         .Z(n33476)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam instr_active_I_0_2_lut_rep_852.init = 16'heeee;
    LUT4 i1_4_lut (.A(n31940), .B(debug_stop_txn_N_2119), .C(is_writing), 
         .D(spi_clk_pos), .Z(stop_txn_now_N_2363)) /* synthesis lut_function=(A (B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(91[18] 99[12])
    defparam i1_4_lut.init = 16'h8808;
    LUT4 i1_2_lut_rep_508_3_lut_4_lut (.A(n31862), .B(start_instr), .C(clk_c_enable_118), 
         .D(n23983), .Z(n31713)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i1_2_lut_rep_508_3_lut_4_lut.init = 16'hd000;
    FD1S3IX instr_fetch_stopped_182 (.D(debug_stop_txn_N_2119), .CK(clk_c), 
            .CD(n8114), .Q(instr_fetch_stopped)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam instr_fetch_stopped_182.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n31862), .B(start_instr), .C(n482), 
         .D(n31977), .Z(clk_c_enable_495)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf0fd;
    LUT4 i8960_2_lut_3_lut_4_lut (.A(n31862), .B(start_instr), .C(n482), 
         .D(n31977), .Z(n11586)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(127[21:46])
    defparam i8960_2_lut_3_lut_4_lut.init = 16'hf020;
    LUT4 i6_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr_23__N_318[7] ), 
         .D(\addr[8] ), .Z(n23)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i13_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[11] ), .D(\addr[12] ), .Z(addr_in[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_557 (.A(start_instr), .B(n31723), .C(\addr[24] ), 
         .D(n27466), .Z(clk_c_enable_118)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_4_lut_adj_557.init = 16'hffbf;
    LUT4 i1_2_lut (.A(instr_active), .B(last_ram_b_sel), .Z(n27466)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_2_lut.init = 16'heeee;
    FD1P3IX instr_active_180 (.D(start_instr), .SP(clk_c_enable_367), .CD(instr_active_N_2106), 
            .CK(clk_c), .Q(instr_active)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(103[12] 109[8])
    defparam instr_active_180.GSR = "DISABLED";
    LUT4 data_addr_24__I_0_i11_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[9] ), .D(\addr[10] ), .Z(addr_in[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i14_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[12] ), .D(\addr[13] ), .Z(addr_in[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i14_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX instr_fetch_started_181 (.D(n31730), .CK(clk_c), .CD(n10500), 
            .Q(instr_fetch_running_N_945)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam instr_fetch_started_181.GSR = "DISABLED";
    LUT4 data_addr_24__I_0_i15_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[13] ), .D(\addr[14] ), .Z(addr_in[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i5_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[3] ), .D(\addr[4] ), .Z(addr_in[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i24_3_lut_rep_518_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[22] ), .D(\addr[23] ), .Z(n31723)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i24_3_lut_rep_518_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i12_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[10] ), .D(\addr[11] ), .Z(addr_in[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i6_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[4] ), .D(\addr[5] ), .Z(addr_in[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 qspi_data_buf_31__I_0_189_3_lut (.A(qspi_data_buf[31]), .B(instr_data[15]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[31] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_31__I_0_189_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_27__I_0_3_lut (.A(qspi_data_buf[27]), .B(instr_data[11]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[27] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_27__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_30__I_0_3_lut (.A(qspi_data_buf[30]), .B(instr_data[14]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[30] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_30__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_26__I_0_3_lut (.A(qspi_data_buf[26]), .B(instr_data[10]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[26] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_26__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_29__I_0_3_lut (.A(qspi_data_buf[29]), .B(instr_data[13]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[29] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_29__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_25__I_0_3_lut (.A(qspi_data_buf[25]), .B(instr_data[9]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[25] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_25__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_28__I_0_3_lut (.A(qspi_data_buf[28]), .B(instr_data[12]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[28] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_28__I_0_3_lut.init = 16'hcaca;
    LUT4 qspi_data_buf_24__I_0_3_lut (.A(qspi_data_buf[24]), .B(instr_data[8]), 
         .C(mem_data_ready), .Z(\mem_data_from_read[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(208[29] 210[85])
    defparam qspi_data_buf_24__I_0_3_lut.init = 16'hcaca;
    LUT4 data_addr_24__I_0_i10_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[8] ), .D(\addr[9] ), .Z(addr_in[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i8_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[6] ), .D(\addr[7] ), .Z(addr_in[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i7_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[5] ), .D(\addr[6] ), .Z(addr_in[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i16_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[14] ), .D(\addr[15] ), .Z(addr_in[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12736_3_lut_4_lut (.A(instr_active), .B(start_instr), .C(\instr_addr_23__N_318[15] ), 
         .D(\addr[16] ), .Z(addr_in[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i12736_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i18_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[16] ), .D(\addr[17] ), .Z(addr_in[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i19_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[17] ), .D(\addr[18] ), .Z(addr_in[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i20_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[18] ), .D(\addr[19] ), .Z(addr_in[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i21_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[19] ), .D(\addr[20] ), .Z(addr_in[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i22_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[20] ), .D(\addr[21] ), .Z(addr_in[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i23_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[21] ), .D(\addr[22] ), .Z(addr_in[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i4_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr_23__N_318[2] ), .D(\addr[3] ), .Z(addr_in[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i3_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr[2] ), .D(\addr[2] ), .Z(addr_in[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 data_addr_24__I_0_i2_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\instr_addr[1] ), .D(\addr[1] ), .Z(addr_in[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam data_addr_24__I_0_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_804 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n32009)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam i1_2_lut_rep_804.init = 16'h4444;
    LUT4 i1_3_lut_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n31881), .D(qspi_data_ready), .Z(clk_c_enable_61)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h44f0;
    LUT4 i1_2_lut_rep_805 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .Z(n32010)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam i1_2_lut_rep_805.init = 16'h8888;
    LUT4 i1_3_lut_3_lut_4_lut_adj_558 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n31881), .D(qspi_data_ready), .Z(clk_c_enable_53)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam i1_3_lut_3_lut_4_lut_adj_558.init = 16'h88f0;
    PFUMX debug_stop_txn_I_182 (.BLUT(debug_stop_txn_N_2120), .ALUT(debug_stop_txn_N_2142), 
          .C0(instr_active), .Z(debug_stop_txn_N_2119)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=132, LSE_RLINE=164 */ ;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(instr_active), .B(start_instr), 
         .C(\addr[24] ), .D(\addr[23] ), .Z(spi_ram_b_select_N_2313)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'hefff;
    LUT4 i4476_2_lut_rep_813 (.A(qspi_data_byte_idx[1]), .B(qspi_data_byte_idx[0]), 
         .Z(n32018)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(153[39:65])
    defparam i4476_2_lut_rep_813.init = 16'h6666;
    LUT4 i1_4_lut_4_lut (.A(qspi_data_byte_idx[1]), .B(qspi_data_byte_idx[0]), 
         .C(\txn_len[1] ), .D(n1), .Z(n174[1])) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(153[39:65])
    defparam i1_4_lut_4_lut.init = 16'h6642;
    LUT4 i1_3_lut_4_lut (.A(qspi_data_ready), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(start_instr), .D(n31857), .Z(clk_c_enable_153)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[26:60])
    defparam i1_3_lut_4_lut.init = 16'hfeff;
    LUT4 qspi_data_byte_idx_1__I_0_i3_2_lut_rep_823 (.A(qspi_data_byte_idx[0]), 
         .B(qspi_data_byte_idx[1]), .Z(n32028)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[144:171])
    defparam qspi_data_byte_idx_1__I_0_i3_2_lut_rep_823.init = 16'heeee;
    LUT4 data_stall_I_0_213_2_lut_3_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(data_stall), .Z(data_ready_N_2113)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[144:171])
    defparam data_stall_I_0_213_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_3_lut_3_lut_4_lut_adj_559 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n31881), .D(qspi_data_ready), .Z(clk_c_enable_76)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[144:171])
    defparam i1_3_lut_3_lut_4_lut_adj_559.init = 16'h11f0;
    LUT4 i26465_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[28]), .D(\mem_data_from_read[20] ), .Z(n29082)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26465_3_lut_4_lut.init = 16'hf960;
    LUT4 i26468_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[29]), .D(\mem_data_from_read[21] ), .Z(n29085)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26468_3_lut_4_lut.init = 16'hf960;
    LUT4 i26471_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[30]), .D(\mem_data_from_read[22] ), .Z(n29088)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26471_3_lut_4_lut.init = 16'hf960;
    LUT4 i26474_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[31]), .D(\mem_data_from_read[23] ), .Z(n29091)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26474_3_lut_4_lut.init = 16'hf960;
    LUT4 i26461_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[11] ), .D(instr_data[3]), .Z(n29078)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26461_3_lut_4_lut.init = 16'hf960;
    LUT4 i26458_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[10] ), .D(instr_data[2]), .Z(n29075)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26458_3_lut_4_lut.init = 16'hf960;
    LUT4 i26455_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[9] ), .D(instr_data[1]), .Z(n29072)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26455_3_lut_4_lut.init = 16'hf960;
    LUT4 n5570_bdd_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[25]), .D(\mem_data_from_read[17] ), .Z(n31594)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n5570_bdd_3_lut_4_lut.init = 16'hf960;
    LUT4 n18610_bdd_3_lut_28602_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[26]), .D(\mem_data_from_read[18] ), .Z(n31583)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n18610_bdd_3_lut_28602_4_lut.init = 16'hf960;
    LUT4 n18610_bdd_3_lut_28528_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[27]), .D(\mem_data_from_read[19] ), .Z(n31577)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n18610_bdd_3_lut_28528_4_lut.init = 16'hf960;
    LUT4 n18610_bdd_3_lut_28424_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[24]), .D(\mem_data_from_read[16] ), .Z(n30603)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam n18610_bdd_3_lut_28424_4_lut.init = 16'hf960;
    LUT4 i26452_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[8]), .D(instr_data[0]), .Z(n29069)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26452_3_lut_4_lut.init = 16'hf960;
    LUT4 i26464_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(qspi_data_buf[12]), .D(instr_data[4]), .Z(n29081)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26464_3_lut_4_lut.init = 16'hf960;
    LUT4 i26467_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[13] ), .D(instr_data[5]), .Z(n29084)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26467_3_lut_4_lut.init = 16'hf960;
    LUT4 i26470_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[14] ), .D(instr_data[6]), .Z(n29087)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26470_3_lut_4_lut.init = 16'hf960;
    LUT4 i26473_3_lut_4_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(\qspi_data_buf[15] ), .D(instr_data[7]), .Z(n29090)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i26473_3_lut_4_lut.init = 16'hf960;
    LUT4 i15264_4_lut (.A(n31958), .B(debug_stop_txn_N_2147), .C(n58), 
         .D(n18588), .Z(debug_stop_txn_N_2142)) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[26] 86[20])
    defparam i15264_4_lut.init = 16'hcccd;
    LUT4 data_ready_I_0_206_4_lut (.A(instr_active), .B(data_ready_N_2108), 
         .C(n31939), .D(data_ready_N_2112), .Z(mem_data_ready)) /* synthesis lut_function=(!(A+!(B+!(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[25:190])
    defparam data_ready_I_0_206_4_lut.init = 16'h4544;
    LUT4 qspi_data_ready_I_0_202_2_lut (.A(qspi_data_ready), .B(data_ready_N_2109), 
         .Z(data_ready_N_2108)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(207[43:98])
    defparam qspi_data_ready_I_0_202_2_lut.init = 16'h8888;
    LUT4 i27679_4_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(data_txn_len[0]), .D(data_txn_len[1]), .Z(data_ready_N_2109)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[64:98])
    defparam i27679_4_lut.init = 16'h8421;
    LUT4 i27884_4_lut (.A(qspi_data_byte_idx[0]), .B(n27644), .C(start_instr), 
         .D(instr_active), .Z(n9)) /* synthesis lut_function=(!(A+!((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(148[12] 160[8])
    defparam i27884_4_lut.init = 16'h5551;
    LUT4 i1_3_lut (.A(data_txn_len[0]), .B(data_txn_len[1]), .C(qspi_data_byte_idx[1]), 
         .Z(n27644)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C)))) */ ;
    defparam i1_3_lut.init = 16'h4141;
    LUT4 i1_4_lut_adj_560 (.A(start_instr), .B(n31723), .C(\addr[24] ), 
         .D(instr_active), .Z(spi_ram_a_select_N_2309)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(55[21:48])
    defparam i1_4_lut_adj_560.init = 16'hffef;
    LUT4 i3925_2_lut (.A(continue_txn), .B(rst_reg_n), .Z(n6085)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i3925_2_lut.init = 16'h4444;
    LUT4 continue_txn_I_189_4_lut (.A(n28716), .B(data_ready_N_2108), .C(n32018), 
         .D(data_txn_len[1]), .Z(data_stall_N_2158)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(190[21] 191[76])
    defparam continue_txn_I_189_4_lut.init = 16'hecce;
    LUT4 i1_3_lut_adj_561 (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .C(data_txn_len[0]), .Z(n28716)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)))) */ ;
    defparam i1_3_lut_adj_561.init = 16'h4848;
    LUT4 data_ready_N_2113_I_0_4_lut (.A(data_ready_N_2113), .B(n31941), 
         .C(n31939), .D(mem_data_ready), .Z(continue_txn_N_2131)) /* synthesis lut_function=(!((B (C)+!B (C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(194[30:139])
    defparam data_ready_N_2113_I_0_4_lut.init = 16'h0a2a;
    LUT4 i1_2_lut_rep_833 (.A(instr_active), .B(\addr[24] ), .Z(n32038)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_833.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_562 (.A(instr_active), .B(\addr[24] ), 
         .C(n31730), .D(n10499), .Z(addr_in[24])) /* synthesis lut_function=(!(A+!(B ((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_562.init = 16'h4404;
    LUT4 i2_2_lut_4_lut (.A(n31908), .B(n31887), .C(rst_reg_n), .D(start_instr), 
         .Z(qspi_data_byte_idx_1__N_2025)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i2_2_lut_4_lut.init = 16'hff7f;
    LUT4 instr_data_7__I_173_i1_3_lut (.A(data_to_write[0]), .B(instr_data[8]), 
         .C(qspi_data_ready), .Z(instr_data_7__N_1969[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i1_3_lut.init = 16'hcaca;
    LUT4 i8815_3_lut (.A(data_to_write[31]), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8815_3_lut.init = 16'hcaca;
    LUT4 i8817_3_lut (.A(data_to_write[30]), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8817_3_lut.init = 16'hcaca;
    LUT4 i8819_3_lut (.A(data_to_write[29]), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8819_3_lut.init = 16'hcaca;
    LUT4 i8821_3_lut (.A(data_to_write[28]), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8821_3_lut.init = 16'hcaca;
    LUT4 i8823_3_lut (.A(data_to_write[27]), .B(instr_data[11]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8823_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i27_4_lut (.A(data_to_write[26]), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n32010), .Z(instr_data_7__N_1969[26])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i27_4_lut.init = 16'hca0a;
    LUT4 i8825_3_lut (.A(data_to_write[23]), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8825_3_lut.init = 16'hcaca;
    LUT4 i8827_3_lut (.A(data_to_write[22]), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8827_3_lut.init = 16'hcaca;
    LUT4 i8829_3_lut (.A(data_to_write[21]), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8829_3_lut.init = 16'hcaca;
    LUT4 i8831_3_lut (.A(data_to_write[20]), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8831_3_lut.init = 16'hcaca;
    LUT4 i8833_3_lut (.A(data_to_write[19]), .B(instr_data[11]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8833_3_lut.init = 16'hcaca;
    LUT4 i8835_3_lut (.A(data_to_write[15]), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8835_3_lut.init = 16'hcaca;
    LUT4 i8837_3_lut (.A(data_to_write[14]), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8837_3_lut.init = 16'hcaca;
    LUT4 i8839_3_lut (.A(data_to_write[13]), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8839_3_lut.init = 16'hcaca;
    LUT4 i8841_3_lut (.A(data_to_write[12]), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8841_3_lut.init = 16'hcaca;
    LUT4 i8843_3_lut (.A(data_to_write[11]), .B(instr_data[11]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8843_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i11_4_lut (.A(data_to_write[10]), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n32052), .Z(instr_data_7__N_1969[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i11_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i10_4_lut (.A(data_to_write[9]), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n32052), .Z(instr_data_7__N_1969[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i10_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i9_4_lut (.A(data_to_write[8]), .B(instr_data[8]), 
         .C(qspi_data_ready), .D(n32052), .Z(instr_data_7__N_1969[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i9_4_lut.init = 16'h0aca;
    LUT4 i8845_3_lut (.A(data_to_write[7]), .B(instr_data[15]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8845_3_lut.init = 16'hcaca;
    LUT4 i8847_3_lut (.A(data_to_write[6]), .B(instr_data[14]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8847_3_lut.init = 16'hcaca;
    LUT4 i8849_3_lut (.A(data_to_write[5]), .B(instr_data[13]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8849_3_lut.init = 16'hcaca;
    LUT4 i8851_3_lut (.A(data_to_write[4]), .B(instr_data[12]), .C(qspi_data_ready), 
         .Z(instr_data_7__N_1969[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam i8851_3_lut.init = 16'hcaca;
    LUT4 instr_data_7__I_173_i4_4_lut (.A(data_to_write[3]), .B(instr_data[11]), 
         .C(qspi_data_ready), .D(n32028), .Z(instr_data_7__N_1969[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i4_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i3_4_lut (.A(data_to_write[2]), .B(instr_data[10]), 
         .C(qspi_data_ready), .D(n32028), .Z(instr_data_7__N_1969[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i3_4_lut.init = 16'h0aca;
    LUT4 instr_data_7__I_173_i2_4_lut (.A(data_to_write[1]), .B(instr_data[9]), 
         .C(qspi_data_ready), .D(n32028), .Z(instr_data_7__N_1969[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(165[18] 167[12])
    defparam instr_data_7__I_173_i2_4_lut.init = 16'h0aca;
    LUT4 addr_23__I_201_2_lut_rep_516_3_lut_4_lut (.A(n31887), .B(n31908), 
         .C(n31977), .D(start_instr), .Z(n31721)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (C))) */ ;
    defparam addr_23__I_201_2_lut_rep_516_3_lut_4_lut.init = 16'h0f07;
    LUT4 i1_3_lut_4_lut_4_lut (.A(continue_txn), .B(data_ready_N_2109), 
         .C(write_qspi_data_byte_idx_1__N_2021[0]), .D(qspi_data_ready), 
         .Z(debug_stop_txn_N_2120)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(87[102:115])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 qspi_data_byte_idx_1__I_0_197_i3_2_lut_rep_847 (.A(qspi_data_byte_idx[0]), 
         .B(qspi_data_byte_idx[1]), .Z(n32052)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam qspi_data_byte_idx_1__I_0_197_i3_2_lut_rep_847.init = 16'hdddd;
    LUT4 i1_3_lut_3_lut_4_lut_adj_563 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(n31881), .D(qspi_data_ready), .Z(clk_c_enable_69)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam i1_3_lut_3_lut_4_lut_adj_563.init = 16'h22f0;
    LUT4 i1_2_lut_rep_771_3_lut (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(instr_active), .Z(n31976)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam i1_2_lut_rep_771_3_lut.init = 16'h2020;
    LUT4 instr_data_7__I_0_i6_3_lut_4_lut (.A(data_txn_len[0]), .B(n31792), 
         .C(instr_data[13]), .D(instr_data[5]), .Z(\mem_data_from_read[5] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_rep_511_3_lut_4_lut (.A(n31887), .B(n31908), .C(n23983), 
         .D(start_instr), .Z(n31716)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_rep_511_3_lut_4_lut.init = 16'hf070;
    LUT4 i1_2_lut_3_lut_4_lut_adj_564 (.A(qspi_data_byte_idx[0]), .B(qspi_data_byte_idx[1]), 
         .C(qspi_data_ready), .D(instr_active), .Z(n27702)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(81[50:77])
    defparam i1_2_lut_3_lut_4_lut_adj_564.init = 16'h0200;
    LUT4 i27721_2_lut_3_lut (.A(read_cycles_count[1]), .B(data_stall), .C(n13146), 
         .Z(data_ready_N_2347)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i27721_2_lut_3_lut.init = 16'h0101;
    LUT4 i27728_3_lut_4_lut (.A(read_cycles_count[1]), .B(data_stall), .C(n13146), 
         .D(n5), .Z(n26722)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i27728_3_lut_4_lut.init = 16'h0001;
    LUT4 instr_data_7__I_0_i2_3_lut_4_lut (.A(data_txn_len[0]), .B(n31792), 
         .C(instr_data[9]), .D(instr_data[1]), .Z(\mem_data_from_read[1] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i5_3_lut_4_lut (.A(data_txn_len[0]), .B(n31792), 
         .C(instr_data[12]), .D(instr_data[4]), .Z(\mem_data_from_read[4] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i1_3_lut_4_lut (.A(data_txn_len[0]), .B(n31792), 
         .C(instr_data[8]), .D(instr_data[0]), .Z(\mem_data_from_read[0] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i4_3_lut_4_lut (.A(data_txn_len[0]), .B(n31792), 
         .C(instr_data[11]), .D(instr_data[3]), .Z(\mem_data_from_read[3] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 instr_data_7__I_0_i8_3_lut_4_lut (.A(data_txn_len[0]), .B(n31792), 
         .C(instr_data[15]), .D(instr_data[7]), .Z(\mem_data_from_read[7] )) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam instr_data_7__I_0_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_adj_565 (.A(start_instr), .B(n31725), .C(n31908), .D(n32038), 
         .Z(is_writing_N_2331)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_565.init = 16'h1000;
    LUT4 i1_2_lut_rep_534 (.A(data_stall), .B(n13146), .Z(n31739)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i1_2_lut_rep_534.init = 16'heeee;
    LUT4 mux_105_i1_3_lut_4_lut (.A(data_stall), .B(n13146), .C(n33479), 
         .D(n31970), .Z(n329[0])) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam mux_105_i1_3_lut_4_lut.init = 16'hf101;
    LUT4 qspi_data_buf_15__I_0_i5_3_lut_4_lut (.A(data_txn_len[0]), .B(n31792), 
         .C(instr_data[12]), .D(qspi_data_buf[12]), .Z(\mem_data_from_read[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam qspi_data_buf_15__I_0_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_rep_526_3_lut_4_lut (.A(data_stall), .B(n13146), .C(n27310), 
         .D(n32041), .Z(n31731)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(185[12] 205[8])
    defparam i1_rep_526_3_lut_4_lut.init = 16'hfef0;
    LUT4 qspi_data_buf_15__I_0_i1_3_lut_4_lut (.A(data_txn_len[0]), .B(n31792), 
         .C(instr_data[8]), .D(qspi_data_buf[8]), .Z(\mem_data_from_read[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam qspi_data_buf_15__I_0_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_566 (.A(instr_fetch_running_N_945), .B(n31741), .C(n8), 
         .D(n27762), .Z(instr_fetch_running_N_943)) /* synthesis lut_function=(A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(138[12] 146[8])
    defparam i1_4_lut_adj_566.init = 16'ha2aa;
    LUT4 i5568_4_lut (.A(n31862), .B(continue_txn_N_2131), .C(continue_txn), 
         .D(data_stall_N_2158), .Z(clk_c_enable_140)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(198[22] 203[16])
    defparam i5568_4_lut.init = 16'h05c5;
    LUT4 equal_58_i1_4_lut (.A(qspi_data_byte_idx[0]), .B(instr_active), 
         .C(start_instr), .D(data_txn_len[0]), .Z(n1)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(155[21:50])
    defparam equal_58_i1_4_lut.init = 16'h5556;
    LUT4 i1_3_lut_rep_652_4_lut (.A(n31939), .B(n31907), .C(rst_reg_n), 
         .D(n31908), .Z(n31857)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i1_3_lut_rep_652_4_lut.init = 16'he000;
    LUT4 i1_2_lut_rep_521_3_lut_4_lut (.A(n31939), .B(n31907), .C(start_instr), 
         .D(n31908), .Z(n31726)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam i1_2_lut_rep_521_3_lut_4_lut.init = 16'hf1ff;
    LUT4 i27708_2_lut_3_lut_4_lut (.A(n31939), .B(n31907), .C(rst_reg_n), 
         .D(n31908), .Z(clk_c_enable_110)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;
    defparam i27708_2_lut_3_lut_4_lut.init = 16'h1fff;
    LUT4 i4455_2_lut (.A(qspi_data_byte_idx[0]), .B(write_qspi_data_byte_idx_1__N_2021[0]), 
         .Z(n6738)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(111[43:95])
    defparam i4455_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_rep_676_4_lut (.A(n31941), .B(n31940), .C(data_stall), 
         .D(n31939), .Z(n31881)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(91[18] 99[12])
    defparam i1_3_lut_rep_676_4_lut.init = 16'h00f2;
    LUT4 data_ready_I_178_2_lut_3_lut_4_lut (.A(n31941), .B(n31940), .C(data_ready_N_2113), 
         .D(n31939), .Z(data_ready_N_2112)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(91[18] 99[12])
    defparam data_ready_I_178_2_lut_3_lut_4_lut.init = 16'hf0f2;
    LUT4 i1_4_lut_adj_567 (.A(n31725), .B(n31721), .C(instr_active), .D(\addr[0] ), 
         .Z(addr_23__N_2188[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_567.init = 16'h0400;
    LUT4 i1_2_lut_rep_587 (.A(mem_data_ready), .B(data_txn_len[1]), .Z(n31792)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_587.init = 16'h2222;
    LUT4 i1_2_lut_rep_565_3_lut (.A(mem_data_ready), .B(data_txn_len[1]), 
         .C(data_txn_len[0]), .Z(n31770)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_565_3_lut.init = 16'h2020;
    qspi_controller q_ctrl (.n31583(n31583), .fsm_state({fsm_state}), .clk_c(clk_c), 
            .clk_c_enable_231(clk_c_enable_231), .n31717(n31717), .n29075(n29075), 
            .clk_c_enable_186(clk_c_enable_186), .n31577(n31577), .qspi_ram_b_select(qspi_ram_b_select), 
            .clk_c_enable_239(clk_c_enable_239), .spi_ram_b_select_N_2313(spi_ram_b_select_N_2313), 
            .n29078(n29078), .qspi_ram_a_select(qspi_ram_a_select), .spi_ram_a_select_N_2309(spi_ram_a_select_N_2309), 
            .spi_clk_pos(spi_clk_pos), .is_writing(is_writing), .clk_c_enable_118(clk_c_enable_118), 
            .n29199(n29199), .clk_c_enable_445(clk_c_enable_445), .\qspi_data_out_3__N_5[0] (\qspi_data_out_3__N_5[0] ), 
            .\instr_data[12] (instr_data[12]), .nibbles_remaining({Open_71, 
            Open_72, \nibbles_remaining[0] }), .n33479(n33479), .n32077(n32077), 
            .\read_cycles_count[1] (read_cycles_count[1]), .clk_c_enable_452(clk_c_enable_452), 
            .n31906(n31906), .n31977(n31977), .n5(n5), .n6228(n6228), 
            .\addr_in[24] (addr_in[24]), .n1084(n1084), .n26722(n26722), 
            .n31716(n31716), .\writing_N_164[3] (\writing_N_164[3] ), .\instr_data[8] (instr_data[8]), 
            .n31971(n31971), .n31970(n31970), .n27464(n27464), .last_ram_b_sel(last_ram_b_sel), 
            .clk_N_45(clk_N_45), .\qspi_data_out_3__N_5[2] (\qspi_data_out_3__N_5[2] ), 
            .\write_qspi_data_byte_idx_1__N_2021[0] (write_qspi_data_byte_idx_1__N_2021[0]), 
            .n27081(n27081), .\qspi_data_oe[0] (\qspi_data_oe[0] ), .clk_c_enable_324(clk_c_enable_324), 
            .clk_c_enable_495(clk_c_enable_495), .\addr_23__N_2188[0] (addr_23__N_2188[0]), 
            .n32041(n32041), .stop_txn_reg(stop_txn_reg), .qspi_data_ready(qspi_data_ready), 
            .n8135(n8135), .n31713(n31713), .instr_active(instr_active), 
            .n32052(n32052), .instr_fetch_running(instr_fetch_running), 
            .n31942(n31942), .debug_stop_txn(debug_stop_txn), .rst_reg_n(rst_reg_n), 
            .clk_c_enable_367(clk_c_enable_367), .qspi_write_done(qspi_write_done), 
            .n8114(n8114), .debug_stop_txn_N_2119(debug_stop_txn_N_2119), 
            .n13146(n13146), .data_stall(data_stall), .n31726(n31726), 
            .\addr_in[7] (addr_in[7]), .\addr_in[6] (addr_in[6]), .\addr_in[5] (addr_in[5]), 
            .n31950(n31950), .n31731(n31731), .\addr_in[4] (addr_in[4]), 
            .\qspi_data_in[0] (\qspi_data_in[0] ), .start_instr(start_instr), 
            .n31723(n31723), .\addr[24] (\addr[24] ), .n23983(n23983), 
            .\addr_in[18] (addr_in[18]), .n23(n23), .\addr_in[9] (addr_in[9]), 
            .\addr_in[10] (addr_in[10]), .n482(n482), .\addr_in[11] (addr_in[11]), 
            .\addr_in[12] (addr_in[12]), .\addr_in[13] (addr_in[13]), .\addr_in[14] (addr_in[14]), 
            .\addr_in[15] (addr_in[15]), .\addr_in[16] (addr_in[16]), .\qspi_data_out_3__N_5[3] (\qspi_data_out_3__N_5[3] ), 
            .\qspi_data_in_3__N_1[0] (\qspi_data_in_3__N_1[0] ), .\addr[21] (\addr[21]_adj_15 ), 
            .\instr_data[9] (instr_data[9]), .n11586(n11586), .\addr_in[3] (addr_in[3]), 
            .\addr_in[2] (addr_in[2]), .\addr_in[1] (addr_in[1]), .\instr_data[10] (instr_data[10]), 
            .\instr_data[11] (instr_data[11]), .\instr_data[13] (instr_data[13]), 
            .\instr_data[14] (instr_data[14]), .\instr_data[15] (instr_data[15]), 
            .\addr_in[17] (addr_in[17]), .\addr_in[19] (addr_in[19]), .\addr_in[20] (addr_in[20]), 
            .\addr_in[21] (addr_in[21]), .\addr_in[22] (addr_in[22]), .n33476(n33476), 
            .data_ready_N_2347(data_ready_N_2347), .n27310(n27310), .n31739(n31739), 
            .n332(n329[0]), .n11527(n11527), .stop_txn_now_N_2363(stop_txn_now_N_2363), 
            .n31736(n31736), .\data_to_write[25] (data_to_write[25]), .n32010(n32010), 
            .\instr_data_7__N_1969[25] (instr_data_7__N_1969[25]), .\data_to_write[24] (data_to_write[24]), 
            .\instr_data_7__N_1969[24] (instr_data_7__N_1969[24]), .\data_to_write[18] (data_to_write[18]), 
            .n32009(n32009), .\instr_data_7__N_1969[18] (instr_data_7__N_1969[18]), 
            .\data_to_write[17] (data_to_write[17]), .\instr_data_7__N_1969[17] (instr_data_7__N_1969[17]), 
            .\data_to_write[16] (data_to_write[16]), .\instr_data_7__N_1969[16] (instr_data_7__N_1969[16]), 
            .spi_clk_pos_derived_59(spi_clk_pos_derived_59), .qspi_clk_N_56(qspi_clk_N_56), 
            .n30603(n30603), .n31712(n31712), .n1176(n1176), .n29085(n29085), 
            .n29088(n29088), .n31940(n31940), .n29069(n29069), .n29081(n29081), 
            .n29084(n29084), .n29087(n29087), .n29090(n29090), .n27030(n27030), 
            .n8(n8_adj_16), .n3(n3), .n6232(n6232), .\qspi_data_byte_idx[1] (qspi_data_byte_idx[1]), 
            .n6738(n6738), .n29082(n29082), .n29091(n29091), .n27620(n27620), 
            .n27183(n27183), .\qspi_data_in[2] (\qspi_data_in[2] ), .\qspi_data_in[3] (\qspi_data_in[3] ), 
            .n31976(n31976), .n32020(n32020), .n27680(n27680), .\instr_addr_23__N_318[0] (\instr_addr_23__N_318[0] ), 
            .n31910(n31910), .n31994(n31994), .n27776(n27776), .n31991(n31991), 
            .n27772(n27772), .n31990(n31990), .n27780(n27780), .n31594(n31594), 
            .n31593(n31593), .n29072(n29072)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(112[21] 136[6])
    
endmodule
//
// Verilog Description of module qspi_controller
//

module qspi_controller (n31583, fsm_state, clk_c, clk_c_enable_231, 
            n31717, n29075, clk_c_enable_186, n31577, qspi_ram_b_select, 
            clk_c_enable_239, spi_ram_b_select_N_2313, n29078, qspi_ram_a_select, 
            spi_ram_a_select_N_2309, spi_clk_pos, is_writing, clk_c_enable_118, 
            n29199, clk_c_enable_445, \qspi_data_out_3__N_5[0] , \instr_data[12] , 
            nibbles_remaining, n33479, n32077, \read_cycles_count[1] , 
            clk_c_enable_452, n31906, n31977, n5, n6228, \addr_in[24] , 
            n1084, n26722, n31716, \writing_N_164[3] , \instr_data[8] , 
            n31971, n31970, n27464, last_ram_b_sel, clk_N_45, \qspi_data_out_3__N_5[2] , 
            \write_qspi_data_byte_idx_1__N_2021[0] , n27081, \qspi_data_oe[0] , 
            clk_c_enable_324, clk_c_enable_495, \addr_23__N_2188[0] , 
            n32041, stop_txn_reg, qspi_data_ready, n8135, n31713, 
            instr_active, n32052, instr_fetch_running, n31942, debug_stop_txn, 
            rst_reg_n, clk_c_enable_367, qspi_write_done, n8114, debug_stop_txn_N_2119, 
            n13146, data_stall, n31726, \addr_in[7] , \addr_in[6] , 
            \addr_in[5] , n31950, n31731, \addr_in[4] , \qspi_data_in[0] , 
            start_instr, n31723, \addr[24] , n23983, \addr_in[18] , 
            n23, \addr_in[9] , \addr_in[10] , n482, \addr_in[11] , 
            \addr_in[12] , \addr_in[13] , \addr_in[14] , \addr_in[15] , 
            \addr_in[16] , \qspi_data_out_3__N_5[3] , \qspi_data_in_3__N_1[0] , 
            \addr[21] , \instr_data[9] , n11586, \addr_in[3] , \addr_in[2] , 
            \addr_in[1] , \instr_data[10] , \instr_data[11] , \instr_data[13] , 
            \instr_data[14] , \instr_data[15] , \addr_in[17] , \addr_in[19] , 
            \addr_in[20] , \addr_in[21] , \addr_in[22] , n33476, data_ready_N_2347, 
            n27310, n31739, n332, n11527, stop_txn_now_N_2363, n31736, 
            \data_to_write[25] , n32010, \instr_data_7__N_1969[25] , \data_to_write[24] , 
            \instr_data_7__N_1969[24] , \data_to_write[18] , n32009, \instr_data_7__N_1969[18] , 
            \data_to_write[17] , \instr_data_7__N_1969[17] , \data_to_write[16] , 
            \instr_data_7__N_1969[16] , spi_clk_pos_derived_59, qspi_clk_N_56, 
            n30603, n31712, n1176, n29085, n29088, n31940, n29069, 
            n29081, n29084, n29087, n29090, n27030, n8, n3, n6232, 
            \qspi_data_byte_idx[1] , n6738, n29082, n29091, n27620, 
            n27183, \qspi_data_in[2] , \qspi_data_in[3] , n31976, n32020, 
            n27680, \instr_addr_23__N_318[0] , n31910, n31994, n27776, 
            n31991, n27772, n31990, n27780, n31594, n31593, n29072) /* synthesis syn_module_defined=1 */ ;
    input n31583;
    output [2:0]fsm_state;
    input clk_c;
    input clk_c_enable_231;
    input n31717;
    input n29075;
    input clk_c_enable_186;
    input n31577;
    output qspi_ram_b_select;
    input clk_c_enable_239;
    input spi_ram_b_select_N_2313;
    input n29078;
    output qspi_ram_a_select;
    input spi_ram_a_select_N_2309;
    output spi_clk_pos;
    output is_writing;
    input clk_c_enable_118;
    input n29199;
    input clk_c_enable_445;
    input \qspi_data_out_3__N_5[0] ;
    output \instr_data[12] ;
    output [2:0]nibbles_remaining;
    output n33479;
    output n32077;
    output \read_cycles_count[1] ;
    input clk_c_enable_452;
    output n31906;
    output n31977;
    output n5;
    output n6228;
    input \addr_in[24] ;
    output n1084;
    input n26722;
    input n31716;
    output \writing_N_164[3] ;
    output \instr_data[8] ;
    output n31971;
    output n31970;
    output n27464;
    output last_ram_b_sel;
    input clk_N_45;
    input \qspi_data_out_3__N_5[2] ;
    output \write_qspi_data_byte_idx_1__N_2021[0] ;
    input n27081;
    output \qspi_data_oe[0] ;
    input clk_c_enable_324;
    input clk_c_enable_495;
    input \addr_23__N_2188[0] ;
    output n32041;
    output stop_txn_reg;
    output qspi_data_ready;
    input n8135;
    input n31713;
    input instr_active;
    input n32052;
    input instr_fetch_running;
    output n31942;
    output debug_stop_txn;
    input rst_reg_n;
    output clk_c_enable_367;
    input qspi_write_done;
    output n8114;
    input debug_stop_txn_N_2119;
    input n13146;
    input data_stall;
    input n31726;
    input \addr_in[7] ;
    input \addr_in[6] ;
    input \addr_in[5] ;
    input n31950;
    input n31731;
    input \addr_in[4] ;
    input \qspi_data_in[0] ;
    input start_instr;
    input n31723;
    input \addr[24] ;
    output n23983;
    input \addr_in[18] ;
    input n23;
    input \addr_in[9] ;
    input \addr_in[10] ;
    output n482;
    input \addr_in[11] ;
    input \addr_in[12] ;
    input \addr_in[13] ;
    input \addr_in[14] ;
    input \addr_in[15] ;
    input \addr_in[16] ;
    input \qspi_data_out_3__N_5[3] ;
    output \qspi_data_in_3__N_1[0] ;
    output \addr[21] ;
    output \instr_data[9] ;
    input n11586;
    input \addr_in[3] ;
    input \addr_in[2] ;
    input \addr_in[1] ;
    output \instr_data[10] ;
    output \instr_data[11] ;
    output \instr_data[13] ;
    output \instr_data[14] ;
    output \instr_data[15] ;
    input \addr_in[17] ;
    input \addr_in[19] ;
    input \addr_in[20] ;
    input \addr_in[21] ;
    input \addr_in[22] ;
    input n33476;
    input data_ready_N_2347;
    output n27310;
    input n31739;
    input n332;
    output n11527;
    input stop_txn_now_N_2363;
    output n31736;
    input \data_to_write[25] ;
    input n32010;
    output \instr_data_7__N_1969[25] ;
    input \data_to_write[24] ;
    output \instr_data_7__N_1969[24] ;
    input \data_to_write[18] ;
    input n32009;
    output \instr_data_7__N_1969[18] ;
    input \data_to_write[17] ;
    output \instr_data_7__N_1969[17] ;
    input \data_to_write[16] ;
    output \instr_data_7__N_1969[16] ;
    output spi_clk_pos_derived_59;
    output qspi_clk_N_56;
    input n30603;
    output n31712;
    input n1176;
    input n29085;
    input n29088;
    output n31940;
    input n29069;
    input n29081;
    input n29084;
    input n29087;
    input n29090;
    output n27030;
    output n8;
    output n3;
    output n6232;
    input \qspi_data_byte_idx[1] ;
    input n6738;
    input n29082;
    input n29091;
    output n27620;
    output n27183;
    input \qspi_data_in[2] ;
    input \qspi_data_in[3] ;
    input n31976;
    input n32020;
    output n27680;
    input \instr_addr_23__N_318[0] ;
    output n31910;
    input n31994;
    output n27776;
    input n31991;
    output n27772;
    input n31990;
    output n27780;
    input n31594;
    input n31593;
    input n29072;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire clk_N_45 /* synthesis is_inv_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(29[9:18])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    
    wire n31584, n31581, n29534;
    wire [7:0]data_out_7__N_2177;
    
    wire n31582, n31877, n1067, n31580, n32056;
    wire [1:0]read_cycles_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(105[15:32])
    wire [1:0]n396;
    
    wire n31578, n31575, n31576, n31574, clk_c_enable_41, n27269;
    wire [1:0]delay_cycles_cfg;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(87[15:31])
    
    wire n31665, n32036, n28732, n31667, n31704, n32073, n32043, 
        n31928;
    wire [23:0]addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(84[31:35])
    
    wire n1076, n6224, n33481;
    wire [2:0]n356;
    
    wire n1069, n1068;
    wire [3:0]spi_in_buffer;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(91[15:28])
    
    wire clk_c_enable_462, clk_c_enable_513, n31895, last_ram_a_sel, 
        spi_clk_neg, spi_clk_use_neg, n6, n31882, data_req_N_2318, 
        n32069, n31931, stop_txn_reg_N_2360, data_ready_N_2338, n32053, 
        n27588, n10, n26213;
    wire [23:0]addr_23__N_2188;
    
    wire n26688, n32068, n30600, n27488, n32059, n4, n10910, n31996, 
        n1027;
    wire [2:0]nibbles_remaining_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(86[15:32])
    
    wire n18667, n31918, clk_c_enable_517;
    wire [1:0]n181;
    wire [1:0]n381;
    wire [0:0]n5164;
    
    wire n1054, n24640;
    wire [1:0]n127;
    wire [2:0]n312;
    
    wire n29271;
    wire [2:0]n4342;
    
    wire n28648, n18029, n30604, n30601, n31951, n30602, n32058, 
        n32067, n31919;
    wire [55:0]instr_data_15__N_1959;
    wire [7:0]data_out_7__N_2273;
    
    wire n28858, n32057, n31591, n31595, n31592;
    
    L6MUX21 i28532 (.D0(n31584), .D1(n31581), .SD(n29534), .Z(data_out_7__N_2177[2]));
    PFUMX i28530 (.BLUT(n31583), .ALUT(n31582), .C0(n31877), .Z(n31584));
    FD1P3IX fsm_state__i0 (.D(n1067), .SP(clk_c_enable_231), .CD(n31717), 
            .CK(clk_c), .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i0.GSR = "DISABLED";
    PFUMX i28526 (.BLUT(n29075), .ALUT(n31580), .C0(n32056), .Z(n31581));
    FD1P3IX read_cycles_count__i0 (.D(n396[0]), .SP(clk_c_enable_186), .CD(n31717), 
            .CK(clk_c), .Q(read_cycles_count[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam read_cycles_count__i0.GSR = "DISABLED";
    L6MUX21 i28523 (.D0(n31578), .D1(n31575), .SD(n29534), .Z(data_out_7__N_2177[3]));
    PFUMX i28521 (.BLUT(n31577), .ALUT(n31576), .C0(n31877), .Z(n31578));
    FD1P3JX spi_ram_b_select_229 (.D(spi_ram_b_select_N_2313), .SP(clk_c_enable_239), 
            .PD(n31717), .CK(clk_c), .Q(qspi_ram_b_select)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_ram_b_select_229.GSR = "DISABLED";
    PFUMX i28518 (.BLUT(n29078), .ALUT(n31574), .C0(n32056), .Z(n31575));
    FD1P3JX spi_ram_a_select_228 (.D(spi_ram_a_select_N_2309), .SP(clk_c_enable_239), 
            .PD(n31717), .CK(clk_c), .Q(qspi_ram_a_select)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_ram_a_select_228.GSR = "DISABLED";
    FD1P3AX spi_clk_pos_225 (.D(n27269), .SP(clk_c_enable_41), .CK(clk_c), 
            .Q(spi_clk_pos)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_clk_pos_225.GSR = "DISABLED";
    FD1P3IX is_writing_222 (.D(n29199), .SP(clk_c_enable_118), .CD(n31717), 
            .CK(clk_c), .Q(is_writing)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam is_writing_222.GSR = "DISABLED";
    FD1P3AX delay_cycles_cfg_i0_i0 (.D(\qspi_data_out_3__N_5[0] ), .SP(clk_c_enable_445), 
            .CK(clk_c), .Q(delay_cycles_cfg[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(112[12] 117[8])
    defparam delay_cycles_cfg_i0_i0.GSR = "DISABLED";
    LUT4 spi_data_out_3__N_2165_0__bdd_4_lut_4_lut_4_lut (.A(is_writing), 
         .B(fsm_state[2]), .C(\instr_data[12] ), .D(nibbles_remaining[0]), 
         .Z(n31665)) /* synthesis lut_function=(A (B (C))+!A (B+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_data_out_3__N_2165_0__bdd_4_lut_4_lut_4_lut.init = 16'hc4d5;
    LUT4 i1_3_lut_4_lut_4_lut (.A(fsm_state[0]), .B(fsm_state[1]), .C(fsm_state[2]), 
         .D(n32036), .Z(n28732)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(266[13:21])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h00e3;
    LUT4 n31665_bdd_4_lut (.A(n31665), .B(fsm_state[1]), .C(n31667), .D(fsm_state[0]), 
         .Z(n31704)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam n31665_bdd_4_lut.init = 16'h22f0;
    LUT4 fsm_state_2__bdd_4_lut_28621 (.A(fsm_state[2]), .B(fsm_state[1]), 
         .C(delay_cycles_cfg[0]), .D(fsm_state[0]), .Z(n32073)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam fsm_state_2__bdd_4_lut_28621.init = 16'h0020;
    LUT4 fsm_state_2__bdd_4_lut_28975 (.A(fsm_state[2]), .B(fsm_state[1]), 
         .C(n33479), .D(fsm_state[0]), .Z(n32077)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;
    defparam fsm_state_2__bdd_4_lut_28975.init = 16'h0009;
    LUT4 i1_2_lut_rep_723_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(n32043), 
         .D(fsm_state[1]), .Z(n31928)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_723_4_lut.init = 16'hfff7;
    FD1P3IX read_cycles_count__i1 (.D(n396[1]), .SP(clk_c_enable_186), .CD(n31717), 
            .CK(clk_c), .Q(\read_cycles_count[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam read_cycles_count__i1.GSR = "DISABLED";
    LUT4 spi_data_out_3__N_2165_0__bdd_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(addr[20]), .Z(n31667)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam spi_data_out_3__N_2165_0__bdd_3_lut.init = 16'h2020;
    FD1P3IX nibbles_remaining__i0 (.D(n1076), .SP(clk_c_enable_452), .CD(n31717), 
            .CK(clk_c), .Q(nibbles_remaining[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i0.GSR = "DISABLED";
    LUT4 i3195_4_lut (.A(n31906), .B(n6224), .C(n31977), .D(n5), .Z(n6228)) /* synthesis lut_function=(A (B+(C (D)))+!A !((C (D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i3195_4_lut.init = 16'haccc;
    LUT4 fsm_state_2__I_0_239_i5_2_lut_rep_857 (.A(fsm_state[2]), .B(fsm_state[1]), 
         .C(fsm_state[0]), .Z(n33481)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state_2__I_0_239_i5_2_lut_rep_857.init = 16'hfbfb;
    LUT4 mux_711_i1_4_lut (.A(n356[0]), .B(\addr_in[24] ), .C(n1084), 
         .D(n26722), .Z(n1067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam mux_711_i1_4_lut.init = 16'hcfca;
    FD1P3IX fsm_state__i2 (.D(n1069), .SP(clk_c_enable_231), .CD(n31717), 
            .CK(clk_c), .Q(fsm_state[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1P3IX fsm_state__i1 (.D(n1068), .SP(clk_c_enable_231), .CD(n31717), 
            .CK(clk_c), .Q(fsm_state[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam fsm_state__i1.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n31716), .B(clk_c_enable_118), .C(n31977), 
         .D(n31717), .Z(clk_c_enable_41)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i1_3_lut_4_lut.init = 16'hfff8;
    FD1P3AX spi_in_buffer_i0_i0 (.D(\qspi_data_out_3__N_5[0] ), .SP(clk_c_enable_462), 
            .CK(clk_c), .Q(spi_in_buffer[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i0.GSR = "DISABLED";
    FD1P3JX spi_flash_select_227 (.D(\addr_in[24] ), .SP(clk_c_enable_239), 
            .PD(n31717), .CK(clk_c), .Q(\writing_N_164[3] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_flash_select_227.GSR = "DISABLED";
    FD1P3AX data_i1 (.D(data_out_7__N_2177[0]), .SP(clk_c_enable_513), .CK(clk_c), 
            .Q(\instr_data[8] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i1.GSR = "DISABLED";
    LUT4 i837_2_lut_rep_690_3_lut_4_lut (.A(nibbles_remaining[0]), .B(n32036), 
         .C(spi_clk_pos), .D(n31971), .Z(n31895)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i837_2_lut_rep_690_3_lut_4_lut.init = 16'hef0f;
    FD1S3JX last_ram_a_sel_235 (.D(qspi_ram_a_select), .CK(clk_c), .PD(clk_c_enable_445), 
            .Q(last_ram_a_sel)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(272[12] 280[8])
    defparam last_ram_a_sel_235.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_538 (.A(nibbles_remaining[0]), .B(n32036), .C(n31970), 
         .D(n26722), .Z(n27464)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_3_lut_4_lut_adj_538.init = 16'h000e;
    FD1S3JX last_ram_b_sel_236 (.D(qspi_ram_b_select), .CK(clk_c), .PD(clk_c_enable_445), 
            .Q(last_ram_b_sel)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(272[12] 280[8])
    defparam last_ram_b_sel_236.GSR = "DISABLED";
    FD1S3AX spi_clk_neg_237 (.D(spi_clk_pos), .CK(clk_N_45), .Q(spi_clk_neg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(286[12:54])
    defparam spi_clk_neg_237.GSR = "DISABLED";
    FD1P3AX spi_clk_use_neg_220 (.D(\qspi_data_out_3__N_5[2] ), .SP(clk_c_enable_445), 
            .CK(clk_c), .Q(spi_clk_use_neg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(112[12] 117[8])
    defparam spi_clk_use_neg_220.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(nibbles_remaining[0]), .B(n32036), .C(spi_clk_pos), 
         .D(n31971), .Z(n6)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h10f0;
    LUT4 i1_2_lut_rep_677_3_lut_4_lut_3_lut_4_lut (.A(nibbles_remaining[0]), 
         .B(n32036), .C(spi_clk_pos), .D(n31971), .Z(n31882)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_2_lut_rep_677_3_lut_4_lut_3_lut_4_lut.init = 16'h00e0;
    FD1S3IX data_req_230 (.D(data_req_N_2318), .CK(clk_c), .CD(n27081), 
            .Q(\write_qspi_data_byte_idx_1__N_2021[0] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam data_req_230.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_539 (.A(nibbles_remaining[0]), .B(n32036), .C(is_writing), 
         .D(n31971), .Z(data_req_N_2318)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_3_lut_4_lut_adj_539.init = 16'h0010;
    FD1P3IX spi_data_oe__i0 (.D(n1084), .SP(clk_c_enable_324), .CD(n31717), 
            .CK(clk_c), .Q(\qspi_data_oe[0] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam spi_data_oe__i0.GSR = "DISABLED";
    FD1P3AX addr_i0 (.D(\addr_23__N_2188[0] ), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i0.GSR = "DISABLED";
    LUT4 mux_113_i3_4_lut_4_lut (.A(fsm_state[1]), .B(n32041), .C(n33479), 
         .D(n32069), .Z(n356[2])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam mux_113_i3_4_lut_4_lut.init = 16'h8f8c;
    LUT4 i3456_2_lut_rep_726_3_lut_4_lut (.A(fsm_state[1]), .B(n32041), 
         .C(n32036), .D(nibbles_remaining[0]), .Z(n31931)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i3456_2_lut_rep_726_3_lut_4_lut.init = 16'h4440;
    FD1S3IX stop_txn_reg_218 (.D(stop_txn_reg_N_2360), .CK(clk_c), .CD(clk_c_enable_445), 
            .Q(stop_txn_reg)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(98[12] 103[8])
    defparam stop_txn_reg_218.GSR = "DISABLED";
    FD1S3IX data_ready_224 (.D(data_ready_N_2338), .CK(clk_c), .CD(n8135), 
            .Q(qspi_data_ready)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam data_ready_224.GSR = "DISABLED";
    LUT4 i15783_3_lut_4_lut (.A(n31713), .B(n31977), .C(n26722), .D(n356[2]), 
         .Z(n1069)) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i15783_3_lut_4_lut.init = 16'hddd0;
    LUT4 i1_3_lut_rep_737_4_lut (.A(instr_active), .B(n32052), .C(instr_fetch_running), 
         .D(qspi_data_ready), .Z(n31942)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_3_lut_rep_737_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_adj_540 (.A(fsm_state[0]), .B(n32053), .C(stop_txn_reg), 
         .D(spi_clk_pos), .Z(n27588)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_3_lut_4_lut_adj_540.init = 16'hfff1;
    LUT4 i1_3_lut_4_lut_adj_541 (.A(fsm_state[0]), .B(n32053), .C(debug_stop_txn), 
         .D(rst_reg_n), .Z(clk_c_enable_367)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_3_lut_4_lut_adj_541.init = 16'hf1ff;
    LUT4 i27662_2_lut_3_lut_4_lut (.A(fsm_state[0]), .B(n32053), .C(rst_reg_n), 
         .D(qspi_write_done), .Z(n8114)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i27662_2_lut_3_lut_4_lut.init = 16'h0f1f;
    LUT4 i15265_2_lut_3_lut_4_lut (.A(fsm_state[0]), .B(n32053), .C(debug_stop_txn_N_2119), 
         .D(qspi_write_done), .Z(debug_stop_txn)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i15265_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_4_lut (.A(n10), .B(n13146), .C(is_writing), .D(data_stall), 
         .Z(data_ready_N_2338)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0002;
    LUT4 i21_4_lut (.A(n32041), .B(\read_cycles_count[1] ), .C(n5), .D(n26213), 
         .Z(n10)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A !(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(165[26] 212[20])
    defparam i21_4_lut.init = 16'ha303;
    LUT4 addr_23__I_0_i8_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[7] ), 
         .D(addr[3]), .Z(addr_23__N_2188[7])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i7_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[6] ), 
         .D(addr[2]), .Z(addr_23__N_2188[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i6_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[5] ), 
         .D(addr[1]), .Z(addr_23__N_2188[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i6_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX delay_cycles_cfg_i0_i1 (.D(n31950), .SP(clk_c_enable_445), .CK(clk_c), 
            .Q(delay_cycles_cfg[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(112[12] 117[8])
    defparam delay_cycles_cfg_i0_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_542 (.A(n31906), .B(n31731), .C(n5), .D(n33479), 
         .Z(n26688)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut_adj_542.init = 16'hff7f;
    LUT4 addr_23__I_0_i5_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[4] ), 
         .D(addr[0]), .Z(addr_23__N_2188[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_95_i3_4_lut_4_lut_then_3_lut (.A(fsm_state[0]), .B(fsm_state[1]), 
         .C(fsm_state[2]), .Z(n32068)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;
    defparam mux_95_i3_4_lut_4_lut_then_3_lut.init = 16'h7c7c;
    LUT4 n9_bdd_4_lut_28423 (.A(n31928), .B(\qspi_data_in[0] ), .C(spi_in_buffer[0]), 
         .D(rst_reg_n), .Z(n30600)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam n9_bdd_4_lut_28423.init = 16'he4a0;
    LUT4 i1_4_lut_adj_543 (.A(start_instr), .B(n31723), .C(\addr[24] ), 
         .D(n27488), .Z(n23983)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(109[49:72])
    defparam i1_4_lut_adj_543.init = 16'hffef;
    LUT4 i1_2_lut (.A(instr_active), .B(last_ram_a_sel), .Z(n27488)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(109[49:72])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 addr_23__I_0_i19_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[18] ), 
         .D(addr[14]), .Z(addr_23__N_2188[18])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_718_i3_4_lut (.A(n32059), .B(\addr_in[24] ), .C(n1084), .D(n4), 
         .Z(n10910)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam mux_718_i3_4_lut.init = 16'h3a35;
    LUT4 i1_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(fsm_state[0]), 
         .Z(n5)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(266[13:21])
    defparam i1_3_lut.init = 16'hf7f7;
    LUT4 i1_4_lut_adj_544 (.A(n23983), .B(clk_c_enable_118), .C(n31726), 
         .D(n31977), .Z(n1084)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i1_4_lut_adj_544.init = 16'h0080;
    LUT4 i10_3_lut_4_lut (.A(n31977), .B(n31726), .C(n23), .D(addr[4]), 
         .Z(addr_23__N_2188[8])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 i3197_3_lut_4_lut_3_lut_4_lut (.A(\writing_N_164[3] ), .B(is_writing), 
         .C(n31996), .D(fsm_state[0]), .Z(n1027)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(187[46] 194[40])
    defparam i3197_3_lut_4_lut_3_lut_4_lut.init = 16'h0f02;
    LUT4 addr_23__I_0_i10_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[9] ), 
         .D(addr[5]), .Z(addr_23__N_2188[9])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i11_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[10] ), 
         .D(addr[6]), .Z(addr_23__N_2188[10])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i11_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX nibbles_remaining__i1 (.D(n18667), .SP(clk_c_enable_452), .CD(n31717), 
            .CK(clk_c), .Q(nibbles_remaining_c[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i1.GSR = "DISABLED";
    LUT4 i806_2_lut_rep_713_3_lut_4_lut (.A(\writing_N_164[3] ), .B(is_writing), 
         .C(n31996), .D(fsm_state[0]), .Z(n31918)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(187[46] 194[40])
    defparam i806_2_lut_rep_713_3_lut_4_lut.init = 16'hfff1;
    LUT4 i1_2_lut_rep_791 (.A(fsm_state[2]), .B(fsm_state[1]), .Z(n31996)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_rep_791.init = 16'hbbbb;
    LUT4 i171_2_lut_3_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(spi_clk_pos), 
         .D(fsm_state[0]), .Z(n482)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i171_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 addr_23__I_0_i12_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[11] ), 
         .D(addr[7]), .Z(addr_23__N_2188[11])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i12_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i13_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[12] ), 
         .D(addr[8]), .Z(addr_23__N_2188[12])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i14_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[13] ), 
         .D(addr[9]), .Z(addr_23__N_2188[13])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i15_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[14] ), 
         .D(addr[10]), .Z(addr_23__N_2188[14])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i16_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[15] ), 
         .D(addr[11]), .Z(addr_23__N_2188[15])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i16_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX nibbles_remaining__i2 (.D(n10910), .SP(clk_c_enable_452), .CD(n31717), 
            .CK(clk_c), .Q(nibbles_remaining_c[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam nibbles_remaining__i2.GSR = "DISABLED";
    LUT4 addr_23__I_0_i17_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[16] ), 
         .D(addr[12]), .Z(addr_23__N_2188[16])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i17_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX spi_in_buffer_i0_i1 (.D(n31950), .SP(clk_c_enable_462), .CK(clk_c), 
            .Q(spi_in_buffer[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i1.GSR = "DISABLED";
    FD1P3AX spi_in_buffer_i0_i2 (.D(\qspi_data_out_3__N_5[2] ), .SP(clk_c_enable_462), 
            .CK(clk_c), .Q(spi_in_buffer[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i2.GSR = "DISABLED";
    FD1P3AX spi_in_buffer_i0_i3 (.D(\qspi_data_out_3__N_5[3] ), .SP(clk_c_enable_462), 
            .CK(clk_c), .Q(spi_in_buffer[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam spi_in_buffer_i0_i3.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_545 (.A(\qspi_data_oe[0] ), .B(n31704), .Z(\qspi_data_in_3__N_1[0] )) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_545.init = 16'h8888;
    FD1P3AX addr_i4 (.D(addr_23__N_2188[4]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i4.GSR = "DISABLED";
    FD1P3AX addr_i5 (.D(addr_23__N_2188[5]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i5.GSR = "DISABLED";
    FD1P3AX addr_i6 (.D(addr_23__N_2188[6]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i6.GSR = "DISABLED";
    FD1P3AX addr_i7 (.D(addr_23__N_2188[7]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i7.GSR = "DISABLED";
    FD1P3AX addr_i8 (.D(addr_23__N_2188[8]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i8.GSR = "DISABLED";
    FD1P3AX addr_i9 (.D(addr_23__N_2188[9]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i9.GSR = "DISABLED";
    FD1P3AX addr_i10 (.D(addr_23__N_2188[10]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i10.GSR = "DISABLED";
    FD1P3AX addr_i11 (.D(addr_23__N_2188[11]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i11.GSR = "DISABLED";
    FD1P3AX addr_i12 (.D(addr_23__N_2188[12]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i12.GSR = "DISABLED";
    FD1P3AX addr_i13 (.D(addr_23__N_2188[13]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i13.GSR = "DISABLED";
    FD1P3AX addr_i14 (.D(addr_23__N_2188[14]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i14.GSR = "DISABLED";
    FD1P3AX addr_i15 (.D(addr_23__N_2188[15]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i15.GSR = "DISABLED";
    FD1P3AX addr_i16 (.D(addr_23__N_2188[16]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i16.GSR = "DISABLED";
    FD1P3AX addr_i17 (.D(addr_23__N_2188[17]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i17.GSR = "DISABLED";
    FD1P3AX addr_i18 (.D(addr_23__N_2188[18]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i18.GSR = "DISABLED";
    FD1P3AX addr_i19 (.D(addr_23__N_2188[19]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i19.GSR = "DISABLED";
    FD1P3AX addr_i20 (.D(addr_23__N_2188[20]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i20.GSR = "DISABLED";
    FD1P3AX addr_i21 (.D(addr_23__N_2188[21]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(\addr[21] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i21.GSR = "DISABLED";
    FD1P3AX addr_i22 (.D(addr_23__N_2188[22]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i22.GSR = "DISABLED";
    FD1P3AX addr_i23 (.D(addr_23__N_2188[23]), .SP(clk_c_enable_495), .CK(clk_c), 
            .Q(addr[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i23.GSR = "DISABLED";
    FD1P3AX data_i2 (.D(data_out_7__N_2177[1]), .SP(clk_c_enable_513), .CK(clk_c), 
            .Q(\instr_data[9] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i2.GSR = "DISABLED";
    FD1P3IX addr_i3 (.D(\addr_in[3] ), .SP(clk_c_enable_495), .CD(n11586), 
            .CK(clk_c), .Q(addr[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i3.GSR = "DISABLED";
    FD1P3IX addr_i2 (.D(\addr_in[2] ), .SP(clk_c_enable_495), .CD(n11586), 
            .CK(clk_c), .Q(addr[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i2.GSR = "DISABLED";
    FD1P3IX addr_i1 (.D(\addr_in[1] ), .SP(clk_c_enable_495), .CD(n11586), 
            .CK(clk_c), .Q(addr[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(219[12] 225[8])
    defparam addr_i1.GSR = "DISABLED";
    FD1P3AX data_i3 (.D(data_out_7__N_2177[2]), .SP(clk_c_enable_513), .CK(clk_c), 
            .Q(\instr_data[10] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i3.GSR = "DISABLED";
    FD1P3AX data_i4 (.D(data_out_7__N_2177[3]), .SP(clk_c_enable_513), .CK(clk_c), 
            .Q(\instr_data[11] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i4.GSR = "DISABLED";
    FD1P3AX data_i5 (.D(data_out_7__N_2177[4]), .SP(clk_c_enable_517), .CK(clk_c), 
            .Q(\instr_data[12] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i5.GSR = "DISABLED";
    FD1P3AX data_i6 (.D(data_out_7__N_2177[5]), .SP(clk_c_enable_517), .CK(clk_c), 
            .Q(\instr_data[13] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i6.GSR = "DISABLED";
    FD1P3AX data_i7 (.D(data_out_7__N_2177[6]), .SP(clk_c_enable_517), .CK(clk_c), 
            .Q(\instr_data[14] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i7.GSR = "DISABLED";
    FD1P3AX data_i8 (.D(data_out_7__N_2177[7]), .SP(clk_c_enable_517), .CK(clk_c), 
            .Q(\instr_data[15] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(227[12] 245[8])
    defparam data_i8.GSR = "DISABLED";
    PFUMX mux_129_i1 (.BLUT(n181[0]), .ALUT(n381[0]), .C0(n5), .Z(n396[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 addr_23__I_0_i18_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[17] ), 
         .D(addr[13]), .Z(addr_23__N_2188[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i18_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i20_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[19] ), 
         .D(addr[15]), .Z(addr_23__N_2188[19])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i20_3_lut_4_lut.init = 16'hfb40;
    PFUMX mux_699_i2 (.BLUT(n356[1]), .ALUT(n5164[0]), .C0(n26722), .Z(n1054));
    LUT4 addr_23__I_0_i21_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[20] ), 
         .D(addr[16]), .Z(addr_23__N_2188[20])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i21_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i22_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[21] ), 
         .D(addr[17]), .Z(addr_23__N_2188[21])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i22_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i23_3_lut_4_lut (.A(n31977), .B(n31726), .C(\addr_in[22] ), 
         .D(addr[18]), .Z(addr_23__N_2188[22])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i23_3_lut_4_lut.init = 16'hfb40;
    LUT4 addr_23__I_0_i24_3_lut_4_lut (.A(n31977), .B(n31726), .C(n31723), 
         .D(addr[19]), .Z(addr_23__N_2188[23])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(220[13:65])
    defparam addr_23__I_0_i24_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_711_i2_3_lut_4_lut (.A(n33476), .B(\addr[24] ), .C(n1084), 
         .D(n1054), .Z(n1068)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_711_i2_3_lut_4_lut.init = 16'hbfb0;
    PFUMX i16095 (.BLUT(n24640), .ALUT(n127[1]), .C0(n26688), .Z(n396[1]));
    LUT4 i3196_3_lut_4_lut (.A(n31716), .B(clk_c_enable_118), .C(n31977), 
         .D(data_ready_N_2347), .Z(n6224)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i3196_3_lut_4_lut.init = 16'hf808;
    LUT4 i16038_2_lut (.A(read_cycles_count[0]), .B(\read_cycles_count[1] ), 
         .Z(n127[1])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(151[22:69])
    defparam i16038_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_546 (.A(delay_cycles_cfg[1]), .B(n27310), .C(n31739), 
         .D(n32041), .Z(n24640)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(264[13:21])
    defparam i1_4_lut_adj_546.init = 16'ha088;
    PFUMX mux_113_i1 (.BLUT(n312[0]), .ALUT(n332), .C0(n29271), .Z(n356[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 equal_120_i4_2_lut_rep_831 (.A(nibbles_remaining_c[1]), .B(nibbles_remaining_c[2]), 
         .Z(n32036)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam equal_120_i4_2_lut_rep_831.init = 16'heeee;
    LUT4 i27941_2_lut_3_lut_4_lut (.A(nibbles_remaining_c[1]), .B(nibbles_remaining_c[2]), 
         .C(n32041), .D(nibbles_remaining[0]), .Z(n29271)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i27941_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i4496_2_lut_3_lut_4_lut (.A(nibbles_remaining_c[1]), .B(nibbles_remaining_c[2]), 
         .C(n4342[1]), .D(nibbles_remaining[0]), .Z(n4)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i4496_2_lut_3_lut_4_lut.init = 16'hfff1;
    LUT4 i8901_1_lut (.A(\write_qspi_data_byte_idx_1__N_2021[0] ), .Z(n11527)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i8901_1_lut.init = 16'h5555;
    LUT4 i27676_4_lut (.A(n5), .B(stop_txn_now_N_2363), .C(n27588), .D(rst_reg_n), 
         .Z(n27269)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i27676_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_836 (.A(fsm_state[2]), .B(fsm_state[0]), .Z(n32041)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_836.init = 16'h8888;
    LUT4 i1_3_lut_3_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(fsm_state[1]), 
         .Z(n28648)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)+!B !(C)))) */ ;
    defparam i1_3_lut_3_lut.init = 16'h3434;
    LUT4 i15962_2_lut_rep_765_3_lut (.A(fsm_state[2]), .B(fsm_state[0]), 
         .C(fsm_state[1]), .Z(n31970)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15962_2_lut_rep_765_3_lut.init = 16'h8080;
    LUT4 i15462_3_lut_4_lut_3_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), 
         .C(is_writing), .D(fsm_state[1]), .Z(n18029)) /* synthesis lut_function=(!(A (B ((D)+!C)))) */ ;
    defparam i15462_3_lut_4_lut_3_lut_4_lut.init = 16'h77f7;
    LUT4 i1_2_lut_rep_766_3_lut (.A(fsm_state[2]), .B(fsm_state[0]), .C(fsm_state[1]), 
         .Z(n31971)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_766_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_rep_531_3_lut_4_lut (.A(fsm_state[2]), .B(fsm_state[0]), 
         .C(n13146), .D(data_stall), .Z(n31736)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_2_lut_rep_531_3_lut_4_lut.init = 16'h8880;
    LUT4 i19311_4_lut (.A(\data_to_write[25] ), .B(\instr_data[9] ), .C(qspi_data_ready), 
         .D(n32010), .Z(\instr_data_7__N_1969[25] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i19311_4_lut.init = 16'hca0a;
    LUT4 i11630_4_lut (.A(\data_to_write[24] ), .B(\instr_data[8] ), .C(qspi_data_ready), 
         .D(n32010), .Z(\instr_data_7__N_1969[24] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i11630_4_lut.init = 16'hca0a;
    LUT4 i19314_4_lut (.A(\data_to_write[18] ), .B(\instr_data[10] ), .C(qspi_data_ready), 
         .D(n32009), .Z(\instr_data_7__N_1969[18] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i19314_4_lut.init = 16'hca0a;
    L6MUX21 i27979 (.D0(n30604), .D1(n30601), .SD(n29534), .Z(data_out_7__N_2177[0]));
    LUT4 i19320_4_lut (.A(\data_to_write[17] ), .B(\instr_data[9] ), .C(qspi_data_ready), 
         .D(n32009), .Z(\instr_data_7__N_1969[17] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i19320_4_lut.init = 16'hca0a;
    LUT4 i19318_4_lut (.A(\data_to_write[16] ), .B(\instr_data[8] ), .C(qspi_data_ready), 
         .D(n32009), .Z(\instr_data_7__N_1969[16] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i19318_4_lut.init = 16'hca0a;
    LUT4 i15216_2_lut_rep_838 (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .Z(n32043)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15216_2_lut_rep_838.init = 16'heeee;
    LUT4 i1_3_lut_rep_746_4_lut (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .C(fsm_state[0]), .D(fsm_state[2]), .Z(n31951)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_3_lut_rep_746_4_lut.init = 16'hefff;
    LUT4 i27_3_lut_4_lut (.A(\read_cycles_count[1] ), .B(read_cycles_count[0]), 
         .C(n18029), .D(spi_clk_pos), .Z(n31906)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam i27_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_95_i1_3_lut_4_lut_4_lut_4_lut (.A(fsm_state[0]), .B(n33481), 
         .C(is_writing), .D(\writing_N_164[3] ), .Z(n312[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(266[13:21])
    defparam mux_95_i1_3_lut_4_lut_4_lut_4_lut.init = 16'h7475;
    LUT4 equal_120_i5_2_lut_rep_855 (.A(nibbles_remaining_c[1]), .B(nibbles_remaining_c[2]), 
         .C(nibbles_remaining[0]), .Z(n33479)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam equal_120_i5_2_lut_rep_855.init = 16'hfefe;
    LUT4 spi_clk_pos_I_0_256_3_lut_rep_842 (.A(spi_clk_pos), .B(spi_clk_neg), 
         .C(spi_clk_use_neg), .Z(spi_clk_pos_derived_59)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(287[26:69])
    defparam spi_clk_pos_I_0_256_3_lut_rep_842.init = 16'hcaca;
    LUT4 qspi_clk_I_0_1_lut_3_lut (.A(spi_clk_pos), .B(spi_clk_neg), .C(spi_clk_use_neg), 
         .Z(qspi_clk_N_56)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(287[26:69])
    defparam qspi_clk_I_0_1_lut_3_lut.init = 16'h3535;
    PFUMX i27977 (.BLUT(n30603), .ALUT(n30602), .C0(n31877), .Z(n30604));
    LUT4 i6412_rep_507_3_lut_4_lut (.A(n23983), .B(n31726), .C(n31977), 
         .D(clk_c_enable_118), .Z(n31712)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(139[21:80])
    defparam i6412_rep_507_3_lut_4_lut.init = 16'h0800;
    LUT4 mux_2877_i3_4_lut_then_2_lut_1_lut (.A(nibbles_remaining_c[2]), .Z(n32058)) /* synthesis lut_function=(A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam mux_2877_i3_4_lut_then_2_lut_1_lut.init = 16'haaaa;
    LUT4 mux_95_i3_4_lut_4_lut_else_3_lut (.A(fsm_state[0]), .B(fsm_state[1]), 
         .C(fsm_state[2]), .D(is_writing), .Z(n32067)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;
    defparam mux_95_i3_4_lut_4_lut_else_3_lut.init = 16'h7c78;
    LUT4 mux_114_i1_4_lut_4_lut (.A(read_cycles_count[0]), .B(n31736), .C(n1176), 
         .D(n32073), .Z(n381[0])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam mux_114_i1_4_lut_4_lut.init = 16'h5f5c;
    LUT4 i1_2_lut_rep_848 (.A(fsm_state[1]), .B(fsm_state[2]), .Z(n32053)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_848.init = 16'heeee;
    LUT4 i1_2_lut_rep_714_3_lut_3_lut_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(fsm_state[0]), .Z(n31919)) /* synthesis lut_function=(!(A (B (C))+!A (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_714_3_lut_3_lut_3_lut.init = 16'h2f2f;
    LUT4 i27381_3_lut_4_lut (.A(\instr_data[9] ), .B(n31882), .C(n31877), 
         .D(n29085), .Z(instr_data_15__N_1959[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(231[22] 237[16])
    defparam i27381_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_rep_772_3_lut (.A(fsm_state[1]), .B(fsm_state[2]), .C(fsm_state[0]), 
         .Z(n31977)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam i1_2_lut_rep_772_3_lut.init = 16'hfefe;
    LUT4 i27383_3_lut_4_lut (.A(\instr_data[10] ), .B(n31882), .C(n31877), 
         .D(n29088), .Z(instr_data_15__N_1959[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(231[22] 237[16])
    defparam i27383_3_lut_4_lut.init = 16'h8f80;
    LUT4 qspi_busy_I_0_2_lut_rep_735_3_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[2]), 
         .C(qspi_write_done), .D(fsm_state[0]), .Z(n31940)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(138[17:38])
    defparam qspi_busy_I_0_2_lut_rep_735_3_lut_4_lut.init = 16'hfffe;
    PFUMX i27974 (.BLUT(n29069), .ALUT(n30600), .C0(n32056), .Z(n30601));
    LUT4 i1_3_lut_4_lut_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(fsm_state[0]), 
         .Z(n27310)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(83[15:25])
    defparam i1_3_lut_4_lut_3_lut.init = 16'h0202;
    LUT4 i10573_1_lut_rep_851 (.A(is_writing), .Z(n32056)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i10573_1_lut_rep_851.init = 16'h5555;
    LUT4 mux_60_i1_4_lut_4_lut_4_lut (.A(is_writing), .B(data_ready_N_2347), 
         .C(delay_cycles_cfg[0]), .D(read_cycles_count[0]), .Z(n181[0])) /* synthesis lut_function=(!(A (B+(D))+!A !(B (C)+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_60_i1_4_lut_4_lut_4_lut.init = 16'h4073;
    LUT4 mux_180_i5_3_lut_3_lut (.A(is_writing), .B(\instr_data[8] ), .C(n29081), 
         .Z(data_out_7__N_2273[4])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i5_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i6_3_lut_3_lut (.A(is_writing), .B(\instr_data[9] ), .C(n29084), 
         .Z(data_out_7__N_2273[5])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i6_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i7_3_lut_3_lut (.A(is_writing), .B(\instr_data[10] ), .C(n29087), 
         .Z(data_out_7__N_2273[6])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i7_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_180_i8_3_lut_3_lut (.A(is_writing), .B(\instr_data[11] ), .C(n29090), 
         .Z(data_out_7__N_2273[7])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam mux_180_i8_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_2_lut (.A(is_writing), .B(delay_cycles_cfg[1]), .Z(n5164[0])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i2_3_lut_4_lut_4_lut (.A(is_writing), .B(\instr_data[14] ), .C(fsm_state[1]), 
         .D(fsm_state[2]), .Z(n27030)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0d00;
    LUT4 i1_2_lut_3_lut (.A(fsm_state[2]), .B(fsm_state[1]), .C(addr[22]), 
         .Z(n8)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_547 (.A(fsm_state[2]), .B(fsm_state[1]), .C(addr[23]), 
         .Z(n3)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_3_lut_adj_547.init = 16'h0404;
    LUT4 i3194_4_lut (.A(n31906), .B(n31713), .C(n31977), .D(n5), .Z(n6232)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i3194_4_lut.init = 16'hac0c;
    LUT4 i15454_4_lut (.A(nibbles_remaining[0]), .B(n1084), .C(n28732), 
         .D(n31919), .Z(n1076)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(149[22] 213[16])
    defparam i15454_4_lut.init = 16'hcddd;
    PFUMX data_out_7__I_0_242_i8 (.BLUT(instr_data_15__N_1959[31]), .ALUT(data_out_7__N_2273[7]), 
          .C0(n29534), .Z(data_out_7__N_2177[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i7 (.BLUT(instr_data_15__N_1959[30]), .ALUT(data_out_7__N_2273[6]), 
          .C0(n29534), .Z(data_out_7__N_2177[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i6 (.BLUT(instr_data_15__N_1959[29]), .ALUT(data_out_7__N_2273[5]), 
          .C0(n29534), .Z(data_out_7__N_2177[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    PFUMX data_out_7__I_0_242_i5 (.BLUT(instr_data_15__N_1959[28]), .ALUT(data_out_7__N_2273[4]), 
          .C0(n29534), .Z(data_out_7__N_2177[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=21, LSE_RCOL=6, LSE_LLINE=112, LSE_RLINE=136 */ ;
    LUT4 i1_4_lut_adj_548 (.A(read_cycles_count[0]), .B(is_writing), .C(fsm_state[0]), 
         .D(n28858), .Z(clk_c_enable_462)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_548.init = 16'h0100;
    LUT4 i1_3_lut_adj_549 (.A(fsm_state[1]), .B(fsm_state[2]), .C(\read_cycles_count[1] ), 
         .Z(n28858)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_549.init = 16'h8080;
    LUT4 i20_4_lut (.A(n31951), .B(n31877), .C(is_writing), .D(n6), 
         .Z(clk_c_enable_513)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (((D)+!C)+!B)) */ ;
    defparam i20_4_lut.init = 16'hf535;
    LUT4 i27796_4_lut (.A(is_writing), .B(n31877), .C(\qspi_data_byte_idx[1] ), 
         .D(n6738), .Z(n29534)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(238[18] 244[12])
    defparam i27796_4_lut.init = 16'h7557;
    LUT4 i1_2_lut_4_lut (.A(spi_clk_pos), .B(n32043), .C(n18029), .D(n33479), 
         .Z(n26213)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[25:140])
    defparam i1_2_lut_4_lut.init = 16'h00a3;
    LUT4 i27379_3_lut_4_lut (.A(\instr_data[8] ), .B(n31931), .C(n31877), 
         .D(n29082), .Z(instr_data_15__N_1959[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam i27379_3_lut_4_lut.init = 16'h8f80;
    LUT4 i27385_3_lut_4_lut (.A(\instr_data[11] ), .B(n31931), .C(n31877), 
         .D(n29091), .Z(instr_data_15__N_1959[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam i27385_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_4_lut_adj_550 (.A(fsm_state[0]), .B(stop_txn_reg), .C(fsm_state[1]), 
         .D(fsm_state[2]), .Z(n27620)) /* synthesis lut_function=(A (B)+!A (B+(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(135[18] 214[12])
    defparam i1_4_lut_adj_550.init = 16'hdccd;
    LUT4 i16036_3_lut_rep_672_4_lut_3_lut (.A(n33479), .B(n5), .C(spi_clk_pos), 
         .Z(n31877)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(231[22] 237[16])
    defparam i16036_3_lut_rep_672_4_lut_3_lut.init = 16'h8c8c;
    LUT4 i1_4_lut_adj_551 (.A(n1027), .B(n26213), .C(n31919), .D(n5), 
         .Z(n27183)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(209[30] 211[24])
    defparam i1_4_lut_adj_551.init = 16'h8000;
    LUT4 mux_2877_i3_4_lut_else_2_lut (.A(nibbles_remaining_c[2]), .B(n33479), 
         .C(fsm_state[2]), .D(fsm_state[0]), .Z(n32057)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_2877_i3_4_lut_else_2_lut.init = 16'h8b88;
    LUT4 n9_bdd_3_lut_28601_4_lut (.A(fsm_state[1]), .B(n31951), .C(spi_in_buffer[1]), 
         .D(n31950), .Z(n31591)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(167[102:126])
    defparam n9_bdd_3_lut_28601_4_lut.init = 16'hf1e0;
    LUT4 n18610_bdd_3_lut_27976_4_lut (.A(n31971), .B(n33479), .C(rst_reg_n), 
         .D(\qspi_data_in[0] ), .Z(n30602)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam n18610_bdd_3_lut_27976_4_lut.init = 16'h4000;
    LUT4 n18610_bdd_3_lut_28529_4_lut (.A(n31971), .B(n33479), .C(rst_reg_n), 
         .D(\qspi_data_in[2] ), .Z(n31582)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam n18610_bdd_3_lut_28529_4_lut.init = 16'h4000;
    LUT4 n18610_bdd_3_lut_28520_4_lut (.A(n31971), .B(n33479), .C(rst_reg_n), 
         .D(\qspi_data_in[3] ), .Z(n31576)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(234[26] 236[20])
    defparam n18610_bdd_3_lut_28520_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_4_lut (.A(n33479), .B(n31918), .C(n31736), .D(n28648), 
         .Z(n356[1])) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(168[29:51])
    defparam i1_4_lut_4_lut.init = 16'h5450;
    LUT4 i1_2_lut_4_lut_adj_552 (.A(qspi_data_ready), .B(n31976), .C(instr_fetch_running), 
         .D(n32020), .Z(n27680)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_4_lut_adj_552.init = 16'h8000;
    LUT4 n9_bdd_4_lut_28525 (.A(n31928), .B(\qspi_data_in[3] ), .C(spi_in_buffer[3]), 
         .D(rst_reg_n), .Z(n31574)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam n9_bdd_4_lut_28525.init = 16'he4a0;
    LUT4 i4811_2_lut_rep_705_4_lut (.A(qspi_data_ready), .B(n31976), .C(instr_fetch_running), 
         .D(\instr_addr_23__N_318[0] ), .Z(n31910)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i4811_2_lut_rep_705_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_553 (.A(qspi_data_ready), .B(n31976), .C(instr_fetch_running), 
         .D(n31994), .Z(n27776)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_4_lut_adj_553.init = 16'hff7f;
    LUT4 i1_2_lut_4_lut_adj_554 (.A(qspi_data_ready), .B(n31976), .C(instr_fetch_running), 
         .D(n31991), .Z(n27772)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_4_lut_adj_554.init = 16'hff7f;
    LUT4 i1_2_lut_4_lut_adj_555 (.A(qspi_data_ready), .B(n31976), .C(instr_fetch_running), 
         .D(n31990), .Z(n27780)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(122[12] 215[8])
    defparam i1_2_lut_4_lut_adj_555.init = 16'hff7f;
    LUT4 i27850_2_lut_4_lut_4_lut (.A(n31951), .B(is_writing), .C(n31877), 
         .D(n31895), .Z(clk_c_enable_517)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (C (D))))) */ ;
    defparam i27850_2_lut_4_lut_4_lut.init = 16'h1ddd;
    LUT4 i1_3_lut_adj_556 (.A(debug_stop_txn), .B(stop_txn_now_N_2363), 
         .C(stop_txn_reg), .Z(stop_txn_reg_N_2360)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_3_lut_adj_556.init = 16'h0202;
    LUT4 i27799_3_lut_4_lut (.A(n32036), .B(nibbles_remaining[0]), .C(n1084), 
         .D(n4342[1]), .Z(n18667)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam i27799_3_lut_4_lut.init = 16'h0d02;
    LUT4 mux_2877_i2_4_lut (.A(n1027), .B(nibbles_remaining_c[1]), .C(n33479), 
         .D(n31919), .Z(n4342[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(205[34] 208[28])
    defparam mux_2877_i2_4_lut.init = 16'hcac0;
    LUT4 n9_bdd_4_lut (.A(n31928), .B(\qspi_data_in[2] ), .C(spi_in_buffer[2]), 
         .D(rst_reg_n), .Z(n31580)) /* synthesis lut_function=(A (C)+!A (B (D))) */ ;
    defparam n9_bdd_4_lut.init = 16'he4a0;
    PFUMX i28609 (.BLUT(n32057), .ALUT(n32058), .C0(fsm_state[1]), .Z(n32059));
    L6MUX21 i28541 (.D0(n31595), .D1(n31592), .SD(n29534), .Z(data_out_7__N_2177[1]));
    PFUMX i28539 (.BLUT(n31594), .ALUT(n31593), .C0(n31877), .Z(n31595));
    PFUMX i28615 (.BLUT(n32067), .ALUT(n32068), .C0(\writing_N_164[3] ), 
          .Z(n32069));
    PFUMX i28537 (.BLUT(n29072), .ALUT(n31591), .C0(n32056), .Z(n31592));
    
endmodule
//
// Verilog Description of module tinyqv_cpu
//

module tinyqv_cpu (clk_c, \data_from_read[2] , counter_hi, was_early_branch, 
            data_to_write, qv_data_write_n, rd, rs1, \instr_addr_23__N_318[0] , 
            addr, \addr[24] , \addr[23] , \addr[22] , \addr[21] , 
            \addr[20] , \addr[19] , \addr[18] , \addr[17] , \addr[16] , 
            \addr[15] , \addr[14] , \addr[13] , \addr[12] , \addr[11] , 
            \addr[10] , \addr[9] , \addr[8] , \addr[7] , \addr[6] , 
            \addr[5] , \addr[4] , \addr[3] , \addr[2] , \addr[1] , 
            \instr_write_offset[3] , debug_data_continue, is_load, n31860, 
            rs2, \instr_len[2] , n31869, debug_instr_valid, \pc[1] , 
            \pc[2] , n2565, n31770, n2208, n31742, \data_out_slice[3] , 
            n31879, n19, n31885, \peri_data_out[9] , n4, \mem_data_from_read[20] , 
            \mem_data_from_read[16] , n31865, n31944, n2524, n2504, 
            n31958, VCC_net, rst_reg_n, n31792, data_txn_len, instr_data, 
            n31997, n18241, n32033, n31902, \pc[5] , \pc[13] , n28964, 
            n10467, \peri_data_out[6] , n31867, n4_adj_11, n26216, 
            n4263, \pc[9] , \imm[23] , \imm[22] , \imm[21] , \imm[20] , 
            \imm[19] , \imm[18] , \imm[17] , \imm[16] , \imm[15] , 
            \imm[14] , \imm[13] , \imm[12] , \imm[11] , \imm[10] , 
            \imm[9] , \imm[8] , \imm[7] , \imm[6] , \imm[5] , \imm[4] , 
            \imm[3] , \imm[2] , \imm[1] , n33488, n10499, n31730, 
            instr_active, \txn_len[1] , n32035, n32019, n31900, n26266, 
            n31901, n80, n31868, n31978, n31847, n27702, n13146, 
            instr_complete_N_1647, instr_fetch_running, n2152, \early_branch_addr[2] , 
            \instr_addr[2] , n31863, \instr_data[1][7] , \instr_data[2][7] , 
            n31853, debug_stop_txn_N_2147, instr_fetch_running_N_945, 
            qspi_data_ready, n32052, n58, n31849, \instr_data[3][7] , 
            n32055, stall_core, start_instr, n31741, n8, \debug_rd_3__N_405[31] , 
            \next_pc_for_core[6] , n2136, n2514, \next_pc_for_core[4] , 
            n31940, n32006, \next_pc_for_core[9] , \next_pc_for_core[13] , 
            \next_pc_for_core[10] , \next_pc_for_core[14] , \peri_data_out[10] , 
            n31761, \mem_data_from_read[19] , \mem_data_from_read[23] , 
            cycle, data_out_3__N_1385, is_ret_de, n31990, n31991, 
            n31994, n31939, n31934, n32027, n26205, clk_c_enable_268, 
            n31941, \next_pc_for_core[8] , \next_pc_for_core[12] , data_ready_r, 
            n31905, n28760, \next_pc_for_core[3] , \pc[23] , \pc[22] , 
            \pc[21] , \pc[20] , \pc[19] , \pc[18] , \pc[17] , \pc[16] , 
            \pc[15] , \pc[14] , \pc[12] , \pc[11] , \pc[10] , \pc[8] , 
            \pc[7] , \next_pc_for_core[5] , \pc[6] , \pc[4] , \next_pc_for_core[7] , 
            n84, \next_pc_for_core[11] , \next_pc_for_core[15] , \pc[3] , 
            \early_branch_addr[5] , n32016, \next_pc_for_core[16] , \early_branch_addr[6] , 
            \next_pc_for_core[17] , \next_pc_for_core[18] , \next_pc_for_core[19] , 
            \next_pc_for_core[20] , \early_branch_addr[4] , \early_branch_addr[3] , 
            \early_branch_addr[7] , \early_branch_addr[8] , \early_branch_addr[9] , 
            \early_branch_addr[10] , \next_pc_for_core[21] , \early_branch_addr[11] , 
            \early_branch_addr[12] , \early_branch_addr[13] , \early_branch_addr[14] , 
            \early_branch_addr[15] , \next_pc_for_core[22] , \early_branch_addr[16] , 
            \early_branch_addr[17] , \next_pc_for_core[23] , n32034, n31880, 
            \gpio_out_sel_7__N_13[0] , n31725, \early_branch_addr[18] , 
            \early_branch_addr[19] , \early_branch_addr[20] , \early_branch_addr[21] , 
            \early_branch_addr[22] , \early_branch_addr[23] , n31864, 
            n1724, n31935, n32020, n27310, n31736, n33479, n31906, 
            n1176, n32021, n32022, n18588, clk_c_enable_36, mem_data_ready, 
            data_ready, n31936, n31962, n31925, n31927, n26282, 
            n31964, n31967, n31735, n31164, n27680, n32017, n31163, 
            clk_c_enable_390, \mem_data_from_read[7] , \data_from_read[7] , 
            \mem_data_from_read[3] , \data_from_read[3] , instr_fetch_running_N_943, 
            \mem_data_from_read[0] , \data_from_read[0] , \mem_data_from_read[4] , 
            \data_from_read[4] , \mem_data_from_read[8] , \data_from_read[8] , 
            \mem_data_from_read[12] , \data_from_read[12] , \mem_data_from_read[1] , 
            \data_from_read[1] , \mem_data_from_read[5] , \data_from_read[5] , 
            n31932, n31922, n31819, \mem_data_from_read[24] , \mem_data_from_read[28] , 
            \mem_data_from_read[25] , \mem_data_from_read[29] , \peri_data_out[11] , 
            \mem_data_from_read[26] , \mem_data_from_read[30] , \mem_data_from_read[27] , 
            \mem_data_from_read[31] , n31910, n31942, \mem_data_from_read[18] , 
            \mem_data_from_read[22] , gpio_out_sel, n14, n14_adj_12, 
            n31961, n5171, n28686, n18680, \qspi_data_buf[9] , \qspi_data_buf[13] , 
            n27776, n27772, n27780, \qspi_data_buf[11] , \qspi_data_buf[15] , 
            \qspi_data_buf[10] , \qspi_data_buf[14] , n31899, clk_c_enable_273, 
            clk_c_enable_357, clk_c_enable_349, n32003, clk_c_enable_259, 
            clk_c_enable_360, n31904, n10573, instr_fetch_stopped, n31841, 
            n15604, n29004, n31798, clk_c_enable_234, \ui_in_sync[0] , 
            n1160, \alu_b_in[3] , debug_rd, \ui_in_sync[1] , \next_fsm_state_3__N_3015[3] , 
            fsm_state, accum, d_3__N_1868, n31929, \mul_out[1] , \mul_out[2] , 
            \mul_out[3] , n31963, next_bit, n28800, n31389, alu_b_in_3__N_1504, 
            \mem_data_from_read[17] , \mem_data_from_read[21] , n29162, 
            n18086, \csr_read_3__N_1447[2] , GND_net, \next_accum[5] , 
            \next_accum[6] , \next_accum[7] , \next_accum[8] , \next_accum[9] , 
            \next_accum[10] , \next_accum[11] , \next_accum[12] , \next_accum[13] , 
            \next_accum[14] , \next_accum[15] , \next_accum[16] , \next_accum[17] , 
            \next_accum[18] , \next_accum[19] , \next_accum[4] , n12, 
            n11, n9, n8_adj_13, \registers[5][7] , \registers[6][7] , 
            \registers[7][7] , n27762, n29747, n4_adj_14) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    input \data_from_read[2] ;
    output [4:2]counter_hi;
    output was_early_branch;
    output [31:0]data_to_write;
    output [1:0]qv_data_write_n;
    output [3:0]rd;
    output [3:0]rs1;
    output \instr_addr_23__N_318[0] ;
    output [27:0]addr;
    output \addr[24] ;
    output \addr[23] ;
    output \addr[22] ;
    output \addr[21] ;
    output \addr[20] ;
    output \addr[19] ;
    output \addr[18] ;
    output \addr[17] ;
    output \addr[16] ;
    output \addr[15] ;
    output \addr[14] ;
    output \addr[13] ;
    output \addr[12] ;
    output \addr[11] ;
    output \addr[10] ;
    output \addr[9] ;
    output \addr[8] ;
    output \addr[7] ;
    output \addr[6] ;
    output \addr[5] ;
    output \addr[4] ;
    output \addr[3] ;
    output \addr[2] ;
    output \addr[1] ;
    output \instr_write_offset[3] ;
    output debug_data_continue;
    output is_load;
    output n31860;
    output [3:0]rs2;
    output \instr_len[2] ;
    output n31869;
    output debug_instr_valid;
    output \pc[1] ;
    output \pc[2] ;
    output n2565;
    input n31770;
    output n2208;
    output n31742;
    input \data_out_slice[3] ;
    output n31879;
    output n19;
    output n31885;
    input \peri_data_out[9] ;
    output n4;
    input \mem_data_from_read[20] ;
    input \mem_data_from_read[16] ;
    output n31865;
    output n31944;
    input n2524;
    input n2504;
    output n31958;
    input VCC_net;
    input rst_reg_n;
    input n31792;
    input [1:0]data_txn_len;
    input [15:0]instr_data;
    output n31997;
    input n18241;
    output n32033;
    output n31902;
    output \pc[5] ;
    output \pc[13] ;
    input n28964;
    output n10467;
    input \peri_data_out[6] ;
    output n31867;
    input n4_adj_11;
    output n26216;
    output n4263;
    output \pc[9] ;
    output \imm[23] ;
    output \imm[22] ;
    output \imm[21] ;
    output \imm[20] ;
    output \imm[19] ;
    output \imm[18] ;
    output \imm[17] ;
    output \imm[16] ;
    output \imm[15] ;
    output \imm[14] ;
    output \imm[13] ;
    output \imm[12] ;
    output \imm[11] ;
    output \imm[10] ;
    output \imm[9] ;
    output \imm[8] ;
    output \imm[7] ;
    output \imm[6] ;
    output \imm[5] ;
    output \imm[4] ;
    output \imm[3] ;
    output \imm[2] ;
    output \imm[1] ;
    input n33488;
    output n10499;
    output n31730;
    input instr_active;
    output \txn_len[1] ;
    output n32035;
    output n32019;
    output n31900;
    output n26266;
    output n31901;
    output n80;
    output n31868;
    output n31978;
    output n31847;
    input n27702;
    output n13146;
    output instr_complete_N_1647;
    output instr_fetch_running;
    input n2152;
    input \early_branch_addr[2] ;
    output \instr_addr[2] ;
    output n31863;
    output \instr_data[1][7] ;
    output \instr_data[2][7] ;
    output n31853;
    output debug_stop_txn_N_2147;
    input instr_fetch_running_N_945;
    input qspi_data_ready;
    input n32052;
    output n58;
    output n31849;
    output \instr_data[3][7] ;
    output n32055;
    output stall_core;
    output start_instr;
    output n31741;
    output n8;
    output \debug_rd_3__N_405[31] ;
    input \next_pc_for_core[6] ;
    output n2136;
    output n2514;
    input \next_pc_for_core[4] ;
    input n31940;
    output n32006;
    input \next_pc_for_core[9] ;
    input \next_pc_for_core[13] ;
    input \next_pc_for_core[10] ;
    input \next_pc_for_core[14] ;
    input \peri_data_out[10] ;
    input n31761;
    input \mem_data_from_read[19] ;
    input \mem_data_from_read[23] ;
    output [1:0]cycle;
    output data_out_3__N_1385;
    input is_ret_de;
    output n31990;
    output n31991;
    output n31994;
    output n31939;
    input n31934;
    input n32027;
    output n26205;
    output clk_c_enable_268;
    output n31941;
    input \next_pc_for_core[8] ;
    input \next_pc_for_core[12] ;
    input data_ready_r;
    input n31905;
    output n28760;
    input \next_pc_for_core[3] ;
    output \pc[23] ;
    output \pc[22] ;
    output \pc[21] ;
    output \pc[20] ;
    output \pc[19] ;
    output \pc[18] ;
    output \pc[17] ;
    output \pc[16] ;
    output \pc[15] ;
    output \pc[14] ;
    output \pc[12] ;
    output \pc[11] ;
    output \pc[10] ;
    output \pc[8] ;
    output \pc[7] ;
    input \next_pc_for_core[5] ;
    output \pc[6] ;
    output \pc[4] ;
    input \next_pc_for_core[7] ;
    input n84;
    input \next_pc_for_core[11] ;
    input \next_pc_for_core[15] ;
    output \pc[3] ;
    input \early_branch_addr[5] ;
    input n32016;
    input \next_pc_for_core[16] ;
    input \early_branch_addr[6] ;
    input \next_pc_for_core[17] ;
    input \next_pc_for_core[18] ;
    input \next_pc_for_core[19] ;
    input \next_pc_for_core[20] ;
    input \early_branch_addr[4] ;
    input \early_branch_addr[3] ;
    input \early_branch_addr[7] ;
    input \early_branch_addr[8] ;
    input \early_branch_addr[9] ;
    input \early_branch_addr[10] ;
    input \next_pc_for_core[21] ;
    input \early_branch_addr[11] ;
    input \early_branch_addr[12] ;
    input \early_branch_addr[13] ;
    input \early_branch_addr[14] ;
    input \early_branch_addr[15] ;
    input \next_pc_for_core[22] ;
    input \early_branch_addr[16] ;
    input \early_branch_addr[17] ;
    input \next_pc_for_core[23] ;
    output n32034;
    input n31880;
    output \gpio_out_sel_7__N_13[0] ;
    output n31725;
    input \early_branch_addr[18] ;
    input \early_branch_addr[19] ;
    input \early_branch_addr[20] ;
    input \early_branch_addr[21] ;
    input \early_branch_addr[22] ;
    input \early_branch_addr[23] ;
    input n31864;
    input n1724;
    output n31935;
    output n32020;
    input n27310;
    input n31736;
    input n33479;
    input n31906;
    output n1176;
    output n32021;
    output n32022;
    output n18588;
    output clk_c_enable_36;
    input mem_data_ready;
    input data_ready;
    output n31936;
    output n31962;
    output n31925;
    output n31927;
    input n26282;
    output n31964;
    output n31967;
    output n31735;
    input n31164;
    input n27680;
    input n32017;
    output n31163;
    output clk_c_enable_390;
    input \mem_data_from_read[7] ;
    input \data_from_read[7] ;
    input \mem_data_from_read[3] ;
    input \data_from_read[3] ;
    input instr_fetch_running_N_943;
    input \mem_data_from_read[0] ;
    input \data_from_read[0] ;
    input \mem_data_from_read[4] ;
    input \data_from_read[4] ;
    input \mem_data_from_read[8] ;
    input \data_from_read[8] ;
    input \mem_data_from_read[12] ;
    input \data_from_read[12] ;
    input \mem_data_from_read[1] ;
    input \data_from_read[1] ;
    input \mem_data_from_read[5] ;
    input \data_from_read[5] ;
    output n31932;
    input n31922;
    output n31819;
    input \mem_data_from_read[24] ;
    input \mem_data_from_read[28] ;
    input \mem_data_from_read[25] ;
    input \mem_data_from_read[29] ;
    input \peri_data_out[11] ;
    input \mem_data_from_read[26] ;
    input \mem_data_from_read[30] ;
    input \mem_data_from_read[27] ;
    input \mem_data_from_read[31] ;
    input n31910;
    input n31942;
    input \mem_data_from_read[18] ;
    input \mem_data_from_read[22] ;
    input [7:6]gpio_out_sel;
    output n14;
    output n14_adj_12;
    input n31961;
    output n5171;
    input n28686;
    output n18680;
    input \qspi_data_buf[9] ;
    input \qspi_data_buf[13] ;
    input n27776;
    input n27772;
    input n27780;
    input \qspi_data_buf[11] ;
    input \qspi_data_buf[15] ;
    input \qspi_data_buf[10] ;
    input \qspi_data_buf[14] ;
    input n31899;
    output clk_c_enable_273;
    output clk_c_enable_357;
    output clk_c_enable_349;
    input n32003;
    output clk_c_enable_259;
    output clk_c_enable_360;
    output n31904;
    input n10573;
    input instr_fetch_stopped;
    output n31841;
    output n15604;
    output n29004;
    output n31798;
    input clk_c_enable_234;
    input \ui_in_sync[0] ;
    output n1160;
    input \alu_b_in[3] ;
    output [3:0]debug_rd;
    input \ui_in_sync[1] ;
    input \next_fsm_state_3__N_3015[3] ;
    input [3:0]fsm_state;
    output [15:0]accum;
    output [19:0]d_3__N_1868;
    output n31929;
    input \mul_out[1] ;
    input \mul_out[2] ;
    input \mul_out[3] ;
    output n31963;
    input next_bit;
    output n28800;
    input n31389;
    output alu_b_in_3__N_1504;
    input \mem_data_from_read[17] ;
    input \mem_data_from_read[21] ;
    input n29162;
    output n18086;
    output \csr_read_3__N_1447[2] ;
    input GND_net;
    input \next_accum[5] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[4] ;
    output n12;
    output n11;
    output n9;
    output n8_adj_13;
    output \registers[5][7] ;
    output \registers[6][7] ;
    output \registers[7][7] ;
    output n27762;
    output n29747;
    input n4_adj_14;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire is_alu_imm, clk_c_enable_358, n31980, is_alu_imm_de, n32277, 
        n32278, interrupt_core, clk_c_enable_134, n31744;
    wire [3:0]alu_op;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(114[15:21])
    
    wire clk_c_enable_347;
    wire [3:0]alu_op_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(64[16:25])
    wire [31:0]imm;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(100[16:19])
    
    wire clk_c_enable_212;
    wire [31:0]n3546;
    
    wire clk_c_enable_20, debug_early_branch, n30773, n30770, n4281, 
        n30774, clk_c_enable_184;
    wire [3:0]data_out_slice;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(230[16:30])
    
    wire clk_c_enable_224;
    wire [1:0]data_write_n_1__N_369;
    wire [2:0]additional_mem_ops;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(120[15:33])
    wire [2:0]additional_mem_ops_2__N_749;
    
    wire clk_c_enable_448;
    wire [3:0]n1764;
    wire [2:1]instr_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(113[15:24])
    
    wire clk_c_enable_30, n31789;
    wire [2:0]mem_op;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(115[15:21])
    
    wire clk_c_enable_325;
    wire [2:0]mem_op_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(65[16:25])
    wire [3:0]n2644;
    wire [1:0]qv_data_read_n;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/tinyqv.v(65[15:29])
    
    wire clk_c_enable_117, n26972;
    wire [15:0]n6;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire clk_c_enable_343;
    wire [63:0]instr_data_0__15__N_638;
    
    wire data_ready_sync, data_ready_core;
    wire [2:0]instr_write_offset_3__N_934;
    
    wire clk_c_enable_107;
    wire [27:0]addr_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(131[17:25])
    
    wire n30765, n30763, n30766;
    wire [27:0]addr_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(52[17:21])
    
    wire n27068;
    wire [1:0]n699;
    
    wire n26290;
    wire [3:1]next_instr_write_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[16:39])
    wire [22:0]instr_addr_23__N_318;
    
    wire clk_c_enable_108, data_continue_N_963, no_write_in_progress, 
        clk_c_enable_109, no_write_in_progress_N_471, is_load_de, n31472, 
        n31471, n31473, n26971;
    wire [3:0]rs1_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(117[15:18])
    
    wire is_store, is_store_de;
    wire [3:0]n2243;
    
    wire n31791;
    wire [3:0]rd_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(119[15:17])
    
    wire n31439, n31438, n19_c, debug_instr_valid_N_436, n31194, n31436, 
        n31845, n31437;
    wire [3:1]next_pc_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[16:30])
    
    wire n31424, n31423, n31425;
    wire [2:0]n4322;
    
    wire n13255, clk_c_enable_157, clk_c_enable_161, clk_c_enable_165, 
        clk_c_enable_169, clk_c_enable_173, clk_c_enable_177, clk_c_enable_181, 
        n26, n31722, n4271, n4279, n29428;
    wire [31:0]n3381;
    wire [15:0]n5223;
    wire [31:0]n3422;
    
    wire n32071, n32070, n32183, n31719, n26764, n4277;
    wire [31:0]n3271;
    
    wire n31813;
    wire [15:0]n2525;
    
    wire n27746, n31852, n32075;
    wire [15:0]n2505;
    
    wire n32074, n31732, n29371;
    wire [15:0]n21;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire n32079, n31416, n31415, n31417;
    wire [15:0]n27;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    wire [15:0]n31;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(372[16:26])
    
    wire n32078, n13, n32184, n29658, n32185, load_started, address_ready, 
        n844, n43, n31838, n2134, n32064, n32065, n32066, n32280, 
        n22, n35, n30803, n31418, n31406, n31405, n31407, n30748, 
        n30747, n30749, n29318, n26119, n24, n22_adj_3135, n9894, 
        n4_adj_3136, n28140, is_jal, is_jal_de, n32063, n29759, 
        n29063;
    wire [15:0]n2163;
    wire [31:0]instr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(47[17:22])
    
    wire n31310, n31311, n30762, n31684;
    wire [15:0]n2143;
    wire [31:0]n3505;
    
    wire n4285, n10068, n31315, n31316, n31743, n31740, n30804, 
        n32072, n31408;
    wire [2:0]c_2__N_1861;
    
    wire n30767, n30775, n31687;
    wire [3:2]addr_offset;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(121[15:26])
    wire [1:0]n33;
    
    wire n31884, n31686, clk_c_enable_214, n30840, clk_c_enable_221, 
        n30709, n27018, n27846, n31748, n26948, n28150, n28152, 
        n30805, n30802, n33484;
    wire [59:0]debug_branch_N_442;
    
    wire n27460;
    wire [30:0]n5121;
    
    wire n31734, is_alu_reg, is_alu_reg_de, n30743, n30742, n30744, 
        n31796, n31846;
    wire [2:0]additional_mem_ops_de;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(70[16:37])
    
    wire clk_c_enable_287, n28006, n28332, n27862, n41;
    wire [3:0]n155;
    
    wire n31820;
    wire [3:0]alu_op_3__N_1170;
    
    wire n32042, n4_adj_3138, n31851, n28260, n9_c, n26770, n27726, 
        n30838, n31866, n1, n30839, n30835, n29023;
    wire [31:0]n3458;
    
    wire is_jalr, is_jalr_de, n27832, n7103, n27604, n29025, n31822, 
        n15_adj_3139, is_branch, is_branch_de, n31747, n27286, debug_ret, 
        n31318, n31319, n29033, n31738, n27750, n29051, n26693, 
        n25, clk_c_enable_289, clk_c_enable_303, clk_c_enable_305, clk_c_enable_319, 
        clk_c_enable_321, clk_c_enable_342, mem_op_increment_reg, mem_op_increment_reg_de, 
        n27942, n31720;
    wire [31:0]n3195;
    
    wire n17976, n37, n27818, n31777, n31760, n24_adj_3140, n30, 
        debug_stop_txn_N_2148, n31745, n27606, n10112, n16;
    wire [31:0]n2982;
    
    wire n30836, n31778;
    wire [31:0]n3304;
    
    wire n28284, n27056, n31965, n12_c, n19_adj_3141, n28018, n31818, 
        n31772, n28020, n31774, n31831, n31972, n30708;
    wire [3:0]alu_op_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[16:25])
    
    wire n32029, n18324, n26175, n32044, n31888, n27796, n2500, 
        is_system, is_system_de, is_lui, is_lui_de, n17, is_auipc, 
        is_auipc_de, n28912, clk_c_enable_370, n6411, data_ready_latch, 
        clk_c_enable_375, n27110, n29597, n30707, n30706, n31718, 
        n29596, n31754;
    wire [3:0]n5677;
    wire [59:0]debug_rd_3__N_405;
    
    wire n32001, n9033;
    wire [59:0]debug_branch_N_446;
    
    wire n31848, n28864, n29595, n27480, n29594, n32054, n29147;
    wire [23:1]return_addr;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(135[17:28])
    wire [1:0]n34;
    
    wire n31809, n27946, debug_rd_3__N_1575, n29049, n29490, n29575, 
        n29028, n31715, n29026, n29574, n29573, n29057, n29020, 
        n29572, n29018, n29568, n29567, n28881, n27724, n29566, 
        n29565, n29561, n29560, n29559, n29558, n31714, n26794, 
        n149, n29392, n31197, n31196, n31835, n31198;
    wire [12:0]n5081;
    
    wire n33486, n29337, n17_adj_3142, n20, n29385, n26782, n15_adj_3143, 
        n20_adj_3144, n31834, n30_adj_3145, n28, n31987, n31892, 
        n31948, n29136, n31894, n32062, n31914, n13_adj_3146, n31875, 
        n26113, n31817, n8_adj_3147, n7, n31786, n32, n31802, 
        n31769, is_lui_N_1365, n31915, n31795;
    wire [59:0]debug_branch_N_840;
    wire [3:0]timer_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(143[16:26])
    
    wire is_timer_addr;
    wire [3:0]debug_branch_N_450;
    
    wire n29148, n209, n31955, n26829;
    wire [3:0]n2630;
    
    wire n2812, n32061, n26478, n17998, n28074, n28080, n29047, 
        n29045, n29027, n28086, n28092, n13248, n29029, n28098, 
        n28104, n31764, n28110, n28116, n31733;
    wire [31:0]n3340;
    
    wire n26788, debug_rd_3__N_413, n29192, n10486, n32039, n28708, 
        n15_adj_3148;
    wire [1:0]cycle_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(58[15:20])
    
    wire n31737, n29160, load_top_bit, n29166;
    wire [2:0]n36;
    
    wire n26776, n28028, n27972, n26648, n29210, n27966, n26800;
    wire [31:0]n3234;
    
    wire n27978, n30171, n30170, n31200, n26310, n31937, n29737, 
        n29739, n29663, n29665, n31762, n31755;
    wire [3:0]n2621;
    
    wire n157_adj_3150, n31999, n29330, n31763, n31441, n29333, 
        n32007, n29240;
    wire [3:0]n234;
    wire [3:0]n2222;
    
    wire n31871;
    wire [31:0]mtimecmp;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(30[16:24])
    
    wire mtimecmp_2__N_1939, mtimecmp_3__N_1935, mtimecmp_1__N_1941, mtimecmp_0__N_1943, 
        clk_c_enable_527;
    wire [1:0]pc_2__N_932;
    
    wire n31766, n32050;
    wire [3:0]n5;
    wire [3:0]n2;
    
    wire n2138, n31975, n6668;
    wire [3:0]n2589;
    wire [3:0]n2597;
    
    wire n2808, n31120, n31121, n26993, n28182;
    wire [20:0]n1742;
    
    wire alu_a_in_3__N_1552, n29220, n31773, n2498, n26871;
    wire [3:0]n2232;
    
    wire n209_adj_3151, n157_adj_3152, n29012, n26889, n26905;
    wire [20:0]pc_23__N_911;
    
    wire n26883, n26877;
    wire [3:0]data_rs2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(84[16:24])
    wire [3:0]n92;
    
    wire n27614, n27994, n32015;
    wire [20:0]n1215;
    
    wire n31117, n31118;
    wire [1:0]n5014;
    
    wire n26827;
    wire [3:0]n1720;
    
    wire n29562, n29563, n26814, n32076, n27672, n31898, n26807, 
        n29569, n29570, n31830;
    wire [3:0]n1725;
    
    wire n26996, n31119, n24_adj_3160, n29043, n31808, n29576, n29577, 
        n29598, n29599, n26995, n26997, n149_adj_3161, n225, n10904;
    wire [3:0]n2607;
    
    wire n2810;
    wire [2:0]additional_mem_ops_2__N_1132;
    
    wire n31803, n28174;
    wire [3:0]n2602;
    
    wire n29400, n26821, n31799, n27998, n31814, n31402, n31807, 
        n27246, n9538;
    wire [3:0]n5624;
    wire [3:0]n5659;
    
    wire n29041, n29019, n8302, n29048, n29375, n32026, load_done, 
        instr_complete_N_1651, n30169, n30168, data_ready_ext, n30167, 
        n31850, n30166, n18518, n30165, n31816, n31815, n28871, 
        n28412, n28400, n28410, n28398, load_done_N_1741, n9710, 
        n28032, n30609, n26202, n31805, n31840, n31823, n28444, 
        n30610, n27804, n24_adj_3162, n28898, n824, n31824, n31821, 
        n31800, n2804, n28060, n4_adj_3163, n28366, n3, n28156, 
        n29193, n10899, n4269, n30611, n27214, n28496, n28498, 
        n28494, n28486, n28474, n28492, n28480, n29194, n31728, 
        n27734, n27744, n31785, n227, n29149, n29656, n29657, 
        n12_adj_3164, n30_adj_3165, n29135, n29733, n29734, n31768, 
        n226, n29137, n8289, n31790, n29, n29652, n29653, n29293, 
        n29654, n29655, n29659, n29660;
    wire [3:0]n108;
    
    wire n32046, n28222, n225_adj_3166, n28204, n29215, n31861, 
        n31903, n32049;
    wire [3:0]csr_read_3__N_1443;
    
    wire n32040;
    wire [3:0]data_rs1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(83[16:24])
    
    wire n31837, n22_adj_3167;
    wire [2:0]mem_op_2__N_1114;
    
    wire n31804, n31806, n32_adj_3168, n10, n23, n31812, n31833, 
        n27688, n29190, n4_adj_3169, n33493, n30950, n31966, n26656, 
        n26899, n28008, n27738, n27728;
    wire [2:0]n1764_adj_3181;
    
    wire n30949, n30837, n16_adj_3171, n26_adj_3172, n32282, n30764, 
        n30772, n27694, n27850, n29006, n30760, n30761, n31685, 
        n29056, n30741, n31784, n30947, n30746, n27576, n31949, 
        n27956, n27960, n32279, n30759, n27892, n27868, n27922, 
        n31682, n27880, n28282, n27928, n27810, n27904, n30771, 
        n28128, n32281, timer_interrupt, time_pulse_r, clk_c_enable_249, 
        n31913;
    wire [3:0]mtime_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(29[16:25])
    
    wire cy, n31876, n31957, n31946, clk_c_enable_449;
    wire [6:0]cycle_count_wide;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(279[16:32])
    
    wire n31870, clk_c_enable_233, n31893, is_double_fault_r, mstatus_mte;
    wire [3:0]\reg_access[3] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(30[16:26])
    
    wire mstatus_mie_N_1709, n31878, mstatus_mie_N_1707, n31872, n31889, 
        n31758, is_jalr_N_1370, n28040, n27790, n27934, n28068, 
        n28054, n12_adj_3176, n27898, n27886, n27910, n27838, n27874, 
        n27824;
    
    FD1P3IX is_alu_imm_394 (.D(is_alu_imm_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_alu_imm)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_alu_imm_394.GSR = "DISABLED";
    PFUMX i28718 (.BLUT(\data_from_read[2] ), .ALUT(n32277), .C0(counter_hi[2]), 
          .Z(n32278));
    FD1P3IX interrupt_core_408 (.D(n31744), .SP(clk_c_enable_134), .CD(n31980), 
            .CK(clk_c), .Q(interrupt_core)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam interrupt_core_408.GSR = "DISABLED";
    FD1P3IX alu_op__i0 (.D(alu_op_de[0]), .SP(clk_c_enable_347), .CD(n31980), 
            .CK(clk_c), .Q(alu_op[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i0.GSR = "DISABLED";
    FD1P3AX imm_i0_i0 (.D(n3546[0]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(imm[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i0.GSR = "DISABLED";
    FD1P3IX was_early_branch_424 (.D(debug_early_branch), .SP(clk_c_enable_20), 
            .CD(n31980), .CK(clk_c), .Q(was_early_branch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(315[12] 320[8])
    defparam was_early_branch_424.GSR = "DISABLED";
    PFUMX i28062 (.BLUT(n30773), .ALUT(n30770), .C0(n4281), .Z(n30774));
    FD1P3IX data_out__i0 (.D(data_out_slice[0]), .SP(clk_c_enable_184), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i0.GSR = "DISABLED";
    FD1P3AX data_write_n_i1 (.D(data_write_n_1__N_369[1]), .SP(clk_c_enable_224), 
            .CK(clk_c), .Q(qv_data_write_n[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_write_n_i1.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i0 (.D(additional_mem_ops_2__N_749[0]), .CK(clk_c), 
            .CD(n31980), .Q(additional_mem_ops[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i0.GSR = "DISABLED";
    FD1P3AX rd_i0_i0 (.D(n1764[0]), .SP(clk_c_enable_448), .CK(clk_c), 
            .Q(rd[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i0.GSR = "DISABLED";
    FD1P3IX instr_len_i1 (.D(n31789), .SP(clk_c_enable_30), .CD(n31980), 
            .CK(clk_c), .Q(instr_len[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_len_i1.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i0 (.D(mem_op_de[0]), .SP(clk_c_enable_325), .CK(clk_c), 
            .Q(mem_op[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i0.GSR = "DISABLED";
    FD1P3AX rs1_i0_i0 (.D(n2644[0]), .SP(clk_c_enable_325), .CK(clk_c), 
            .Q(rs1[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i0.GSR = "DISABLED";
    FD1P3AX data_read_n_i0_i0 (.D(n26972), .SP(clk_c_enable_117), .CK(clk_c), 
            .Q(qv_data_read_n[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_read_n_i0_i0.GSR = "DISABLED";
    FD1P3AX instr_data_3__i1 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_343), 
            .CK(clk_c), .Q(n6[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i1.GSR = "DISABLED";
    FD1S3IX data_ready_sync_415 (.D(data_ready_core), .CK(clk_c), .CD(n31980), 
            .Q(data_ready_sync)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(235[12] 256[8])
    defparam data_ready_sync_415.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i1 (.D(instr_write_offset_3__N_934[0]), .CK(clk_c), 
            .CD(n31980), .Q(\instr_addr_23__N_318[0] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i1.GSR = "DISABLED";
    FD1P3IX data_addr__i0 (.D(addr_out[0]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(addr[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i0.GSR = "DISABLED";
    PFUMX i28058 (.BLUT(n30765), .ALUT(n30763), .C0(n4281), .Z(n30766));
    FD1P3IX data_addr__i27 (.D(addr_out[27]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(addr[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i27.GSR = "DISABLED";
    FD1P3IX data_addr__i26 (.D(addr_out[26]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(addr_c[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i26.GSR = "DISABLED";
    FD1P3IX data_addr__i25 (.D(addr_out[25]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(addr_c[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i25.GSR = "DISABLED";
    FD1P3IX data_addr__i24 (.D(addr_out[24]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[24] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i24.GSR = "DISABLED";
    FD1P3IX data_addr__i23 (.D(addr_out[23]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i23.GSR = "DISABLED";
    FD1P3IX data_addr__i22 (.D(addr_out[22]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i22.GSR = "DISABLED";
    FD1P3IX data_addr__i21 (.D(addr_out[21]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i21.GSR = "DISABLED";
    FD1P3IX data_addr__i20 (.D(addr_out[20]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i20.GSR = "DISABLED";
    FD1P3IX data_addr__i19 (.D(addr_out[19]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i19.GSR = "DISABLED";
    FD1P3IX data_addr__i18 (.D(addr_out[18]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i18.GSR = "DISABLED";
    FD1P3IX data_addr__i17 (.D(addr_out[17]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[17] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i17.GSR = "DISABLED";
    FD1P3IX data_addr__i16 (.D(addr_out[16]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[16] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i16.GSR = "DISABLED";
    FD1P3IX data_addr__i15 (.D(addr_out[15]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[15] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i15.GSR = "DISABLED";
    FD1P3IX data_addr__i14 (.D(addr_out[14]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[14] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i14.GSR = "DISABLED";
    FD1P3IX data_addr__i13 (.D(addr_out[13]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[13] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i13.GSR = "DISABLED";
    FD1P3IX data_addr__i12 (.D(addr_out[12]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[12] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i12.GSR = "DISABLED";
    FD1P3IX data_addr__i11 (.D(addr_out[11]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[11] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i11.GSR = "DISABLED";
    FD1P3IX data_addr__i10 (.D(addr_out[10]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[10] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i10.GSR = "DISABLED";
    FD1P3IX data_addr__i9 (.D(addr_out[9]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[9] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i9.GSR = "DISABLED";
    FD1P3IX data_addr__i8 (.D(addr_out[8]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[8] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i8.GSR = "DISABLED";
    FD1P3IX data_addr__i7 (.D(addr_out[7]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i7.GSR = "DISABLED";
    FD1P3IX data_addr__i6 (.D(addr_out[6]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[6] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i6.GSR = "DISABLED";
    FD1P3IX data_addr__i5 (.D(addr_out[5]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[5] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i5.GSR = "DISABLED";
    FD1P3IX data_addr__i4 (.D(addr_out[4]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[4] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i4.GSR = "DISABLED";
    FD1P3IX data_addr__i3 (.D(n27068), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[3] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i3.GSR = "DISABLED";
    FD1P3IX data_addr__i2 (.D(n699[0]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[2] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i2.GSR = "DISABLED";
    FD1P3IX data_addr__i1 (.D(addr_out[1]), .SP(clk_c_enable_107), .CD(n31980), 
            .CK(clk_c), .Q(\addr[1] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam data_addr__i1.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i3 (.D(next_instr_write_offset[3]), .CK(clk_c), 
            .CD(n26290), .Q(\instr_write_offset[3] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i3.GSR = "DISABLED";
    FD1S3IX instr_write_offset__i2 (.D(instr_write_offset_3__N_934[1]), .CK(clk_c), 
            .CD(n31980), .Q(instr_addr_23__N_318[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_write_offset__i2.GSR = "DISABLED";
    FD1P3AX data_continue_420 (.D(data_continue_N_963), .SP(clk_c_enable_108), 
            .CK(clk_c), .Q(debug_data_continue)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_continue_420.GSR = "DISABLED";
    FD1P3JX no_write_in_progress_419 (.D(no_write_in_progress_N_471), .SP(clk_c_enable_109), 
            .PD(n31980), .CK(clk_c), .Q(no_write_in_progress)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam no_write_in_progress_419.GSR = "DISABLED";
    FD1P3IX is_load_393 (.D(is_load_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_load)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_load_393.GSR = "DISABLED";
    PFUMX i28474 (.BLUT(n31472), .ALUT(n31471), .C0(n31860), .Z(n31473));
    FD1P3AX data_read_n_i0_i1 (.D(n26971), .SP(clk_c_enable_117), .CK(clk_c), 
            .Q(qv_data_read_n[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_read_n_i0_i1.GSR = "DISABLED";
    FD1P3AX rs1_i0_i3 (.D(n2644[3]), .SP(clk_c_enable_325), .CK(clk_c), 
            .Q(rs1_c[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i3.GSR = "DISABLED";
    FD1P3IX is_store_396 (.D(is_store_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_store)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_store_396.GSR = "DISABLED";
    FD1P3AX rs1_i0_i2 (.D(n2644[2]), .SP(clk_c_enable_325), .CK(clk_c), 
            .Q(rs1_c[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i2.GSR = "DISABLED";
    FD1P3AX rs1_i0_i1 (.D(n2644[1]), .SP(clk_c_enable_325), .CK(clk_c), 
            .Q(rs1_c[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs1_i0_i1.GSR = "DISABLED";
    FD1P3AX rs2_i0_i0 (.D(n2243[0]), .SP(clk_c_enable_448), .CK(clk_c), 
            .Q(rs2[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i0.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i2 (.D(mem_op_de[2]), .SP(clk_c_enable_325), .CK(clk_c), 
            .Q(mem_op[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i2.GSR = "DISABLED";
    FD1P3AX mem_op_i0_i1 (.D(mem_op_de[1]), .SP(clk_c_enable_325), .CK(clk_c), 
            .Q(mem_op[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_i0_i1.GSR = "DISABLED";
    FD1P3AX instr_len_i2 (.D(n31791), .SP(clk_c_enable_347), .CK(clk_c), 
            .Q(\instr_len[2] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_len_i2.GSR = "DISABLED";
    FD1P3AX rd_i0_i3 (.D(n1764[3]), .SP(clk_c_enable_448), .CK(clk_c), 
            .Q(rd_c[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i3.GSR = "DISABLED";
    PFUMX i28456 (.BLUT(n31439), .ALUT(n31438), .C0(n31869), .Z(n19_c));
    FD1P3IX instr_valid_392 (.D(debug_instr_valid_N_436), .SP(clk_c_enable_134), 
            .CD(n31980), .CK(clk_c), .Q(debug_instr_valid)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam instr_valid_392.GSR = "DISABLED";
    FD1P3AX rd_i0_i2 (.D(n1764[2]), .SP(clk_c_enable_448), .CK(clk_c), 
            .Q(rd_c[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i2.GSR = "DISABLED";
    FD1P3AX rd_i0_i1 (.D(n1764[1]), .SP(clk_c_enable_448), .CK(clk_c), 
            .Q(rd_c[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rd_i0_i1.GSR = "DISABLED";
    PFUMX i28454 (.BLUT(n31194), .ALUT(n31436), .C0(n31845), .Z(n31437));
    LUT4 instr_len_2__bdd_4_lut (.A(\instr_len[2] ), .B(\pc[1] ), .C(instr_len[1]), 
         .D(\pc[2] ), .Z(next_pc_offset[3])) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B (C (D)))) */ ;
    defparam instr_len_2__bdd_4_lut.init = 16'hea80;
    LUT4 i1835_2_lut_3_lut_4_lut_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), 
         .C(\instr_len[2] ), .D(\pc[2] ), .Z(n2565)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A ((C (D)+!C !(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1835_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h0660;
    PFUMX i28449 (.BLUT(n31424), .ALUT(n31423), .C0(n31770), .Z(n31425));
    LUT4 i1546_2_lut_3_lut_4_lut_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), 
         .C(\instr_len[2] ), .D(\pc[2] ), .Z(n2208)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1546_2_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h6006;
    LUT4 i8_2_lut_4_lut (.A(n31742), .B(n4322[0]), .C(n4322[1]), .D(additional_mem_ops[2]), 
         .Z(n13255)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(120[15:33])
    defparam i8_2_lut_4_lut.init = 16'hfd02;
    FD1S3IX additional_mem_ops__i2 (.D(additional_mem_ops_2__N_749[2]), .CK(clk_c), 
            .CD(n31980), .Q(additional_mem_ops[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i2.GSR = "DISABLED";
    FD1S3IX additional_mem_ops__i1 (.D(additional_mem_ops_2__N_749[1]), .CK(clk_c), 
            .CD(n31980), .Q(additional_mem_ops[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam additional_mem_ops__i1.GSR = "DISABLED";
    FD1P3IX data_out__i31 (.D(\data_out_slice[3] ), .SP(clk_c_enable_157), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i31.GSR = "DISABLED";
    FD1P3IX data_out__i30 (.D(data_out_slice[2]), .SP(clk_c_enable_157), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i30.GSR = "DISABLED";
    FD1P3IX data_out__i29 (.D(data_out_slice[1]), .SP(clk_c_enable_157), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i29.GSR = "DISABLED";
    FD1P3IX data_out__i28 (.D(data_out_slice[0]), .SP(clk_c_enable_157), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i28.GSR = "DISABLED";
    FD1P3IX data_out__i27 (.D(\data_out_slice[3] ), .SP(clk_c_enable_161), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i27.GSR = "DISABLED";
    FD1P3IX data_out__i26 (.D(data_out_slice[2]), .SP(clk_c_enable_161), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i26.GSR = "DISABLED";
    FD1P3IX data_out__i25 (.D(data_out_slice[1]), .SP(clk_c_enable_161), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i25.GSR = "DISABLED";
    FD1P3IX data_out__i24 (.D(data_out_slice[0]), .SP(clk_c_enable_161), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i24.GSR = "DISABLED";
    FD1P3IX data_out__i23 (.D(\data_out_slice[3] ), .SP(clk_c_enable_165), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[23])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i23.GSR = "DISABLED";
    FD1P3IX data_out__i22 (.D(data_out_slice[2]), .SP(clk_c_enable_165), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[22])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i22.GSR = "DISABLED";
    FD1P3IX data_out__i21 (.D(data_out_slice[1]), .SP(clk_c_enable_165), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[21])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i21.GSR = "DISABLED";
    FD1P3IX data_out__i20 (.D(data_out_slice[0]), .SP(clk_c_enable_165), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[20])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i20.GSR = "DISABLED";
    FD1P3IX data_out__i19 (.D(\data_out_slice[3] ), .SP(clk_c_enable_169), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[19])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i19.GSR = "DISABLED";
    FD1P3IX data_out__i18 (.D(data_out_slice[2]), .SP(clk_c_enable_169), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[18])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i18.GSR = "DISABLED";
    FD1P3IX data_out__i17 (.D(data_out_slice[1]), .SP(clk_c_enable_169), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[17])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i17.GSR = "DISABLED";
    FD1P3IX data_out__i16 (.D(data_out_slice[0]), .SP(clk_c_enable_169), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[16])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i16.GSR = "DISABLED";
    FD1P3IX data_out__i15 (.D(\data_out_slice[3] ), .SP(clk_c_enable_173), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i15.GSR = "DISABLED";
    FD1P3IX data_out__i14 (.D(data_out_slice[2]), .SP(clk_c_enable_173), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i14.GSR = "DISABLED";
    FD1P3IX data_out__i13 (.D(data_out_slice[1]), .SP(clk_c_enable_173), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i13.GSR = "DISABLED";
    FD1P3IX data_out__i12 (.D(data_out_slice[0]), .SP(clk_c_enable_173), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i12.GSR = "DISABLED";
    FD1P3IX data_out__i11 (.D(\data_out_slice[3] ), .SP(clk_c_enable_177), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i11.GSR = "DISABLED";
    FD1P3IX data_out__i10 (.D(data_out_slice[2]), .SP(clk_c_enable_177), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i10.GSR = "DISABLED";
    FD1P3IX data_out__i9 (.D(data_out_slice[1]), .SP(clk_c_enable_177), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i9.GSR = "DISABLED";
    FD1P3IX data_out__i8 (.D(data_out_slice[0]), .SP(clk_c_enable_177), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i8.GSR = "DISABLED";
    FD1P3IX data_out__i7 (.D(\data_out_slice[3] ), .SP(clk_c_enable_181), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i7.GSR = "DISABLED";
    FD1P3IX data_out__i6 (.D(data_out_slice[2]), .SP(clk_c_enable_181), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i6.GSR = "DISABLED";
    FD1P3IX data_out__i5 (.D(data_out_slice[1]), .SP(clk_c_enable_181), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i5.GSR = "DISABLED";
    FD1P3IX data_out__i4 (.D(data_out_slice[0]), .SP(clk_c_enable_181), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i4.GSR = "DISABLED";
    LUT4 i27881_3_lut_4_lut (.A(n26), .B(n31722), .C(n4271), .D(n4279), 
         .Z(n29428)) /* synthesis lut_function=(!(A (B (C+(D))))) */ ;
    defparam i27881_3_lut_4_lut.init = 16'h777f;
    FD1P3IX data_out__i3 (.D(\data_out_slice[3] ), .SP(clk_c_enable_184), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i3.GSR = "DISABLED";
    FD1P3IX data_out__i2 (.D(data_out_slice[2]), .SP(clk_c_enable_184), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i2.GSR = "DISABLED";
    FD1P3IX data_out__i1 (.D(data_out_slice[1]), .SP(clk_c_enable_184), 
            .CD(n31980), .CK(clk_c), .Q(data_to_write[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam data_out__i1.GSR = "DISABLED";
    LUT4 mux_2119_i14_3_lut_4_lut (.A(n26), .B(n31722), .C(n3381[11]), 
         .D(n5223[12]), .Z(n3422[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_2119_i14_3_lut_4_lut.init = 16'hf870;
    LUT4 data_from_read_9__bdd_3_lut_then_3_lut (.A(n31879), .B(n19), .C(n31885), 
         .Z(n32071)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam data_from_read_9__bdd_3_lut_then_3_lut.init = 16'hcece;
    LUT4 data_from_read_9__bdd_3_lut_else_3_lut (.A(n31879), .B(n19), .C(\peri_data_out[9] ), 
         .D(n4), .Z(n32070)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam data_from_read_9__bdd_3_lut_else_3_lut.init = 16'heeec;
    LUT4 n31958_bdd_3_lut (.A(counter_hi[2]), .B(\mem_data_from_read[20] ), 
         .C(\mem_data_from_read[16] ), .Z(n32183)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n31958_bdd_3_lut.init = 16'hd8d8;
    LUT4 i27591_3_lut_4_lut_4_lut (.A(n31719), .B(n26764), .C(n4277), 
         .D(n31865), .Z(n3381[7])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i27591_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_2119_i12_3_lut_4_lut (.A(n26), .B(n31722), .C(n3381[11]), 
         .D(n3271[11]), .Z(n3422[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_2119_i12_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_4_lut_then_4_lut (.A(n31813), .B(n2525[2]), .C(n27746), .D(n31852), 
         .Z(n32075)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h4010;
    LUT4 i1_4_lut_else_4_lut (.A(n31813), .B(n2505[2]), .C(n27746), .D(n31852), 
         .Z(n32074)) /* synthesis lut_function=(!(A+!(B (C (D))+!B !((D)+!C)))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h4010;
    LUT4 i27903_3_lut (.A(n4281), .B(n31732), .C(n31944), .Z(n29371)) /* synthesis lut_function=(A+!((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27903_3_lut.init = 16'haeae;
    LUT4 mux_1538_i16_3_lut_then_3_lut (.A(n21[15]), .B(n6[15]), .C(n2524), 
         .Z(n32079)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1538_i16_3_lut_then_3_lut.init = 16'hacac;
    PFUMX i28444 (.BLUT(n31416), .ALUT(n31415), .C0(n31770), .Z(n31417));
    LUT4 mux_1538_i16_3_lut_else_3_lut (.A(n27[15]), .B(n31[15]), .C(n2504), 
         .Z(n32078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1538_i16_3_lut_else_3_lut.init = 16'hcaca;
    LUT4 n32183_bdd_3_lut (.A(n32183), .B(n13), .C(n31958), .Z(n32184)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n32183_bdd_3_lut.init = 16'hcaca;
    LUT4 n29658_bdd_3_lut (.A(n29658), .B(n32184), .C(counter_hi[4]), 
         .Z(n32185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n29658_bdd_3_lut.init = 16'hcaca;
    FD1P3IX load_started_422 (.D(VCC_net), .SP(address_ready), .CD(n844), 
            .CK(clk_c), .Q(load_started)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam load_started_422.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(rst_reg_n), .B(clk_c_enable_30), .C(n43), 
         .D(n31838), .Z(n2134)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h8880;
    PFUMX i28613 (.BLUT(n32064), .ALUT(n32065), .C0(counter_hi[2]), .Z(n32066));
    LUT4 n31792_bdd_4_lut_29319 (.A(n31792), .B(data_txn_len[0]), .C(instr_data[10]), 
         .D(instr_data[2]), .Z(n32280)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam n31792_bdd_4_lut_29319.init = 16'hfd20;
    LUT4 i1_2_lut_rep_514_3_lut_4_lut (.A(rst_reg_n), .B(clk_c_enable_30), 
         .C(n22), .D(n31838), .Z(n31719)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_514_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(rst_reg_n), .B(clk_c_enable_30), .C(n35), 
         .D(n31838), .Z(n4277)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_697_3_lut_4_lut (.A(addr[27]), .B(n31997), .C(n18241), 
         .D(n32033), .Z(n31902)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_697_3_lut_4_lut.init = 16'h000e;
    LUT4 pc_1__bdd_3_lut_28084 (.A(\pc[5] ), .B(\pc[13] ), .C(counter_hi[3]), 
         .Z(n30803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_1__bdd_3_lut_28084.init = 16'hcaca;
    LUT4 n31417_bdd_3_lut_4_lut (.A(addr[27]), .B(n31997), .C(n32066), 
         .D(n31417), .Z(n31418)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n31417_bdd_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i28436 (.BLUT(n31406), .ALUT(n31405), .C0(n31770), .Z(n31407));
    LUT4 mux_2119_i13_3_lut_4_lut (.A(n26), .B(n31722), .C(n3381[11]), 
         .D(n5223[11]), .Z(n3422[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_2119_i13_3_lut_4_lut.init = 16'hf870;
    LUT4 data_from_read_2__bdd_4_lut_29318 (.A(n28964), .B(n31879), .C(n10467), 
         .D(\peri_data_out[6] ), .Z(n32277)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam data_from_read_2__bdd_4_lut_29318.init = 16'hfefa;
    PFUMX i28051 (.BLUT(n30748), .ALUT(n30747), .C0(counter_hi[2]), .Z(n30749));
    LUT4 i27945_3_lut_4_lut (.A(addr[27]), .B(n31997), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n29318)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i27945_3_lut_4_lut.init = 16'hefff;
    LUT4 i43_3_lut (.A(n31860), .B(n31867), .C(n26119), .Z(n24)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;
    defparam i43_3_lut.init = 16'h6464;
    LUT4 i1_4_lut (.A(n22_adj_3135), .B(n9894), .C(n4_adj_3136), .D(n31791), 
         .Z(n28140)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0002;
    FD1P3IX is_jal_401 (.D(is_jal_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_jal)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_jal_401.GSR = "DISABLED";
    FD1P3AX imm_i0_i31 (.D(n3546[31]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(imm[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i31.GSR = "DISABLED";
    LUT4 n31425_bdd_3_lut_4_lut (.A(addr[27]), .B(n31997), .C(n32063), 
         .D(n31425), .Z(n29759)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n31425_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1538_i3_3_lut (.A(n29063), .B(n2163[2]), .C(n31944), .Z(instr[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1538_i3_3_lut.init = 16'hcaca;
    LUT4 n31310_bdd_3_lut_4_lut (.A(addr[27]), .B(n31997), .C(n13), .D(n31310), 
         .Z(n31311)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n31310_bdd_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX imm_i0_i30 (.D(n30762), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(imm[30])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i30.GSR = "DISABLED";
    FD1P3AX imm_i0_i29 (.D(n3546[29]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(imm[29])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i29.GSR = "DISABLED";
    FD1P3AX imm_i0_i28 (.D(n3546[28]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(imm[28])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i28.GSR = "DISABLED";
    FD1P3AX imm_i0_i27 (.D(n3546[27]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(imm[27])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i27.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_398 (.A(addr[27]), .B(n31997), .C(\addr[7] ), 
         .D(n4_adj_11), .Z(n26216)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_3_lut_4_lut_adj_398.init = 16'h00e0;
    LUT4 n31683_bdd_3_lut (.A(instr[17]), .B(instr[31]), .C(n4263), .Z(n31684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31683_bdd_3_lut.init = 16'hcaca;
    LUT4 n17863_bdd_3_lut_28598 (.A(n2143[1]), .B(n2163[1]), .C(n31944), 
         .Z(instr[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n17863_bdd_3_lut_28598.init = 16'hcaca;
    FD1P3AX imm_i0_i26 (.D(n3546[26]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(imm[26])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i26.GSR = "DISABLED";
    LUT4 mux_2147_i32_4_lut (.A(n3505[17]), .B(instr[31]), .C(n4285), 
         .D(n10068), .Z(n3546[31])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i32_4_lut.init = 16'hca0a;
    FD1P3AX imm_i0_i25 (.D(n3546[25]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(imm[25])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i25.GSR = "DISABLED";
    LUT4 n31315_bdd_3_lut_4_lut (.A(addr[27]), .B(n31997), .C(n13), .D(n31315), 
         .Z(n31316)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n31315_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_rep_535 (.A(address_ready), .B(n31743), .C(is_load), 
         .Z(n31740)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(291[13:39])
    defparam i1_3_lut_rep_535.init = 16'h2020;
    LUT4 pc_1__bdd_3_lut_28560 (.A(\pc[1] ), .B(\pc[9] ), .C(counter_hi[3]), 
         .Z(n30804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_1__bdd_3_lut_28560.init = 16'hcaca;
    LUT4 n31407_bdd_3_lut_4_lut (.A(addr[27]), .B(n31997), .C(n32072), 
         .D(n31407), .Z(n31408)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam n31407_bdd_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX imm_i0_i24 (.D(n3546[24]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(imm[24])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i24.GSR = "DISABLED";
    FD1S3IX counter_hi_3563__i2 (.D(c_2__N_1861[0]), .CK(clk_c), .CD(n31980), 
            .Q(counter_hi[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3563__i2.GSR = "DISABLED";
    FD1P3AX imm_i0_i23 (.D(n3546[23]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[23] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i23.GSR = "DISABLED";
    FD1P3AX imm_i0_i22 (.D(n3546[22]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[22] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i22.GSR = "DISABLED";
    FD1P3AX imm_i0_i21 (.D(n3546[21]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[21] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i21.GSR = "DISABLED";
    FD1P3AX imm_i0_i20 (.D(n3546[20]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[20] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i20.GSR = "DISABLED";
    FD1P3AX imm_i0_i19 (.D(n30767), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[19] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i19.GSR = "DISABLED";
    FD1P3AX imm_i0_i18 (.D(n30775), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[18] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i18.GSR = "DISABLED";
    FD1P3AX imm_i0_i17 (.D(n31687), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[17] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i17.GSR = "DISABLED";
    FD1S3IX addr_offset_3564__i2 (.D(n33[0]), .CK(clk_c), .CD(n31980), 
            .Q(addr_offset[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam addr_offset_3564__i2.GSR = "DISABLED";
    FD1P3AX imm_i0_i16 (.D(n3546[16]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[16] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i16.GSR = "DISABLED";
    FD1P3AX imm_i0_i15 (.D(n3546[15]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[15] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i15.GSR = "DISABLED";
    FD1P3AX imm_i0_i14 (.D(n3546[14]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[14] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i14.GSR = "DISABLED";
    FD1P3AX imm_i0_i13 (.D(n3546[13]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[13] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i13.GSR = "DISABLED";
    FD1P3AX imm_i0_i12 (.D(n3546[12]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[12] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i12.GSR = "DISABLED";
    FD1P3AX imm_i0_i11 (.D(n3546[11]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[11] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i11.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(address_ready), .B(n31743), .C(is_load), .D(n31884), 
         .Z(clk_c_enable_108)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(291[13:39])
    defparam i1_2_lut_4_lut.init = 16'hff20;
    LUT4 n3520_bdd_3_lut (.A(n3505[17]), .B(n31686), .C(n4285), .Z(n31687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3520_bdd_3_lut.init = 16'hcaca;
    FD1P3AX imm_i0_i10 (.D(n3546[10]), .SP(clk_c_enable_212), .CK(clk_c), 
            .Q(\imm[10] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i10.GSR = "DISABLED";
    FD1P3AX imm_i0_i9 (.D(n30840), .SP(clk_c_enable_214), .CK(clk_c), 
            .Q(\imm[9] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i9.GSR = "DISABLED";
    FD1P3AX imm_i0_i8 (.D(n3546[8]), .SP(clk_c_enable_214), .CK(clk_c), 
            .Q(\imm[8] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i8.GSR = "DISABLED";
    FD1P3AX imm_i0_i7 (.D(n3546[7]), .SP(clk_c_enable_221), .CK(clk_c), 
            .Q(\imm[7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i7.GSR = "DISABLED";
    FD1P3AX imm_i0_i6 (.D(n3546[6]), .SP(clk_c_enable_221), .CK(clk_c), 
            .Q(\imm[6] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i6.GSR = "DISABLED";
    FD1P3AX imm_i0_i5 (.D(n3546[5]), .SP(clk_c_enable_221), .CK(clk_c), 
            .Q(\imm[5] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i5.GSR = "DISABLED";
    FD1P3AX imm_i0_i4 (.D(n3546[4]), .SP(clk_c_enable_221), .CK(clk_c), 
            .Q(\imm[4] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i4.GSR = "DISABLED";
    FD1P3AX imm_i0_i3 (.D(n3546[3]), .SP(clk_c_enable_221), .CK(clk_c), 
            .Q(\imm[3] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i3.GSR = "DISABLED";
    FD1P3AX imm_i0_i2 (.D(n30709), .SP(clk_c_enable_221), .CK(clk_c), 
            .Q(\imm[2] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i2.GSR = "DISABLED";
    FD1P3AX imm_i0_i1 (.D(n3546[1]), .SP(clk_c_enable_221), .CK(clk_c), 
            .Q(\imm[1] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam imm_i0_i1.GSR = "DISABLED";
    LUT4 mux_1822_i1_3_lut (.A(n21[0]), .B(n27[0]), .C(n2504), .Z(n2505[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1532_i14_3_lut (.A(n6[13]), .B(n21[13]), .C(n2524), .Z(n2163[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i14_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_399 (.A(n27018), .B(n31743), .C(n27846), 
         .D(n31748), .Z(n26948)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[22:78])
    defparam i1_2_lut_3_lut_4_lut_adj_399.init = 16'h0f0d;
    LUT4 i1_2_lut_3_lut (.A(n27018), .B(n31743), .C(n28150), .Z(n28152)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[22:78])
    defparam i1_2_lut_3_lut.init = 16'hd0d0;
    LUT4 mux_1528_i14_3_lut (.A(n27[13]), .B(n31[13]), .C(n2504), .Z(n2143[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1826_i1_3_lut (.A(n31[0]), .B(n6[0]), .C(n2524), .Z(n2525[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1532_i13_3_lut (.A(n6[12]), .B(n21[12]), .C(n2524), .Z(n2163[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i13_3_lut.init = 16'hcaca;
    LUT4 mux_1528_i13_3_lut (.A(n27[12]), .B(n31[12]), .C(n2504), .Z(n2143[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i13_3_lut.init = 16'hcaca;
    LUT4 n30805_bdd_3_lut (.A(n30805), .B(n30802), .C(n33484), .Z(debug_branch_N_442[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30805_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_1532_i12_3_lut (.A(n6[11]), .B(n21[11]), .C(n2524), .Z(n2163[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1528_i12_3_lut (.A(n27[11]), .B(n31[11]), .C(n2504), .Z(n2143[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i12_3_lut.init = 16'hcaca;
    LUT4 mux_1532_i10_3_lut (.A(n6[9]), .B(n21[9]), .C(n2524), .Z(n2163[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1528_i10_3_lut (.A(n27[9]), .B(n31[9]), .C(n2504), .Z(n2143[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1532_i9_3_lut (.A(n6[8]), .B(n21[8]), .C(n2524), .Z(n2163[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i9_3_lut.init = 16'hcaca;
    LUT4 mux_1528_i9_3_lut (.A(n27[8]), .B(n31[8]), .C(n2504), .Z(n2143[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_400 (.A(n27018), .B(n31743), .C(n33488), .Z(n27460)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[22:78])
    defparam i1_2_lut_3_lut_adj_400.init = 16'hd0d0;
    LUT4 mux_1532_i4_3_lut (.A(n6[3]), .B(n21[3]), .C(n2524), .Z(n2163[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1528_i4_3_lut (.A(n27[3]), .B(n31[3]), .C(n2504), .Z(n2143[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i4_3_lut.init = 16'hcaca;
    LUT4 mux_2147_i30_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n5121[29]), .Z(n3546[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i30_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_2_lut_rep_529_3_lut_4_lut (.A(n27018), .B(n31743), .C(n27846), 
         .D(n31748), .Z(n31734)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[22:78])
    defparam i1_2_lut_rep_529_3_lut_4_lut.init = 16'hf0f2;
    FD1P3AX data_write_n_i0 (.D(data_write_n_1__N_369[0]), .SP(clk_c_enable_224), 
            .CK(clk_c), .Q(qv_data_write_n[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam data_write_n_i0.GSR = "DISABLED";
    FD1P3IX is_alu_reg_397 (.D(is_alu_reg_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_alu_reg)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_alu_reg_397.GSR = "DISABLED";
    PFUMX i28047 (.BLUT(n30743), .ALUT(n30742), .C0(counter_hi[2]), .Z(n30744));
    LUT4 mux_2147_i26_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n5121[25]), .Z(n3546[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i26_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_3_lut_4_lut_adj_401 (.A(n10499), .B(n31730), .C(data_txn_len[1]), 
         .D(instr_active), .Z(\txn_len[1] )) /* synthesis lut_function=(!(A ((D)+!C)+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(435[34:115])
    defparam i1_3_lut_4_lut_adj_401.init = 16'h00b0;
    LUT4 mux_2147_i29_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n5121[28]), .Z(n3546[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i29_3_lut_4_lut.init = 16'hf870;
    LUT4 i5725_4_lut_4_lut (.A(clk_c_enable_30), .B(n31796), .C(additional_mem_ops[0]), 
         .D(n31846), .Z(additional_mem_ops_de[0])) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i5725_4_lut_4_lut.init = 16'hd850;
    FD1P3AX instr_data_3__i64 (.D(instr_data[15]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i64.GSR = "DISABLED";
    LUT4 mux_1822_i16_3_lut (.A(n21[15]), .B(n27[15]), .C(n2504), .Z(n2505[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i16_3_lut.init = 16'hcaca;
    LUT4 mux_2147_i28_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n5121[27]), .Z(n3546[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i28_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_2_lut_rep_695_3_lut_4_lut (.A(\addr[5] ), .B(n32035), .C(n32019), 
         .D(\addr[4] ), .Z(n31900)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_695_3_lut_4_lut.init = 16'hfdff;
    LUT4 i1_4_lut_4_lut (.A(n31845), .B(n24), .C(n28006), .D(n28332), 
         .Z(n27862)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_4_lut.init = 16'hf040;
    LUT4 i1_2_lut_rep_696_3_lut_4_lut (.A(\addr[5] ), .B(n32035), .C(n26266), 
         .D(\addr[4] ), .Z(n31901)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_696_3_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_402 (.A(\addr[5] ), .B(n32035), .C(n32019), 
         .D(\addr[4] ), .Z(n80)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_4_lut_adj_402.init = 16'hfffd;
    LUT4 i46_3_lut_4_lut_3_lut (.A(n31845), .B(n31868), .C(n31867), .Z(n41)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;
    defparam i46_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 mux_2147_i25_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n5121[24]), .Z(n3546[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i25_3_lut_4_lut.init = 16'hf870;
    FD1P3AX instr_data_3__i63 (.D(instr_data[14]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i63.GSR = "DISABLED";
    LUT4 mux_2096_i6_4_lut_4_lut (.A(n31845), .B(n4271), .C(n31868), .D(n31846), 
         .Z(n3271[5])) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C+(D))+!B (D))) */ ;
    defparam mux_2096_i6_4_lut_4_lut.init = 16'hddc0;
    LUT4 mux_2096_i2_4_lut_4_lut (.A(n31845), .B(n4271), .C(n31868), .D(n31852), 
         .Z(n3271[1])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_2096_i2_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_29_i3_3_lut_4_lut_4_lut (.A(n31845), .B(n155[2]), .C(n31813), 
         .D(n31820), .Z(alu_op_3__N_1170[2])) /* synthesis lut_function=(A (B (C+(D)))+!A (B+!(C+(D)))) */ ;
    defparam mux_29_i3_3_lut_4_lut_4_lut.init = 16'hccc5;
    LUT4 n31194_bdd_4_lut_4_lut (.A(n31845), .B(n31860), .C(n31867), .D(n31868), 
         .Z(n31439)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam n31194_bdd_4_lut_4_lut.init = 16'h0040;
    LUT4 i4589_3_lut_4_lut (.A(\instr_addr_23__N_318[0] ), .B(n32042), .C(n31978), 
         .D(instr_addr_23__N_318[1]), .Z(n4_adj_3138)) /* synthesis lut_function=(A ((D)+!C)+!A !(B (C+!(D))+!B !((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i4589_3_lut_4_lut.init = 16'hbf0b;
    LUT4 mux_2096_i4_4_lut_4_lut (.A(n31845), .B(n4271), .C(n31868), .D(n31851), 
         .Z(n3271[3])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_2096_i4_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i1_4_lut_4_lut_adj_403 (.A(\instr_write_offset[3] ), .B(instr_addr_23__N_318[1]), 
         .C(\pc[2] ), .D(n28260), .Z(n9_c)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A !(B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam i1_4_lut_4_lut_adj_403.init = 16'h4124;
    LUT4 mux_2096_i3_4_lut_4_lut (.A(n31845), .B(n4271), .C(n31868), .D(n31847), 
         .Z(n3271[2])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam mux_2096_i3_4_lut_4_lut.init = 16'hd1c0;
    LUT4 n4271_bdd_4_lut_28549 (.A(n31719), .B(n4277), .C(n26770), .D(n27726), 
         .Z(n30838)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam n4271_bdd_4_lut_28549.init = 16'hd1c0;
    LUT4 i1_4_lut_adj_404 (.A(n31866), .B(next_instr_write_offset[3]), .C(n1), 
         .D(n27702), .Z(n13146)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_404.init = 16'h0400;
    LUT4 n30839_bdd_3_lut (.A(n30839), .B(n30835), .C(n4285), .Z(n30840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30839_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_2123_i21_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n29023), .Z(n3458[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2123_i21_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_1826_i16_3_lut (.A(n31[15]), .B(n6[15]), .C(n2524), .Z(n2525[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i16_3_lut.init = 16'hcaca;
    FD1P3IX is_jalr_400 (.D(is_jalr_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_jalr)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_jalr_400.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_405 (.A(n31851), .B(rst_reg_n), .C(n31867), 
         .Z(n27832)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_405.init = 16'h0808;
    LUT4 mux_1822_i14_3_lut (.A(n21[13]), .B(n27[13]), .C(n2504), .Z(n2505[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i14_3_lut.init = 16'hcaca;
    LUT4 mux_1826_i14_3_lut (.A(n31[13]), .B(n6[13]), .C(n2524), .Z(n2525[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i14_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_406 (.A(n7103), .B(n27604), .C(\instr_write_offset[3] ), 
         .D(instr_complete_N_1647), .Z(next_instr_write_offset[3])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i1_4_lut_adj_406.init = 16'h965a;
    LUT4 mux_2123_i22_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n29025), .Z(n3458[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2123_i22_3_lut_4_lut.init = 16'hf870;
    LUT4 i15832_2_lut_3_lut_4_lut (.A(n31845), .B(n31867), .C(n31847), 
         .D(n31822), .Z(n15_adj_3139)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15832_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3IX is_branch_399 (.D(is_branch_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_branch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_branch_399.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_525_4_lut (.A(n31747), .B(instr_fetch_running), .C(n27286), 
         .D(debug_ret), .Z(n31730)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_3_lut_rep_525_4_lut.init = 16'h0002;
    PFUMX i28387 (.BLUT(n31318), .ALUT(n31316), .C0(counter_hi[4]), .Z(n31319));
    LUT4 mux_2123_i23_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n29033), .Z(n3458[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2123_i23_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_2123_i24_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n2152), .Z(n3458[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2123_i24_3_lut_4_lut.init = 16'hf870;
    LUT4 i1_4_lut_adj_407 (.A(n31744), .B(n31738), .C(n31742), .D(n27750), 
         .Z(n4281)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_407.init = 16'h0400;
    LUT4 mux_2123_i27_3_lut_4_lut (.A(n4285), .B(n4281), .C(n5121[21]), 
         .D(n29051), .Z(n3458[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2123_i27_3_lut_4_lut.init = 16'hf870;
    LUT4 instr_addr_23__I_0_i2_3_lut (.A(instr_addr_23__N_318[1]), .B(\early_branch_addr[2] ), 
         .C(was_early_branch), .Z(\instr_addr[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(438[25:119])
    defparam instr_addr_23__I_0_i2_3_lut.init = 16'hcaca;
    FD1P3AX instr_data_3__i62 (.D(instr_data[13]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i62.GSR = "DISABLED";
    LUT4 i1_3_lut_3_lut_4_lut (.A(n22), .B(n31722), .C(n31863), .D(rst_reg_n), 
         .Z(n26693)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam i1_3_lut_3_lut_4_lut.init = 16'h7000;
    LUT4 i31_4_lut_4_lut (.A(n31845), .B(n31868), .C(n26119), .D(n31867), 
         .Z(n25)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam i31_4_lut_4_lut.init = 16'h11fa;
    FD1P3AX instr_data_3__i61 (.D(instr_data[12]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i61.GSR = "DISABLED";
    FD1P3AX instr_data_3__i60 (.D(instr_data[11]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i60.GSR = "DISABLED";
    FD1P3AX instr_data_3__i59 (.D(instr_data[10]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i59.GSR = "DISABLED";
    FD1P3AX instr_data_3__i58 (.D(instr_data[9]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i58.GSR = "DISABLED";
    FD1P3AX instr_data_3__i57 (.D(instr_data[8]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i57.GSR = "DISABLED";
    FD1P3AX instr_data_3__i56 (.D(instr_data[7]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[7])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i56.GSR = "DISABLED";
    FD1P3AX instr_data_3__i55 (.D(instr_data[6]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i55.GSR = "DISABLED";
    FD1P3AX instr_data_3__i54 (.D(instr_data[5]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i54.GSR = "DISABLED";
    FD1P3AX instr_data_3__i53 (.D(instr_data[4]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i53.GSR = "DISABLED";
    FD1P3AX instr_data_3__i52 (.D(instr_data[3]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i52.GSR = "DISABLED";
    FD1P3AX instr_data_3__i51 (.D(instr_data[2]), .SP(clk_c_enable_287), 
            .CK(clk_c), .Q(n21[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i51.GSR = "DISABLED";
    FD1P3AX instr_data_3__i50 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_289), 
            .CK(clk_c), .Q(n21[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i50.GSR = "DISABLED";
    FD1P3AX instr_data_3__i49 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_289), 
            .CK(clk_c), .Q(n21[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i49.GSR = "DISABLED";
    FD1P3AX instr_data_3__i48 (.D(instr_data[15]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i48.GSR = "DISABLED";
    FD1P3AX instr_data_3__i47 (.D(instr_data[14]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i47.GSR = "DISABLED";
    FD1P3AX instr_data_3__i46 (.D(instr_data[13]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i46.GSR = "DISABLED";
    FD1P3AX instr_data_3__i45 (.D(instr_data[12]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i45.GSR = "DISABLED";
    FD1P3AX instr_data_3__i44 (.D(instr_data[11]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i44.GSR = "DISABLED";
    FD1P3AX instr_data_3__i43 (.D(instr_data[10]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i43.GSR = "DISABLED";
    FD1P3AX instr_data_3__i42 (.D(instr_data[9]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i42.GSR = "DISABLED";
    FD1P3AX instr_data_3__i41 (.D(instr_data[8]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i41.GSR = "DISABLED";
    FD1P3AX instr_data_3__i40 (.D(instr_data[7]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(\instr_data[1][7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i40.GSR = "DISABLED";
    FD1P3AX instr_data_3__i39 (.D(instr_data[6]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i39.GSR = "DISABLED";
    FD1P3AX instr_data_3__i38 (.D(instr_data[5]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i38.GSR = "DISABLED";
    FD1P3AX instr_data_3__i37 (.D(instr_data[4]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i37.GSR = "DISABLED";
    FD1P3AX instr_data_3__i36 (.D(instr_data[3]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i36.GSR = "DISABLED";
    FD1P3AX instr_data_3__i35 (.D(instr_data[2]), .SP(clk_c_enable_303), 
            .CK(clk_c), .Q(n27[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i35.GSR = "DISABLED";
    FD1P3AX instr_data_3__i34 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_305), 
            .CK(clk_c), .Q(n27[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i34.GSR = "DISABLED";
    FD1P3AX instr_data_3__i33 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_305), 
            .CK(clk_c), .Q(n27[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i33.GSR = "DISABLED";
    FD1P3AX instr_data_3__i32 (.D(instr_data[15]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i32.GSR = "DISABLED";
    FD1P3AX instr_data_3__i31 (.D(instr_data[14]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i31.GSR = "DISABLED";
    FD1P3AX instr_data_3__i30 (.D(instr_data[13]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i30.GSR = "DISABLED";
    FD1P3AX instr_data_3__i29 (.D(instr_data[12]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i29.GSR = "DISABLED";
    FD1P3AX instr_data_3__i28 (.D(instr_data[11]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i28.GSR = "DISABLED";
    FD1P3AX instr_data_3__i27 (.D(instr_data[10]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i27.GSR = "DISABLED";
    FD1P3AX instr_data_3__i26 (.D(instr_data[9]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i26.GSR = "DISABLED";
    FD1P3AX instr_data_3__i25 (.D(instr_data[8]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i25.GSR = "DISABLED";
    FD1P3AX instr_data_3__i24 (.D(instr_data[7]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(\instr_data[2][7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i24.GSR = "DISABLED";
    FD1P3AX instr_data_3__i23 (.D(instr_data[6]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i23.GSR = "DISABLED";
    FD1P3AX instr_data_3__i22 (.D(instr_data[5]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i22.GSR = "DISABLED";
    FD1P3AX instr_data_3__i21 (.D(instr_data[4]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i21.GSR = "DISABLED";
    FD1P3AX instr_data_3__i20 (.D(instr_data[3]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i20.GSR = "DISABLED";
    FD1P3AX instr_data_3__i19 (.D(instr_data[2]), .SP(clk_c_enable_319), 
            .CK(clk_c), .Q(n31[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i19.GSR = "DISABLED";
    FD1P3AX instr_data_3__i18 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(n31[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i18.GSR = "DISABLED";
    FD1P3AX instr_data_3__i17 (.D(instr_data_0__15__N_638[0]), .SP(clk_c_enable_321), 
            .CK(clk_c), .Q(n31[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i17.GSR = "DISABLED";
    FD1P3AX instr_data_3__i16 (.D(instr_data[15]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[15])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i16.GSR = "DISABLED";
    FD1P3AX instr_data_3__i15 (.D(instr_data[14]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[14])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i15.GSR = "DISABLED";
    FD1P3AX mem_op_increment_reg_413 (.D(mem_op_increment_reg_de), .SP(clk_c_enable_325), 
            .CK(clk_c), .Q(mem_op_increment_reg)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam mem_op_increment_reg_413.GSR = "DISABLED";
    LUT4 i1_3_lut_3_lut_4_lut_adj_408 (.A(n31845), .B(n31868), .C(n33488), 
         .D(n31838), .Z(n27942)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_3_lut_4_lut_adj_408.init = 16'h0010;
    LUT4 i15374_2_lut_3_lut_4_lut (.A(n22), .B(n31722), .C(n31853), .D(n31720), 
         .Z(n3195[5])) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (C)) */ ;
    defparam i15374_2_lut_3_lut_4_lut.init = 16'hf070;
    LUT4 i52_4_lut_4_lut (.A(n31869), .B(n31867), .C(n17976), .D(n31845), 
         .Z(n37)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B (D)+!B !(C+(D))))) */ ;
    defparam i52_4_lut_4_lut.init = 16'h4403;
    LUT4 mux_1822_i13_3_lut (.A(n21[12]), .B(n27[12]), .C(n2504), .Z(n2505[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i13_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_409 (.A(n31847), .B(n33488), .C(n31867), .Z(n27818)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_409.init = 16'h0808;
    LUT4 i1_2_lut_rep_572_3_lut (.A(n31869), .B(n31867), .C(n31860), .Z(n31777)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_572_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_555_3_lut_4_lut (.A(n31869), .B(n31867), .C(n31845), 
         .D(n31860), .Z(n31760)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_555_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_4_lut_4_lut_4_lut (.A(n31869), .B(n31867), .C(n31868), 
         .D(n31845), .Z(n24_adj_3140)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A (B (C (D))+!B (C+(D)))) */ ;
    defparam i1_4_lut_4_lut_4_lut_4_lut.init = 16'hf130;
    FD1P3AX instr_data_3__i14 (.D(instr_data[13]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[13])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i14.GSR = "DISABLED";
    LUT4 i15995_2_lut_3_lut_4_lut (.A(n31869), .B(n31867), .C(n31868), 
         .D(n31845), .Z(n30)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i15995_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_410 (.A(debug_ret), .B(n27286), .C(debug_stop_txn_N_2148), 
         .D(n31745), .Z(debug_stop_txn_N_2147)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_410.init = 16'h1000;
    FD1P3AX instr_data_3__i13 (.D(instr_data[12]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[12])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i13.GSR = "DISABLED";
    FD1P3AX instr_data_3__i12 (.D(instr_data[11]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[11])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i12.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(instr_fetch_running_N_945), .B(n13146), .Z(debug_stop_txn_N_2148)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i1_2_lut.init = 16'hdddd;
    FD1P3AX instr_data_3__i11 (.D(instr_data[10]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[10])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i11.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_411 (.A(qspi_data_ready), .B(n27606), .C(n32052), 
         .D(next_instr_write_offset[3]), .Z(n58)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_4_lut_adj_411.init = 16'hc4f5;
    LUT4 i1_4_lut_adj_412 (.A(was_early_branch), .B(n10112), .C(n16), 
         .D(n31838), .Z(n9894)) /* synthesis lut_function=(A+(B (C (D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[82:120])
    defparam i1_4_lut_adj_412.init = 16'hfaba;
    LUT4 n4271_bdd_3_lut_4_lut (.A(n31849), .B(n31845), .C(n2982[13]), 
         .D(n4271), .Z(n30836)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam n4271_bdd_3_lut_4_lut.init = 16'hf022;
    FD1P3AX instr_data_3__i10 (.D(instr_data[9]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[9])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i10.GSR = "DISABLED";
    LUT4 i15859_2_lut_rep_573_3_lut (.A(n31860), .B(n31845), .C(n31853), 
         .Z(n31778)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15859_2_lut_rep_573_3_lut.init = 16'h4040;
    FD1P3AX instr_data_3__i9 (.D(instr_data[8]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[8])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i9.GSR = "DISABLED";
    FD1P3AX instr_data_3__i8 (.D(instr_data[7]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(\instr_data[3][7] )) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i8.GSR = "DISABLED";
    FD1P3AX instr_data_3__i7 (.D(instr_data[6]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[6])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i7.GSR = "DISABLED";
    FD1P3AX instr_data_3__i6 (.D(instr_data[5]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[5])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i6.GSR = "DISABLED";
    FD1P3AX instr_data_3__i5 (.D(instr_data[4]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[4])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i5.GSR = "DISABLED";
    FD1P3AX instr_data_3__i4 (.D(instr_data[3]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i4.GSR = "DISABLED";
    FD1P3AX instr_data_3__i3 (.D(instr_data[2]), .SP(clk_c_enable_342), 
            .CK(clk_c), .Q(n6[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i3.GSR = "DISABLED";
    FD1P3AX instr_data_3__i2 (.D(instr_data_0__15__N_638[49]), .SP(clk_c_enable_343), 
            .CK(clk_c), .Q(n6[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_data_3__i2.GSR = "DISABLED";
    LUT4 i15858_2_lut_3_lut (.A(n31860), .B(n31845), .C(n31852), .Z(n3304[1])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15858_2_lut_3_lut.init = 16'h4040;
    LUT4 mux_2096_i12_4_lut_4_lut_4_lut (.A(n31860), .B(n31845), .C(n4279), 
         .D(n31853), .Z(n3271[11])) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (C (D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2096_i12_4_lut_4_lut_4_lut.init = 16'h4300;
    LUT4 i1_4_lut_adj_413 (.A(n28284), .B(n27056), .C(n31965), .D(n32055), 
         .Z(n12_c)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !((C (D)+!C !(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(224[82:120])
    defparam i1_4_lut_adj_413.init = 16'h8448;
    LUT4 i1_4_lut_adj_414 (.A(n19_adj_3141), .B(n28018), .C(n31818), .D(n31772), 
         .Z(n28020)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A ((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_414.init = 16'h0c88;
    LUT4 i1_4_lut_adj_415 (.A(n9894), .B(n31774), .C(n31831), .D(rst_reg_n), 
         .Z(n28018)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_415.init = 16'h0400;
    LUT4 stall_core_I_0_438_2_lut_rep_767 (.A(stall_core), .B(interrupt_core), 
         .Z(n31972)) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(340[19:48])
    defparam stall_core_I_0_438_2_lut_rep_767.init = 16'h1111;
    L6MUX21 i28034 (.D0(n30708), .D1(n3458[2]), .SD(n4285), .Z(n30709));
    FD1P3IX alu_op__i3 (.D(alu_op_de[3]), .SP(clk_c_enable_347), .CD(n31980), 
            .CK(clk_c), .Q(alu_op[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i3.GSR = "DISABLED";
    FD1P3IX alu_op__i2 (.D(alu_op_de[2]), .SP(clk_c_enable_347), .CD(n31980), 
            .CK(clk_c), .Q(alu_op_in[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i2.GSR = "DISABLED";
    FD1P3IX alu_op__i1 (.D(alu_op_de[1]), .SP(clk_c_enable_347), .CD(n31980), 
            .CK(clk_c), .Q(alu_op[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam alu_op__i1.GSR = "DISABLED";
    LUT4 i15756_2_lut_3_lut (.A(stall_core), .B(interrupt_core), .C(n32029), 
         .Z(n18324)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(340[19:48])
    defparam i15756_2_lut_3_lut.init = 16'h1f1f;
    LUT4 i1_2_lut_rep_683_3_lut_4_lut_4_lut (.A(stall_core), .B(interrupt_core), 
         .C(n26175), .D(n32044), .Z(n31888)) /* synthesis lut_function=((B+!((D)+!C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(340[19:48])
    defparam i1_2_lut_rep_683_3_lut_4_lut_4_lut.init = 16'hddfd;
    LUT4 i1_4_lut_adj_416 (.A(clk_c_enable_448), .B(n31742), .C(n27796), 
         .D(n31738), .Z(n2500)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_416.init = 16'ha888;
    FD1P3IX is_system_402 (.D(is_system_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_system)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_system_402.GSR = "DISABLED";
    FD1P3IX is_lui_398 (.D(is_lui_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_lui)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_lui_398.GSR = "DISABLED";
    LUT4 i3_2_lut_3_lut_3_lut_4_lut (.A(n31869), .B(n31868), .C(n31867), 
         .D(n31845), .Z(n17)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_2_lut_3_lut_3_lut_4_lut.init = 16'h0010;
    FD1P3IX is_auipc_395 (.D(is_auipc_de), .SP(clk_c_enable_358), .CD(n31980), 
            .CK(clk_c), .Q(is_auipc)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam is_auipc_395.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_417 (.A(debug_ret), .B(n27286), .C(n31747), .D(n28912), 
         .Z(start_instr)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_417.init = 16'h0010;
    FD1P3AX instr_fetch_running_429 (.D(n6411), .SP(clk_c_enable_370), .CK(clk_c), 
            .Q(instr_fetch_running)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam instr_fetch_running_429.GSR = "DISABLED";
    FD1P3AX data_ready_latch_416 (.D(n27110), .SP(clk_c_enable_375), .CK(clk_c), 
            .Q(data_ready_latch)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(235[12] 256[8])
    defparam data_ready_latch_416.GSR = "DISABLED";
    LUT4 i26980_3_lut (.A(imm[27]), .B(imm[31]), .C(counter_hi[2]), .Z(n29597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26980_3_lut.init = 16'hcaca;
    PFUMX i28032 (.BLUT(n30707), .ALUT(n30706), .C0(n31718), .Z(n30708));
    LUT4 i26354_2_lut (.A(n10499), .B(instr_fetch_running), .Z(n28912)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26354_2_lut.init = 16'heeee;
    LUT4 i26979_3_lut (.A(\imm[19] ), .B(\imm[23] ), .C(counter_hi[2]), 
         .Z(n29596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26979_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_418 (.A(n31741), .B(n8), .C(n31748), .D(n31754), 
         .Z(debug_ret)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_418.init = 16'h0200;
    LUT4 i1_4_lut_adj_419 (.A(n31748), .B(n27460), .C(is_jal_de), .D(n8), 
         .Z(n27286)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_419.init = 16'h0040;
    LUT4 next_pc_for_core_23__I_0_i270_4_lut (.A(n5677[1]), .B(debug_rd_3__N_405[29]), 
         .C(n32001), .D(n9033), .Z(debug_branch_N_446[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i270_4_lut.init = 16'hcac0;
    LUT4 i26308_4_lut (.A(n31777), .B(n31848), .C(n31868), .D(n31845), 
         .Z(n28864)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i26308_4_lut.init = 16'hfaea;
    LUT4 next_pc_for_core_23__I_0_i271_4_lut (.A(n5677[2]), .B(debug_rd_3__N_405[30]), 
         .C(n32001), .D(n9033), .Z(debug_branch_N_446[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i271_4_lut.init = 16'hcac0;
    LUT4 next_pc_for_core_23__I_0_i272_4_lut (.A(n5677[3]), .B(\debug_rd_3__N_405[31] ), 
         .C(n32001), .D(n9033), .Z(debug_branch_N_446[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i272_4_lut.init = 16'hcac0;
    LUT4 i26978_3_lut (.A(\imm[11] ), .B(\imm[15] ), .C(counter_hi[2]), 
         .Z(n29595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26978_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_420 (.A(n27480), .B(n31742), .C(n9894), .D(instr_complete_N_1647), 
         .Z(n8)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_420.init = 16'hfefc;
    LUT4 i26977_3_lut (.A(\imm[3] ), .B(\imm[7] ), .C(counter_hi[2]), 
         .Z(n29594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26977_3_lut.init = 16'hcaca;
    LUT4 i26530_3_lut_4_lut (.A(n32055), .B(n32054), .C(counter_hi[2]), 
         .D(\next_pc_for_core[6] ), .Z(n29147)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i26530_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_347_i2_3_lut_4_lut (.A(n32055), .B(n32054), .C(debug_ret), 
         .D(return_addr[2]), .Z(n34[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam mux_347_i2_3_lut_4_lut.init = 16'hf606;
    LUT4 i1_4_lut_adj_421 (.A(n9894), .B(n31867), .C(n27942), .D(n31809), 
         .Z(n27946)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_421.init = 16'h4000;
    LUT4 i1_4_lut_adj_422 (.A(no_write_in_progress), .B(data_ready_core), 
         .C(debug_instr_valid), .D(is_load), .Z(debug_rd_3__N_1575)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_4_lut_adj_422.init = 16'h8000;
    L6MUX21 mux_2147_i1 (.D0(n3505[0]), .D1(n3458[0]), .SD(n4285), .Z(n3546[0]));
    PFUMX mux_2147_i27 (.BLUT(n29049), .ALUT(n3458[26]), .C0(n29490), 
          .Z(n3546[26]));
    LUT4 i26958_3_lut (.A(imm[26]), .B(imm[30]), .C(counter_hi[2]), .Z(n29575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26958_3_lut.init = 16'hcaca;
    PFUMX mux_2147_i24 (.BLUT(n29028), .ALUT(n3458[23]), .C0(n29490), 
          .Z(n3546[23]));
    LUT4 mux_2138_i12_3_lut_4_lut (.A(n31718), .B(n31715), .C(n3422[11]), 
         .D(n2982[13]), .Z(n3505[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2138_i12_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_1826_i13_3_lut (.A(n31[12]), .B(n6[12]), .C(n2524), .Z(n2525[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i13_3_lut.init = 16'hcaca;
    PFUMX mux_2147_i23 (.BLUT(n29026), .ALUT(n3458[22]), .C0(n29490), 
          .Z(n3546[22]));
    LUT4 i26957_3_lut (.A(\imm[18] ), .B(\imm[22] ), .C(counter_hi[2]), 
         .Z(n29574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26957_3_lut.init = 16'hcaca;
    LUT4 i26956_3_lut (.A(\imm[10] ), .B(\imm[14] ), .C(counter_hi[2]), 
         .Z(n29573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26956_3_lut.init = 16'hcaca;
    LUT4 mux_1528_i1_3_lut (.A(n27[0]), .B(n31[0]), .C(n2504), .Z(n2143[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1538_i1_rep_111_3_lut (.A(n2163[0]), .B(instr[31]), .C(n4263), 
         .Z(n29057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1538_i1_rep_111_3_lut.init = 16'hcaca;
    LUT4 mux_1532_i1_3_lut (.A(n6[0]), .B(n21[0]), .C(n2524), .Z(n2163[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i1_3_lut.init = 16'hcaca;
    LUT4 mux_1538_i1_3_lut (.A(n2143[0]), .B(n2163[0]), .C(n31944), .Z(instr[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1538_i1_3_lut.init = 16'hcaca;
    PFUMX mux_2147_i22 (.BLUT(n29020), .ALUT(n3458[21]), .C0(n29490), 
          .Z(n3546[21]));
    LUT4 i26955_3_lut (.A(\imm[2] ), .B(\imm[6] ), .C(counter_hi[2]), 
         .Z(n29572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26955_3_lut.init = 16'hcaca;
    PFUMX mux_2147_i21 (.BLUT(n29018), .ALUT(n3458[20]), .C0(n29490), 
          .Z(n3546[20]));
    LUT4 i26951_3_lut (.A(imm[25]), .B(imm[29]), .C(counter_hi[2]), .Z(n29568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26951_3_lut.init = 16'hcaca;
    L6MUX21 mux_2147_i5 (.D0(n3505[4]), .D1(n3458[4]), .SD(n4285), .Z(n3546[4]));
    LUT4 i26950_3_lut (.A(\imm[17] ), .B(\imm[21] ), .C(counter_hi[2]), 
         .Z(n29567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26950_3_lut.init = 16'hcaca;
    PFUMX mux_2138_i1 (.BLUT(n3381[0]), .ALUT(n28881), .C0(n31718), .Z(n3505[0]));
    LUT4 mux_1822_i9_3_lut (.A(n21[8]), .B(n27[8]), .C(n2504), .Z(n2505[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i9_3_lut.init = 16'hcaca;
    L6MUX21 mux_2138_i6 (.D0(n3381[5]), .D1(n3422[5]), .SD(n31718), .Z(n3505[5]));
    LUT4 mux_1826_i9_3_lut (.A(n31[8]), .B(n6[8]), .C(n2524), .Z(n2525[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i9_3_lut.init = 16'hcaca;
    PFUMX mux_2138_i5 (.BLUT(n3381[4]), .ALUT(n3422[4]), .C0(n31718), 
          .Z(n3505[4]));
    LUT4 i1_4_lut_adj_423 (.A(clk_c_enable_448), .B(n31742), .C(n27724), 
         .D(n31738), .Z(n2136)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_423.init = 16'ha888;
    FD1P3AX rs2_i0_i1 (.D(n2243[1]), .SP(clk_c_enable_448), .CK(clk_c), 
            .Q(rs2[1])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i1.GSR = "DISABLED";
    FD1P3AX rs2_i0_i2 (.D(n2243[2]), .SP(clk_c_enable_448), .CK(clk_c), 
            .Q(rs2[2])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i2.GSR = "DISABLED";
    FD1P3AX rs2_i0_i3 (.D(n2243[3]), .SP(clk_c_enable_448), .CK(clk_c), 
            .Q(rs2[3])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam rs2_i0_i3.GSR = "DISABLED";
    LUT4 i26949_3_lut (.A(\imm[9] ), .B(\imm[13] ), .C(counter_hi[2]), 
         .Z(n29566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26949_3_lut.init = 16'hcaca;
    LUT4 i26948_3_lut (.A(\imm[1] ), .B(\imm[5] ), .C(counter_hi[2]), 
         .Z(n29565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26948_3_lut.init = 16'hcaca;
    LUT4 mux_1822_i8_3_lut (.A(n21[7]), .B(\instr_data[1][7] ), .C(n2504), 
         .Z(n2514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i8_3_lut.init = 16'hcaca;
    L6MUX21 mux_2147_i17 (.D0(n3505[16]), .D1(n3458[16]), .SD(n4285), 
            .Z(n3546[16]));
    LUT4 i26944_3_lut (.A(imm[24]), .B(imm[28]), .C(counter_hi[2]), .Z(n29561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26944_3_lut.init = 16'hcaca;
    PFUMX mux_2147_i16 (.BLUT(n3505[15]), .ALUT(n3458[15]), .C0(n4285), 
          .Z(n3546[15]));
    LUT4 i26943_3_lut (.A(\imm[16] ), .B(\imm[20] ), .C(counter_hi[2]), 
         .Z(n29560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26943_3_lut.init = 16'hcaca;
    LUT4 i26942_3_lut (.A(\imm[8] ), .B(\imm[12] ), .C(counter_hi[2]), 
         .Z(n29559)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26942_3_lut.init = 16'hcaca;
    LUT4 mux_1822_i10_3_lut (.A(n21[9]), .B(n27[9]), .C(n2504), .Z(n2505[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i10_3_lut.init = 16'hcaca;
    LUT4 i26941_3_lut (.A(imm[0]), .B(\imm[4] ), .C(counter_hi[2]), .Z(n29558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26941_3_lut.init = 16'hcaca;
    LUT4 mux_1826_i10_3_lut (.A(n31[9]), .B(n6[9]), .C(n2524), .Z(n2525[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i10_3_lut.init = 16'hcaca;
    LUT4 mux_1822_i4_3_lut (.A(n21[3]), .B(n27[3]), .C(n2504), .Z(n2505[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i4_3_lut.init = 16'hcaca;
    LUT4 mux_1826_i4_3_lut (.A(n31[3]), .B(n6[3]), .C(n2524), .Z(n2525[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i4_3_lut.init = 16'hcaca;
    PFUMX mux_2147_i15 (.BLUT(n3505[14]), .ALUT(n3458[14]), .C0(n4285), 
          .Z(n3546[14]));
    LUT4 i27618_3_lut_4_lut (.A(n31848), .B(n31714), .C(n4277), .D(n26794), 
         .Z(n3381[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27618_3_lut_4_lut.init = 16'hf808;
    PFUMX mux_2147_i14 (.BLUT(n3505[13]), .ALUT(n3458[13]), .C0(n4285), 
          .Z(n3546[13]));
    PFUMX mux_2147_i13 (.BLUT(n3505[12]), .ALUT(n3458[12]), .C0(n4285), 
          .Z(n3546[12]));
    PFUMX mux_2147_i12 (.BLUT(n3505[11]), .ALUT(n3458[11]), .C0(n4285), 
          .Z(n3546[11]));
    LUT4 i15415_2_lut (.A(\next_pc_for_core[4] ), .B(counter_hi[2]), .Z(n149)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i15415_2_lut.init = 16'h8888;
    PFUMX mux_2147_i11 (.BLUT(n3422[10]), .ALUT(n3505[10]), .C0(n29392), 
          .Z(n3546[10]));
    PFUMX i28321 (.BLUT(n31197), .ALUT(n31196), .C0(n31835), .Z(n31198));
    LUT4 mux_3126_i9_3_lut (.A(n31868), .B(instr[31]), .C(n4263), .Z(n5081[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3126_i9_3_lut.init = 16'hcaca;
    LUT4 i27922_2_lut (.A(counter_hi[4]), .B(n33486), .Z(n29337)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam i27922_2_lut.init = 16'heeee;
    LUT4 i2_2_lut_3_lut (.A(n31869), .B(n31860), .C(n31867), .Z(n17_adj_3142)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    defparam i2_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_3_lut_4_lut_3_lut (.A(n31869), .B(n31860), .C(n31868), .Z(n20)) /* synthesis lut_function=(A (B+(C))+!A !(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    defparam i1_3_lut_4_lut_3_lut.init = 16'hb9b9;
    LUT4 mux_3126_i8_3_lut (.A(n31845), .B(instr[31]), .C(n4263), .Z(n5081[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3126_i8_3_lut.init = 16'hcaca;
    PFUMX mux_2147_i9 (.BLUT(n3422[8]), .ALUT(n3505[8]), .C0(n29385), 
          .Z(n3546[8]));
    LUT4 mux_3126_i7_3_lut (.A(n31867), .B(instr[31]), .C(n4263), .Z(n5081[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3126_i7_3_lut.init = 16'hcaca;
    L6MUX21 mux_2147_i8 (.D0(n3505[7]), .D1(n3458[7]), .SD(n4285), .Z(n3546[7]));
    LUT4 mux_3126_i6_3_lut (.A(n31853), .B(instr[31]), .C(n4263), .Z(n5081[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3126_i6_3_lut.init = 16'hcaca;
    PFUMX mux_2110_i6 (.BLUT(n3195[5]), .ALUT(n26782), .C0(n4277), .Z(n3381[5]));
    LUT4 i2_4_lut (.A(n31940), .B(n31958), .C(n32033), .D(n32006), .Z(n10499)) /* synthesis lut_function=(A+!(B+(C (D)))) */ ;
    defparam i2_4_lut.init = 16'habbb;
    LUT4 i15570_2_lut_3_lut (.A(n31869), .B(n31860), .C(n15_adj_3143), 
         .Z(mem_op_de[0])) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    defparam i15570_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i2_2_lut_3_lut_adj_424 (.A(n31869), .B(n31860), .C(n31868), .Z(n20_adj_3144)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    defparam i2_2_lut_3_lut_adj_424.init = 16'h4040;
    LUT4 mux_1538_i11_3_lut (.A(n29051), .B(n2163[10]), .C(n31944), .Z(instr[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1538_i11_3_lut.init = 16'hcaca;
    LUT4 i15833_2_lut_3_lut_4_lut (.A(n31869), .B(n31845), .C(n31863), 
         .D(n31834), .Z(n30_adj_3145)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i15833_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i49_3_lut_3_lut (.A(n31869), .B(n31845), .C(n31860), .Z(n28)) /* synthesis lut_function=(!(A (C)+!A (B+!(C)))) */ ;
    defparam i49_3_lut_3_lut.init = 16'h1a1a;
    LUT4 is_system_I_0_481_2_lut_rep_782 (.A(is_system), .B(debug_instr_valid), 
         .Z(n31987)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam is_system_I_0_481_2_lut_rep_782.init = 16'h8888;
    LUT4 i1_2_lut_rep_687_3_lut_3_lut_4_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[1]), .D(alu_op[0]), .Z(n31892)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_687_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 additional_mem_ops_2__N_1132_0__bdd_2_lut_28320_3_lut_4_lut (.A(n31869), 
         .B(n31845), .C(n31865), .D(n31834), .Z(n31196)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam additional_mem_ops_2__N_1132_0__bdd_2_lut_28320_3_lut_4_lut.init = 16'h1000;
    LUT4 mux_1822_i2_3_lut (.A(n21[1]), .B(n27[1]), .C(n2504), .Z(n2505[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i2_3_lut.init = 16'hcaca;
    LUT4 is_system_I_0_3_lut_rep_743_4_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[1]), .D(alu_op[0]), .Z(n31948)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam is_system_I_0_3_lut_rep_743_4_lut.init = 16'h8880;
    LUT4 i26519_3_lut (.A(\next_pc_for_core[9] ), .B(\next_pc_for_core[13] ), 
         .C(counter_hi[2]), .Z(n29136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26519_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_689_3_lut_3_lut_4_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[1]), .D(alu_op[0]), .Z(n31894)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_689_3_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 data_from_read_10__bdd_3_lut_then_3_lut (.A(n31879), .B(n19), .C(n31885), 
         .Z(n32062)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam data_from_read_10__bdd_3_lut_then_3_lut.init = 16'hcece;
    LUT4 i1_2_lut_rep_709_2_lut_3_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[1]), .Z(n31914)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_709_2_lut_3_lut.init = 16'h8080;
    LUT4 i30_3_lut_4_lut_3_lut (.A(n31869), .B(n31868), .C(n31860), .Z(n13_adj_3146)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam i30_3_lut_4_lut_3_lut.init = 16'h1818;
    LUT4 i1_2_lut_rep_670_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut (.A(is_system), 
         .B(debug_instr_valid), .C(alu_op[1]), .D(alu_op[0]), .Z(n31875)) /* synthesis lut_function=(!(((C (D)+!C !(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam i1_2_lut_rep_670_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h0880;
    LUT4 i22_4_lut_4_lut (.A(n31868), .B(n31869), .C(n26113), .D(n31817), 
         .Z(n8_adj_3147)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam i22_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i1_3_lut_4_lut_4_lut_4_lut (.A(n31868), .B(n7), .C(n31786), .D(n31845), 
         .Z(n32)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_4_lut_4_lut.init = 16'h55fd;
    LUT4 i1_4_lut_4_lut_adj_425 (.A(n31868), .B(n31802), .C(n31809), .D(n31769), 
         .Z(is_lui_N_1365)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_425.init = 16'h4000;
    PFUMX mux_2138_i17 (.BLUT(n3271[16]), .ALUT(n3422[16]), .C0(n29428), 
          .Z(n3505[16]));
    LUT4 is_csr_I_0_573_2_lut_rep_710_4_lut_3_lut_4_lut (.A(is_system), .B(debug_instr_valid), 
         .C(alu_op[1]), .D(alu_op[0]), .Z(n31915)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(338[20:44])
    defparam is_csr_I_0_573_2_lut_rep_710_4_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_rep_590_3_lut_4_lut (.A(n31867), .B(n31868), .C(n31845), 
         .D(n31869), .Z(n31795)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_rep_590_3_lut_4_lut.init = 16'h0002;
    LUT4 debug_branch_I_48_i4_3_lut (.A(debug_branch_N_840[31]), .B(timer_data[3]), 
         .C(is_timer_addr), .Z(debug_branch_N_450[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_48_i4_3_lut.init = 16'hcaca;
    LUT4 i26531_3_lut (.A(\next_pc_for_core[10] ), .B(\next_pc_for_core[14] ), 
         .C(counter_hi[2]), .Z(n29148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26531_3_lut.init = 16'hcaca;
    PFUMX mux_2138_i8 (.BLUT(n3381[7]), .ALUT(n3422[7]), .C0(n31718), 
          .Z(n3505[7]));
    L6MUX21 mux_2138_i7 (.D0(n3381[6]), .D1(n3422[6]), .SD(n31718), .Z(n3505[6]));
    L6MUX21 mux_2138_i4 (.D0(n3381[3]), .D1(n3422[3]), .SD(n31718), .Z(n3505[3]));
    LUT4 next_pc_for_core_23__I_0_i269_4_lut (.A(n209), .B(n5677[0]), .C(n31955), 
         .D(n9033), .Z(debug_branch_N_446[28])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i269_4_lut.init = 16'haca0;
    L6MUX21 mux_2138_i2 (.D0(n3381[1]), .D1(n3422[1]), .SD(n31718), .Z(n3505[1]));
    PFUMX mux_1889_i3 (.BLUT(n26829), .ALUT(n2630[2]), .C0(n2812), .Z(n2644[2]));
    LUT4 data_from_read_10__bdd_3_lut_else_3_lut (.A(n31879), .B(n19), .C(\peri_data_out[10] ), 
         .D(n4), .Z(n32061)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam data_from_read_10__bdd_3_lut_else_3_lut.init = 16'heeec;
    LUT4 mux_1826_i2_3_lut (.A(n31[1]), .B(n6[1]), .C(n2524), .Z(n2525[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_426 (.A(n9894), .B(n26478), .C(n17998), .D(n28074), 
         .Z(n28080)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_426.init = 16'h0100;
    LUT4 i1_4_lut_adj_427 (.A(n2152), .B(n33488), .C(n29047), .D(n31944), 
         .Z(n28074)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_427.init = 16'hc088;
    LUT4 mux_1538_i7_rep_81_3_lut_3_lut (.A(n31732), .B(n31863), .C(n29045), 
         .Z(n29027)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1538_i7_rep_81_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_4_lut_adj_428 (.A(n9894), .B(n26478), .C(n17998), .D(n28086), 
         .Z(n28092)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_428.init = 16'h0100;
    LUT4 i1_4_lut_adj_429 (.A(n29033), .B(n33488), .C(n29045), .D(n31944), 
         .Z(n28086)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_429.init = 16'hc088;
    PFUMX i23915 (.BLUT(n13255), .ALUT(n13248), .C0(n26948), .Z(additional_mem_ops_2__N_749[2]));
    PFUMX i28611 (.BLUT(n32061), .ALUT(n32062), .C0(counter_hi[2]), .Z(n32063));
    LUT4 mux_1538_i8_rep_83_3_lut_3_lut (.A(n31732), .B(n31849), .C(n29047), 
         .Z(n29029)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1538_i8_rep_83_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_4_lut_adj_430 (.A(n9894), .B(n26478), .C(n17998), .D(n28098), 
         .Z(n28104)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_430.init = 16'h0100;
    LUT4 n4271_bdd_2_lut_4_lut (.A(n31838), .B(n31764), .C(n4281), .D(instr[29]), 
         .Z(n30835)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n4271_bdd_2_lut_4_lut.init = 16'hca00;
    LUT4 i1_4_lut_adj_431 (.A(n9894), .B(n26478), .C(n17998), .D(n28110), 
         .Z(n28116)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_431.init = 16'h0100;
    LUT4 mux_2101_i17_3_lut_4_lut (.A(n31733), .B(n31761), .C(n5081[9]), 
         .D(n2143[0]), .Z(n3340[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2101_i17_3_lut_4_lut.init = 16'hf870;
    PFUMX mux_2110_i9 (.BLUT(n26693), .ALUT(n26788), .C0(n4277), .Z(n3381[8]));
    LUT4 i1_3_lut (.A(no_write_in_progress), .B(debug_instr_valid), .C(is_store), 
         .Z(debug_rd_3__N_413)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i26575_3_lut (.A(\mem_data_from_read[19] ), .B(\mem_data_from_read[23] ), 
         .C(counter_hi[2]), .Z(n29192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26575_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_432 (.A(cycle[0]), .B(n10486), .C(n32039), .D(n28708), 
         .Z(n15_adj_3148)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_4_lut_adj_432.init = 16'hfffd;
    LUT4 i1_2_lut_adj_433 (.A(n33484), .B(cycle_c[1]), .Z(n28708)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(311[13:33])
    defparam i1_2_lut_adj_433.init = 16'heeee;
    LUT4 i2_2_lut_rep_515_3_lut_4_lut (.A(n31737), .B(n31742), .C(n31760), 
         .D(rst_reg_n), .Z(n31720)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i2_2_lut_rep_515_3_lut_4_lut.init = 16'h2000;
    LUT4 debug_branch_I_48_i1_3_lut (.A(n29160), .B(load_top_bit), .C(data_out_3__N_1385), 
         .Z(debug_branch_N_450[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_48_i1_3_lut.init = 16'hcaca;
    LUT4 debug_branch_I_48_i2_3_lut (.A(n29166), .B(load_top_bit), .C(data_out_3__N_1385), 
         .Z(debug_branch_N_450[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[18:66])
    defparam debug_branch_I_48_i2_3_lut.init = 16'hcaca;
    FD1S3IX counter_hi_3563__i3 (.D(n36[1]), .CK(clk_c), .CD(n31980), 
            .Q(counter_hi[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3563__i3.GSR = "DISABLED";
    FD1S3IX counter_hi_3563__i4 (.D(n36[2]), .CK(clk_c), .CD(n31980), 
            .Q(counter_hi[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3563__i4.GSR = "DISABLED";
    FD1S3IX addr_offset_3564__i3 (.D(n33[1]), .CK(clk_c), .CD(n31980), 
            .Q(addr_offset[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam addr_offset_3564__i3.GSR = "DISABLED";
    LUT4 n3301_bdd_4_lut_28031 (.A(n3271[2]), .B(n4279), .C(n31845), .D(n31847), 
         .Z(n30706)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B (C (D)))) */ ;
    defparam n3301_bdd_4_lut_28031.init = 16'he222;
    LUT4 i1_2_lut_rep_549 (.A(is_ret_de), .B(n33488), .Z(n31754)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_549.init = 16'h8888;
    PFUMX mux_2110_i7 (.BLUT(n3195[6]), .ALUT(n26776), .C0(n4277), .Z(n3381[6]));
    LUT4 i1_2_lut_3_lut_4_lut_adj_434 (.A(is_ret_de), .B(n33488), .C(n31743), 
         .D(n27018), .Z(n28028)) /* synthesis lut_function=(A (B (C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_434.init = 16'h8088;
    LUT4 i1_2_lut_rep_785 (.A(\instr_addr_23__N_318[0] ), .B(instr_addr_23__N_318[1]), 
         .Z(n31990)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_rep_785.init = 16'hbbbb;
    LUT4 i1_2_lut_2_lut_3_lut (.A(\instr_addr_23__N_318[0] ), .B(instr_addr_23__N_318[1]), 
         .C(n33488), .Z(n27972)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i1_2_lut_rep_786 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .Z(n31991)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_rep_786.init = 16'hbbbb;
    PFUMX mux_2110_i4 (.BLUT(n3195[3]), .ALUT(n26648), .C0(n4277), .Z(n3381[3]));
    LUT4 i27773_2_lut_3_lut (.A(n31737), .B(n31742), .C(n31860), .Z(n29210)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i27773_2_lut_3_lut.init = 16'hdfdf;
    LUT4 i1_2_lut_2_lut_3_lut_adj_435 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .C(n33488), .Z(n27966)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_2_lut_3_lut_adj_435.init = 16'hbfbf;
    PFUMX mux_2110_i2 (.BLUT(n26800), .ALUT(n3234[1]), .C0(n4277), .Z(n3381[1]));
    LUT4 i1_2_lut_rep_789 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .Z(n31994)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_rep_789.init = 16'heeee;
    LUT4 i1_2_lut_2_lut_3_lut_adj_436 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .C(n33488), .Z(n27978)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(428[21:56])
    defparam i1_2_lut_2_lut_3_lut_adj_436.init = 16'hefef;
    LUT4 i1_2_lut_rep_519_3_lut (.A(n31737), .B(n31742), .C(n33488), .Z(clk_c_enable_325)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i1_2_lut_rep_519_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_792 (.A(addr_c[26]), .B(addr_c[25]), .Z(n31997)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_792.init = 16'heeee;
    LUT4 i1_rep_132_2_lut_3_lut (.A(addr_c[26]), .B(addr_c[25]), .C(addr[27]), 
         .Z(n30171)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_rep_132_2_lut_3_lut.init = 16'hfefe;
    LUT4 i15666_2_lut_rep_734_3_lut_4_lut (.A(addr_c[26]), .B(addr_c[25]), 
         .C(n32033), .D(addr[27]), .Z(n31939)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i15666_2_lut_rep_734_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_rep_131_2_lut_3_lut (.A(addr_c[26]), .B(addr_c[25]), .C(addr[27]), 
         .Z(n30170)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_rep_131_2_lut_3_lut.init = 16'hfefe;
    PFUMX mux_2119_i7 (.BLUT(n3271[6]), .ALUT(n3304[6]), .C0(n4279), .Z(n3422[6]));
    LUT4 i1_2_lut_rep_517_3_lut_4_lut (.A(n31737), .B(n31742), .C(n31838), 
         .D(n33488), .Z(n31722)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam i1_2_lut_rep_517_3_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_753_3_lut (.A(addr_c[26]), .B(addr_c[25]), .C(addr[27]), 
         .Z(n31958)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_753_3_lut.init = 16'hfefe;
    LUT4 additional_mem_ops_1__bdd_3_lut_4_lut (.A(n31737), .B(n31742), 
         .C(n31200), .D(additional_mem_ops[1]), .Z(n4322[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(222[22:82])
    defparam additional_mem_ops_1__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 i26314_4_lut (.A(n31934), .B(n10467), .C(n26310), .D(n32027), 
         .Z(n13)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(352[54:66])
    defparam i26314_4_lut.init = 16'hcddd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_437 (.A(addr_c[26]), .B(addr_c[25]), .C(n32006), 
         .D(addr[27]), .Z(n26205)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_4_lut_adj_437.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_728_3_lut_4_lut (.A(addr_c[26]), .B(addr_c[25]), .C(n32033), 
         .D(addr[27]), .Z(clk_c_enable_268)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_728_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i27898_2_lut_rep_510 (.A(n4279), .B(n4271), .Z(n31715)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27898_2_lut_rep_510.init = 16'hbbbb;
    LUT4 i27598_3_lut_4_lut (.A(n4279), .B(n4271), .C(n3271[8]), .D(n2982[8]), 
         .Z(n3422[8])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27598_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i27924_2_lut_rep_732_3_lut_4_lut (.A(addr_c[26]), .B(addr_c[25]), 
         .C(counter_hi[4]), .D(addr[27]), .Z(n31937)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i27924_2_lut_rep_732_3_lut_4_lut.init = 16'hffef;
    LUT4 i27122_3_lut (.A(n29737), .B(n31418), .C(counter_hi[3]), .Z(n29739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27122_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_736_3_lut_4_lut (.A(addr_c[26]), .B(addr_c[25]), .C(n32006), 
         .D(addr[27]), .Z(n31941)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_736_3_lut_4_lut.init = 16'hfffe;
    LUT4 i27048_3_lut (.A(n29663), .B(n31408), .C(counter_hi[3]), .Z(n29665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27048_3_lut.init = 16'hcaca;
    PFUMX mux_2119_i6 (.BLUT(n3271[5]), .ALUT(n3304[5]), .C0(n4279), .Z(n3422[5]));
    PFUMX mux_2119_i4 (.BLUT(n3271[3]), .ALUT(n3304[3]), .C0(n4279), .Z(n3422[3]));
    LUT4 i1_2_lut_rep_550_4_lut (.A(n31817), .B(n31762), .C(n31868), .D(n31831), 
         .Z(n31755)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_550_4_lut.init = 16'h1000;
    PFUMX mux_2119_i2 (.BLUT(n3271[1]), .ALUT(n3304[1]), .C0(n4279), .Z(n3422[1]));
    LUT4 i27893_2_lut_3_lut_4_lut (.A(n4279), .B(n4271), .C(n4285), .D(n31718), 
         .Z(n29392)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27893_2_lut_3_lut_4_lut.init = 16'hf4f0;
    L6MUX21 mux_1889_i2 (.D0(n2621[1]), .D1(n2630[1]), .SD(n2812), .Z(n2644[1]));
    LUT4 is_lui_I_0_473_2_lut_rep_796 (.A(is_lui), .B(debug_instr_valid), 
         .Z(n32001)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam is_lui_I_0_473_2_lut_rep_796.init = 16'h8888;
    PFUMX mux_1889_i1 (.BLUT(n2621[0]), .ALUT(n2630[0]), .C0(n2812), .Z(n2644[0]));
    LUT4 next_pc_for_core_23__I_0_i157_3_lut (.A(\next_pc_for_core[8] ), .B(\next_pc_for_core[12] ), 
         .C(counter_hi[2]), .Z(n157_adj_3150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(351[34:46])
    defparam next_pc_for_core_23__I_0_i157_3_lut.init = 16'hcaca;
    PFUMX mux_2096_i8 (.BLUT(n5223[6]), .ALUT(n2982[7]), .C0(n4271), .Z(n3271[7]));
    LUT4 i26713_3_lut_4_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(n29337), 
         .D(n31999), .Z(n29330)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i26713_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 is_jalr_N_1372_bdd_2_lut_28458_4_lut (.A(n31817), .B(n31762), .C(n31868), 
         .D(n31763), .Z(n31441)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam is_jalr_N_1372_bdd_2_lut_28458_4_lut.init = 16'h1000;
    LUT4 i27920_2_lut_3_lut_4_lut_4_lut (.A(is_lui), .B(debug_instr_valid), 
         .C(is_jalr), .D(is_jal), .Z(n29333)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i27920_2_lut_3_lut_4_lut_4_lut.init = 16'hbbbf;
    LUT4 i27949_3_lut_4_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(n32007), 
         .D(n31999), .Z(n29240)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam i27949_3_lut_4_lut_4_lut.init = 16'hc888;
    PFUMX mux_2096_i5 (.BLUT(n5223[3]), .ALUT(n2982[4]), .C0(n4271), .Z(n3271[4]));
    LUT4 i27814_3_lut_4_lut (.A(n31764), .B(n31944), .C(n4281), .D(n4285), 
         .Z(n29490)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27814_3_lut_4_lut.init = 16'h1fff;
    LUT4 mux_91_i1_3_lut_4_lut (.A(is_lui), .B(debug_instr_valid), .C(debug_rd_3__N_405[28]), 
         .D(n157_adj_3150), .Z(n234[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(334[17:38])
    defparam mux_91_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1551_i1_4_lut (.A(n31846), .B(rs2[0]), .C(n31742), .D(mem_op_increment_reg), 
         .Z(n2222[0])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1551_i1_4_lut.init = 16'h3aca;
    LUT4 mtimecmp_6__I_0_3_lut_4_lut (.A(\addr[2] ), .B(n31871), .C(data_out_slice[2]), 
         .D(mtimecmp[6]), .Z(mtimecmp_2__N_1939)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(449[27:65])
    defparam mtimecmp_6__I_0_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_2123_i4 (.BLUT(n29029), .ALUT(n3340[3]), .C0(n29371), .Z(n3458[3]));
    LUT4 mtimecmp_7__I_0_3_lut_4_lut (.A(\addr[2] ), .B(n31871), .C(\data_out_slice[3] ), 
         .D(mtimecmp[7]), .Z(mtimecmp_3__N_1935)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(449[27:65])
    defparam mtimecmp_7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 mtimecmp_5__I_0_3_lut_4_lut (.A(\addr[2] ), .B(n31871), .C(data_out_slice[1]), 
         .D(mtimecmp[5]), .Z(mtimecmp_1__N_1941)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(449[27:65])
    defparam mtimecmp_5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 mtimecmp_4__I_0_3_lut_4_lut (.A(\addr[2] ), .B(n31871), .C(data_out_slice[0]), 
         .D(mtimecmp[4]), .Z(mtimecmp_0__N_1943)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(449[27:65])
    defparam mtimecmp_4__I_0_3_lut_4_lut.init = 16'hf780;
    FD1P3IX pc_offset__i1 (.D(pc_2__N_932[0]), .SP(clk_c_enable_527), .CD(n31980), 
            .CK(clk_c), .Q(\pc[1] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i1.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_438 (.A(n31766), .B(n31764), .C(n27746), .D(n9894), 
         .Z(n27750)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_adj_438.init = 16'h0070;
    LUT4 mux_1551_i2_4_lut (.A(n31852), .B(rs2[1]), .C(n31742), .D(n32050), 
         .Z(n2222[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1551_i2_4_lut.init = 16'h3aca;
    PFUMX mux_2123_i3 (.BLUT(n29027), .ALUT(n3340[2]), .C0(n29371), .Z(n3458[2]));
    L6MUX21 mux_1153_i4 (.D0(n5[3]), .D1(n2[3]), .SD(n2138), .Z(n1764[3]));
    LUT4 mux_1551_i3_4_lut (.A(n31847), .B(rs2[2]), .C(n31742), .D(n31975), 
         .Z(n2222[2])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1551_i3_4_lut.init = 16'h3aca;
    L6MUX21 mux_1153_i3 (.D0(n5[2]), .D1(n2[2]), .SD(n2138), .Z(n1764[2]));
    LUT4 mux_1551_i4_4_lut (.A(n31851), .B(rs2[3]), .C(n31742), .D(n6668), 
         .Z(n2222[3])) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1551_i4_4_lut.init = 16'h3aca;
    L6MUX21 mux_1153_i2 (.D0(n5[1]), .D1(n2[1]), .SD(n2138), .Z(n1764[1]));
    PFUMX mux_1874_i2 (.BLUT(n2589[1]), .ALUT(n2597[1]), .C0(n2808), .Z(n2621[1]));
    LUT4 i1_2_lut_rep_801 (.A(qv_data_read_n[0]), .B(qv_data_read_n[1]), 
         .Z(n32006)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_801.init = 16'h8888;
    LUT4 n31120_bdd_3_lut_4_lut (.A(n31764), .B(n31865), .C(n4281), .D(n31120), 
         .Z(n31121)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n31120_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_3_lut_4_lut_adj_439 (.A(qv_data_read_n[0]), .B(qv_data_read_n[1]), 
         .C(data_ready_r), .D(n31905), .Z(n28760)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_439.init = 16'h0700;
    LUT4 i1_4_lut_adj_440 (.A(n31743), .B(n26993), .C(n31744), .D(n28182), 
         .Z(clk_c_enable_134)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;
    defparam i1_4_lut_adj_440.init = 16'h3332;
    LUT4 mux_345_i1_3_lut (.A(\next_pc_for_core[3] ), .B(return_addr[3]), 
         .C(debug_ret), .Z(n1742[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i1_3_lut.init = 16'hcaca;
    LUT4 i26628_2_lut_rep_802 (.A(counter_hi[4]), .B(counter_hi[3]), .Z(n32007)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam i26628_2_lut_rep_802.init = 16'h4444;
    LUT4 i26603_2_lut_3_lut (.A(n33484), .B(n33486), .C(alu_a_in_3__N_1552), 
         .Z(n29220)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam i26603_2_lut_3_lut.init = 16'h4040;
    LUT4 i27537_3_lut_4_lut (.A(n31846), .B(n31773), .C(n2498), .D(n26871), 
         .Z(n2232[0])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27537_3_lut_4_lut.init = 16'hefe0;
    LUT4 i2_2_lut_3_lut_4_lut (.A(n33488), .B(clk_c_enable_30), .C(n22_adj_3135), 
         .D(n31838), .Z(n2808)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 pc_23__I_0_450_i269_rep_66_3_lut_4_lut (.A(counter_hi[4]), .B(counter_hi[3]), 
         .C(n209_adj_3151), .D(n157_adj_3152), .Z(n29012)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam pc_23__I_0_450_i269_rep_66_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i27557_3_lut_4_lut_4_lut (.A(n31773), .B(n26889), .C(n2498), 
         .D(n31851), .Z(n2232[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam i27557_3_lut_4_lut_4_lut.init = 16'hfc5c;
    PFUMX mux_1889_i4 (.BLUT(n26905), .ALUT(n2630[3]), .C0(n2812), .Z(n2644[3]));
    FD1P3IX pc_offset__i23 (.D(pc_23__N_911[20]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[23] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i23.GSR = "DISABLED";
    FD1P3IX pc_offset__i22 (.D(pc_23__N_911[19]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[22] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i22.GSR = "DISABLED";
    FD1P3IX pc_offset__i21 (.D(pc_23__N_911[18]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[21] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i21.GSR = "DISABLED";
    FD1P3IX pc_offset__i20 (.D(pc_23__N_911[17]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[20] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i20.GSR = "DISABLED";
    FD1P3IX pc_offset__i19 (.D(pc_23__N_911[16]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[19] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i19.GSR = "DISABLED";
    FD1P3IX pc_offset__i18 (.D(pc_23__N_911[15]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[18] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i18.GSR = "DISABLED";
    FD1P3IX pc_offset__i17 (.D(pc_23__N_911[14]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[17] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i17.GSR = "DISABLED";
    FD1P3IX pc_offset__i16 (.D(pc_23__N_911[13]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[16] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i16.GSR = "DISABLED";
    FD1P3IX pc_offset__i15 (.D(pc_23__N_911[12]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[15] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i15.GSR = "DISABLED";
    FD1P3IX pc_offset__i14 (.D(pc_23__N_911[11]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[14] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i14.GSR = "DISABLED";
    FD1P3IX pc_offset__i13 (.D(pc_23__N_911[10]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[13] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i13.GSR = "DISABLED";
    FD1P3IX pc_offset__i12 (.D(pc_23__N_911[9]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[12] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i12.GSR = "DISABLED";
    FD1P3IX pc_offset__i11 (.D(pc_23__N_911[8]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[11] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i11.GSR = "DISABLED";
    FD1P3IX pc_offset__i10 (.D(pc_23__N_911[7]), .SP(clk_c_enable_527), 
            .CD(n31980), .CK(clk_c), .Q(\pc[10] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i10.GSR = "DISABLED";
    FD1P3IX pc_offset__i9 (.D(pc_23__N_911[6]), .SP(clk_c_enable_527), .CD(n31980), 
            .CK(clk_c), .Q(\pc[9] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i9.GSR = "DISABLED";
    FD1P3IX pc_offset__i8 (.D(pc_23__N_911[5]), .SP(clk_c_enable_527), .CD(n31980), 
            .CK(clk_c), .Q(\pc[8] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i8.GSR = "DISABLED";
    LUT4 i27555_3_lut_4_lut_4_lut (.A(n31773), .B(n26883), .C(n2498), 
         .D(n31847), .Z(n2232[2])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam i27555_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_345_i2_3_lut (.A(\next_pc_for_core[4] ), .B(return_addr[4]), 
         .C(debug_ret), .Z(n1742[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i2_3_lut.init = 16'hcaca;
    FD1P3IX pc_offset__i7 (.D(pc_23__N_911[4]), .SP(clk_c_enable_527), .CD(n31980), 
            .CK(clk_c), .Q(\pc[7] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i7.GSR = "DISABLED";
    LUT4 mux_345_i3_3_lut (.A(\next_pc_for_core[5] ), .B(return_addr[5]), 
         .C(debug_ret), .Z(n1742[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i3_3_lut.init = 16'hcaca;
    FD1P3IX pc_offset__i6 (.D(pc_23__N_911[3]), .SP(clk_c_enable_527), .CD(n31980), 
            .CK(clk_c), .Q(\pc[6] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i6.GSR = "DISABLED";
    FD1P3IX pc_offset__i5 (.D(pc_23__N_911[2]), .SP(clk_c_enable_527), .CD(n31980), 
            .CK(clk_c), .Q(\pc[5] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i5.GSR = "DISABLED";
    FD1P3IX pc_offset__i4 (.D(pc_23__N_911[1]), .SP(clk_c_enable_527), .CD(n31980), 
            .CK(clk_c), .Q(\pc[4] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i4.GSR = "DISABLED";
    LUT4 i27553_3_lut_4_lut_4_lut (.A(n31773), .B(n26877), .C(n2498), 
         .D(n31852), .Z(n2232[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam i27553_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_345_i4_3_lut (.A(\next_pc_for_core[6] ), .B(return_addr[6]), 
         .C(debug_ret), .Z(n1742[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i4_3_lut.init = 16'hcaca;
    LUT4 mux_345_i5_3_lut (.A(\next_pc_for_core[7] ), .B(return_addr[7]), 
         .C(debug_ret), .Z(n1742[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i5_3_lut.init = 16'hcaca;
    LUT4 mux_345_i6_3_lut (.A(\next_pc_for_core[8] ), .B(return_addr[8]), 
         .C(debug_ret), .Z(n1742[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i6_3_lut.init = 16'hcaca;
    LUT4 mux_345_i7_3_lut (.A(\next_pc_for_core[9] ), .B(return_addr[9]), 
         .C(debug_ret), .Z(n1742[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i7_3_lut.init = 16'hcaca;
    LUT4 mux_345_i8_3_lut (.A(\next_pc_for_core[10] ), .B(return_addr[10]), 
         .C(debug_ret), .Z(n1742[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i8_3_lut.init = 16'hcaca;
    LUT4 mux_40_i1_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[28]), 
         .D(data_rs2[0]), .Z(n92[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i24_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(\debug_rd_3__N_405[31] ), 
         .D(n84), .Z(n92[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam i24_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i9_3_lut (.A(\next_pc_for_core[11] ), .B(return_addr[11]), 
         .C(debug_ret), .Z(n1742[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i9_3_lut.init = 16'hcaca;
    LUT4 mux_40_i3_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[30]), 
         .D(data_rs2[2]), .Z(n92[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i10_3_lut (.A(\next_pc_for_core[12] ), .B(return_addr[12]), 
         .C(debug_ret), .Z(n1742[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i10_3_lut.init = 16'hcaca;
    LUT4 i16_4_lut (.A(n27614), .B(clk_c_enable_30), .C(rst_reg_n), .D(n31719), 
         .Z(clk_c_enable_212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i16_4_lut.init = 16'hcfca;
    LUT4 mux_40_i2_3_lut_4_lut (.A(is_alu_imm), .B(debug_instr_valid), .C(debug_rd_3__N_405[29]), 
         .D(data_rs2[1]), .Z(n92[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(330[21:46])
    defparam mux_40_i2_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_1564_i4 (.BLUT(n2232[3]), .ALUT(n2222[3]), .C0(n2500), .Z(n2243[3]));
    LUT4 mux_345_i11_3_lut (.A(\next_pc_for_core[13] ), .B(return_addr[13]), 
         .C(debug_ret), .Z(n1742[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i11_3_lut.init = 16'hcaca;
    PFUMX mux_1564_i3 (.BLUT(n2232[2]), .ALUT(n2222[2]), .C0(n2500), .Z(n2243[2]));
    LUT4 mux_345_i12_3_lut (.A(\next_pc_for_core[14] ), .B(return_addr[14]), 
         .C(debug_ret), .Z(n1742[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i12_3_lut.init = 16'hcaca;
    PFUMX mux_1564_i2 (.BLUT(n2232[1]), .ALUT(n2222[1]), .C0(n2500), .Z(n2243[1]));
    LUT4 mux_345_i13_3_lut (.A(\next_pc_for_core[15] ), .B(return_addr[15]), 
         .C(debug_ret), .Z(n1742[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i13_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_441 (.A(n4285), .B(n31744), .C(n31738), .D(n27994), 
         .Z(n27614)) /* synthesis lut_function=(A+!(B+!(C (D)))) */ ;
    defparam i1_4_lut_adj_441.init = 16'hbaaa;
    FD1P3IX pc_offset__i3 (.D(pc_23__N_911[0]), .SP(clk_c_enable_527), .CD(n31980), 
            .CK(clk_c), .Q(\pc[3] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i3.GSR = "DISABLED";
    FD1P3IX pc_offset__i2 (.D(pc_2__N_932[1]), .SP(clk_c_enable_527), .CD(n31980), 
            .CK(clk_c), .Q(\pc[2] ));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam pc_offset__i2.GSR = "DISABLED";
    LUT4 is_branch_I_0_475_2_lut_rep_810 (.A(is_branch), .B(debug_instr_valid), 
         .Z(n32015)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam is_branch_I_0_475_2_lut_rep_810.init = 16'h8888;
    LUT4 mux_844_i3_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[5] ), 
         .D(addr_out[5]), .Z(n1215[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 n31117_bdd_3_lut (.A(n31117), .B(n31865), .C(n4263), .Z(n31118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31117_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_442 (.A(n31742), .B(n35), .C(n28006), .D(n26), 
         .Z(n27994)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i1_4_lut_adj_442.init = 16'h5040;
    LUT4 mux_3079_i1_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(n32016), .D(addr_out[1]), .Z(n5014[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_3079_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i14_3_lut (.A(\next_pc_for_core[16] ), .B(return_addr[16]), 
         .C(debug_ret), .Z(n1742[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i14_3_lut.init = 16'hcaca;
    PFUMX mux_1143_i4 (.BLUT(n26827), .ALUT(n1720[3]), .C0(n2134), .Z(n5[3]));
    LUT4 mux_844_i4_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[6] ), 
         .D(addr_out[6]), .Z(n1215[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i15_3_lut (.A(\next_pc_for_core[17] ), .B(return_addr[17]), 
         .C(debug_ret), .Z(n1742[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i15_3_lut.init = 16'hcaca;
    L6MUX21 i26947 (.D0(n29562), .D1(n29563), .SD(counter_hi[4]), .Z(debug_rd_3__N_405[28]));
    PFUMX mux_1143_i3 (.BLUT(n26814), .ALUT(n1720[2]), .C0(n2134), .Z(n5[2]));
    LUT4 i1_3_lut_3_lut (.A(n31742), .B(n32076), .C(n9894), .Z(n27672)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i1_3_lut_3_lut.init = 16'h0404;
    LUT4 mux_345_i16_3_lut (.A(\next_pc_for_core[18] ), .B(return_addr[18]), 
         .C(debug_ret), .Z(n1742[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i16_3_lut.init = 16'hcaca;
    LUT4 mux_3079_i2_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[2] ), .D(n31898), .Z(n5014[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_3079_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i17_3_lut (.A(\next_pc_for_core[19] ), .B(return_addr[19]), 
         .C(debug_ret), .Z(n1742[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i17_3_lut.init = 16'hcaca;
    LUT4 mux_345_i18_3_lut (.A(\next_pc_for_core[20] ), .B(return_addr[20]), 
         .C(debug_ret), .Z(n1742[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i18_3_lut.init = 16'hcaca;
    PFUMX mux_1143_i2 (.BLUT(n26807), .ALUT(n1720[1]), .C0(n2134), .Z(n5[1]));
    LUT4 i1_3_lut_adj_443 (.A(n31867), .B(n31473), .C(n28), .Z(n26)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_adj_443.init = 16'hecec;
    LUT4 mux_844_i2_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[4] ), 
         .D(addr_out[4]), .Z(n1215[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i2_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_2123_i17 (.BLUT(n3340[16]), .ALUT(n5121[16]), .C0(n4281), 
          .Z(n3458[16]));
    LUT4 mux_844_i1_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[3] ), 
         .D(addr_out[3]), .Z(n1215[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_844_i5_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[7] ), 
         .D(addr_out[7]), .Z(n1215[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i14129_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[8] ), 
         .D(addr_out[8]), .Z(n1215[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam i14129_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_844_i7_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[9] ), 
         .D(addr_out[9]), .Z(n1215[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_844_i8_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[10] ), 
         .D(addr_out[10]), .Z(n1215[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i19_3_lut (.A(\next_pc_for_core[21] ), .B(return_addr[21]), 
         .C(debug_ret), .Z(n1742[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i19_3_lut.init = 16'hcaca;
    LUT4 mux_844_i9_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), .C(\early_branch_addr[11] ), 
         .D(addr_out[11]), .Z(n1215[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_844_i10_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[12] ), .D(addr_out[12]), .Z(n1215[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i10_3_lut_4_lut.init = 16'hf780;
    L6MUX21 i26954 (.D0(n29569), .D1(n29570), .SD(n33484), .Z(debug_rd_3__N_405[29]));
    LUT4 mux_844_i11_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[13] ), .D(addr_out[13]), .Z(n1215[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i11_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_2123_i5 (.BLUT(n3340[4]), .ALUT(n5121[4]), .C0(n4281), .Z(n3458[4]));
    LUT4 mux_844_i12_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[14] ), .D(addr_out[14]), .Z(n1215[11])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_844_i13_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[15] ), .D(addr_out[15]), .Z(n1215[12])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i20_3_lut (.A(\next_pc_for_core[22] ), .B(return_addr[22]), 
         .C(debug_ret), .Z(n1742[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i20_3_lut.init = 16'hcaca;
    LUT4 mux_844_i14_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[16] ), .D(addr_out[16]), .Z(n1215[13])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_844_i15_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[17] ), .D(addr_out[17]), .Z(n1215[14])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_345_i21_3_lut (.A(\next_pc_for_core[23] ), .B(return_addr[23]), 
         .C(debug_ret), .Z(n1742[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(416[18] 430[16])
    defparam mux_345_i21_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_444 (.A(n31838), .B(clk_c_enable_325), .C(n31831), 
         .D(n31830), .Z(n4285)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;
    defparam i2_4_lut_adj_444.init = 16'hc888;
    LUT4 i1_2_lut_4_lut_adj_445 (.A(n32034), .B(n31880), .C(n32027), .D(data_to_write[6]), 
         .Z(\gpio_out_sel_7__N_13[0] )) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_4_lut_adj_445.init = 16'h4000;
    LUT4 i6902_4_lut (.A(n29051), .B(instr[26]), .C(n4281), .D(n31764), 
         .Z(n3340[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i6902_4_lut.init = 16'hca0a;
    LUT4 i1_rep_520_4_lut (.A(debug_ret), .B(n27286), .C(n31745), .D(n10499), 
         .Z(n31725)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_rep_520_4_lut.init = 16'h0010;
    LUT4 mux_844_i16_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[18] ), .D(addr_out[18]), .Z(n1215[15])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1832_i15_3_lut_rep_640 (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .Z(n31845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i15_3_lut_rep_640.init = 16'hcaca;
    LUT4 i1_2_lut_rep_597_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31867), .Z(n31802)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_597_4_lut.init = 16'hca00;
    PFUMX mux_1147_i4 (.BLUT(n1725[3]), .ALUT(n26996), .C0(n2136), .Z(n2[3]));
    PFUMX i28265 (.BLUT(n31119), .ALUT(n31118), .C0(n31733), .Z(n31120));
    LUT4 i38_3_lut (.A(n31869), .B(n31860), .C(n24_adj_3160), .Z(n22)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;
    defparam i38_3_lut.init = 16'h9898;
    LUT4 mux_844_i17_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[19] ), .D(addr_out[19]), .Z(n1215[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 n4263_bdd_3_lut_28267 (.A(n29043), .B(n29025), .C(n31944), .Z(n31117)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n4263_bdd_3_lut_28267.init = 16'hacac;
    LUT4 i27604_3_lut (.A(n3340[12]), .B(n5121[12]), .C(n4281), .Z(n3458[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27604_3_lut.init = 16'hcaca;
    LUT4 i27841_2_lut_rep_603_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31860), .Z(n31808)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i27841_2_lut_rep_603_4_lut.init = 16'h00ca;
    L6MUX21 i26961 (.D0(n29576), .D1(n29577), .SD(n33484), .Z(debug_rd_3__N_405[30]));
    LUT4 mux_844_i18_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[20] ), .D(addr_out[20]), .Z(n1215[17])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i18_3_lut_4_lut.init = 16'hf780;
    L6MUX21 i26983 (.D0(n29598), .D1(n29599), .SD(n33484), .Z(\debug_rd_3__N_405[31] ));
    LUT4 i27606_3_lut (.A(n3340[13]), .B(n5121[13]), .C(n4281), .Z(n3458[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27606_3_lut.init = 16'hcaca;
    LUT4 mux_844_i19_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[21] ), .D(addr_out[21]), .Z(n1215[18])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i19_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_1147_i3 (.BLUT(n1725[2]), .ALUT(n26995), .C0(n2136), .Z(n2[2]));
    LUT4 i27608_3_lut (.A(n3340[14]), .B(n5121[14]), .C(n4281), .Z(n3458[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27608_3_lut.init = 16'hcaca;
    PFUMX mux_1147_i2 (.BLUT(n1725[1]), .ALUT(n26997), .C0(n2136), .Z(n2[1]));
    LUT4 mux_2101_i12_3_lut_4_lut (.A(n4281), .B(n31733), .C(n5081[4]), 
         .D(n29023), .Z(n3340[11])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2101_i12_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i27610_3_lut (.A(n3340[15]), .B(n5121[15]), .C(n4281), .Z(n3458[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27610_3_lut.init = 16'hcaca;
    PFUMX pc_23__I_0_450_i209 (.BLUT(n149_adj_3161), .ALUT(n225), .C0(n33484), 
          .Z(n209_adj_3151)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 mux_844_i20_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[22] ), .D(addr_out[22]), .Z(n1215[19])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i20_3_lut_4_lut.init = 16'hf780;
    PFUMX mux_1879_i2 (.BLUT(n10904), .ALUT(n2607[1]), .C0(n2810), .Z(n2630[1]));
    LUT4 additional_mem_ops_2__N_1132_0__bdd_2_lut_28323_4_lut (.A(n2505[14]), 
         .B(n2525[14]), .C(n31944), .D(additional_mem_ops_2__N_1132[0]), 
         .Z(n31197)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam additional_mem_ops_2__N_1132_0__bdd_2_lut_28323_4_lut.init = 16'hca00;
    LUT4 i15612_2_lut_rep_612_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31867), .Z(n31817)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15612_2_lut_rep_612_4_lut.init = 16'hffca;
    PFUMX mux_1564_i1 (.BLUT(n2232[0]), .ALUT(n2222[0]), .C0(n2500), .Z(n2243[0]));
    LUT4 i15394_2_lut (.A(\pc[4] ), .B(counter_hi[2]), .Z(n149_adj_3161)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam i15394_2_lut.init = 16'h8888;
    LUT4 i23825_2_lut_rep_598_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31868), .Z(n31803)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i23825_2_lut_rep_598_4_lut.init = 16'hffca;
    LUT4 i1_4_lut_adj_446 (.A(n31741), .B(n8), .C(n31748), .D(n28174), 
         .Z(debug_early_branch)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_446.init = 16'h0200;
    LUT4 i1_2_lut_adj_447 (.A(is_jal_de), .B(rst_reg_n), .Z(n28174)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_447.init = 16'h8888;
    LUT4 mux_844_i21_3_lut_4_lut (.A(is_branch), .B(debug_instr_valid), 
         .C(\early_branch_addr[23] ), .D(addr_out[23]), .Z(n1215[20])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(335[20:44])
    defparam mux_844_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_448 (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31864), .Z(n2602[0])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_448.init = 16'h3500;
    LUT4 i27891_3_lut_4_lut (.A(n4263), .B(n31944), .C(n31733), .D(n4281), 
         .Z(n29400)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27891_3_lut_4_lut.init = 16'hff1f;
    PFUMX mux_1143_i1 (.BLUT(n26821), .ALUT(n1724), .C0(n2134), .Z(n5[0]));
    LUT4 i1_2_lut_2_lut_rep_594_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31867), .Z(n31799)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_2_lut_rep_594_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_814 (.A(\addr[2] ), .B(\addr[3] ), .Z(n32019)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_814.init = 16'hdddd;
    LUT4 n4263_bdd_4_lut_28270 (.A(n31838), .B(n29043), .C(n29025), .D(n31944), 
         .Z(n31119)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n4263_bdd_4_lut_28270.init = 16'h88a0;
    LUT4 i1_2_lut_rep_730_3_lut_4_lut (.A(\addr[2] ), .B(\addr[3] ), .C(n32034), 
         .D(n32035), .Z(n31935)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_730_3_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_815 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .Z(n32020)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_815.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_449 (.A(n27310), .B(n31736), .C(n33479), .D(n31906), 
         .Z(n1176)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/mem_ctrl.v(61[10:25])
    defparam i1_3_lut_4_lut_adj_449.init = 16'hf1ff;
    LUT4 i1_2_lut_3_lut_adj_450 (.A(instr_addr_23__N_318[1]), .B(\instr_addr_23__N_318[0] ), 
         .C(n33488), .Z(n27998)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_450.init = 16'h8080;
    LUT4 i1_2_lut_rep_816 (.A(qv_data_write_n[1]), .B(qv_data_read_n[1]), 
         .Z(n32021)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(270[12] 304[8])
    defparam i1_2_lut_rep_816.init = 16'h8888;
    LUT4 i15582_2_lut_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31863), .Z(n2602[2])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15582_2_lut_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_rep_609_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31868), .Z(n31814)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_609_4_lut.init = 16'hcaff;
    LUT4 additional_mem_ops_2__N_1132_0__bdd_2_lut_4_lut (.A(n2505[14]), .B(n2525[14]), 
         .C(n31944), .D(additional_mem_ops_2__N_1132[0]), .Z(n31402)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam additional_mem_ops_2__N_1132_0__bdd_2_lut_4_lut.init = 16'h00ca;
    LUT4 mux_2101_i5_3_lut (.A(n31848), .B(instr[24]), .C(n31732), .Z(n3340[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2101_i5_3_lut.init = 16'hcaca;
    LUT4 i15583_2_lut_rep_602_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31849), .Z(n31807)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15583_2_lut_rep_602_4_lut.init = 16'h3500;
    LUT4 i1_2_lut_rep_817 (.A(qv_data_write_n[0]), .B(qv_data_read_n[0]), 
         .Z(n32022)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_817.init = 16'h8888;
    PFUMX mux_2123_i1 (.BLUT(n27246), .ALUT(n5121[0]), .C0(n4281), .Z(n3458[0]));
    LUT4 i15372_2_lut_3_lut_4_lut (.A(qv_data_write_n[0]), .B(qv_data_read_n[0]), 
         .C(qv_data_read_n[1]), .D(qv_data_write_n[1]), .Z(n18588)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15372_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i27317_3_lut_3_lut (.A(\imm[10] ), .B(n9538), .C(n5624[2]), .Z(n5659[2])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i27317_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_1538_i5_rep_73_3_lut (.A(n29041), .B(n31864), .C(n4263), 
         .Z(n29019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1538_i5_rep_73_3_lut.init = 16'hcaca;
    PFUMX mux_55_i1 (.BLUT(n8302), .ALUT(additional_mem_ops_de[0]), .C0(n29210), 
          .Z(n4322[0])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i27602_3_lut (.A(n29019), .B(n3340[11]), .C(n29400), .Z(n3458[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i27602_3_lut.init = 16'hcaca;
    PFUMX mux_2123_i7 (.BLUT(n29048), .ALUT(n3340[6]), .C0(n29375), .Z(n3458[6]));
    LUT4 i1_2_lut_rep_821 (.A(debug_instr_valid), .B(no_write_in_progress), 
         .Z(n32026)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_2_lut_rep_821.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_451 (.A(debug_instr_valid), .B(no_write_in_progress), 
         .C(load_done), .D(is_load), .Z(instr_complete_N_1651)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_3_lut_4_lut_adj_451.init = 16'h8000;
    PFUMX mux_845_i21 (.BLUT(n1742[20]), .ALUT(n1215[20]), .C0(n31748), 
          .Z(pc_23__N_911[20]));
    PFUMX mux_845_i20 (.BLUT(n1742[19]), .ALUT(n1215[19]), .C0(n30169), 
          .Z(pc_23__N_911[19]));
    PFUMX mux_845_i19 (.BLUT(n1742[18]), .ALUT(n1215[18]), .C0(n30169), 
          .Z(pc_23__N_911[18]));
    PFUMX mux_845_i18 (.BLUT(n1742[17]), .ALUT(n1215[17]), .C0(n30169), 
          .Z(pc_23__N_911[17]));
    PFUMX mux_845_i17 (.BLUT(n1742[16]), .ALUT(n1215[16]), .C0(n30169), 
          .Z(pc_23__N_911[16]));
    PFUMX mux_845_i16 (.BLUT(n1742[15]), .ALUT(n1215[15]), .C0(n30168), 
          .Z(pc_23__N_911[15]));
    LUT4 i26433_3_lut_rep_824 (.A(counter_hi[2]), .B(counter_hi[3]), .C(counter_hi[4]), 
         .Z(n32029)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i26433_3_lut_rep_824.init = 16'h8080;
    LUT4 i27670_2_lut_4_lut (.A(counter_hi[2]), .B(counter_hi[3]), .C(counter_hi[4]), 
         .D(rst_reg_n), .Z(clk_c_enable_20)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;
    defparam i27670_2_lut_4_lut.init = 16'h80ff;
    PFUMX mux_845_i15 (.BLUT(n1742[14]), .ALUT(n1215[14]), .C0(n30168), 
          .Z(pc_23__N_911[14]));
    LUT4 i21218_3_lut_4_lut (.A(n27846), .B(n31738), .C(addr_offset[2]), 
         .D(n31742), .Z(n33[0])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (D)+!B !(C (D)+!C !(D))))) */ ;
    defparam i21218_3_lut_4_lut.init = 16'h4fb0;
    PFUMX mux_845_i14 (.BLUT(n1742[13]), .ALUT(n1215[13]), .C0(n30168), 
          .Z(pc_23__N_911[13]));
    LUT4 i1_2_lut_rep_625_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31868), .Z(n31830)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_625_4_lut.init = 16'hca00;
    PFUMX mux_845_i13 (.BLUT(n1742[12]), .ALUT(n1215[12]), .C0(n30168), 
          .Z(pc_23__N_911[12]));
    LUT4 i1_4_lut_adj_452 (.A(n31884), .B(data_ready_ext), .C(data_ready_sync), 
         .D(clk_c_enable_36), .Z(clk_c_enable_224)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_452.init = 16'hfeee;
    PFUMX mux_845_i12 (.BLUT(n1742[11]), .ALUT(n1215[11]), .C0(n30167), 
          .Z(pc_23__N_911[11]));
    PFUMX mux_845_i11 (.BLUT(n1742[10]), .ALUT(n1215[10]), .C0(n30167), 
          .Z(pc_23__N_911[10]));
    LUT4 i15804_2_lut_2_lut_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31850), .Z(n5223[6])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15804_2_lut_2_lut_4_lut.init = 16'h3500;
    LUT4 i15802_2_lut_2_lut_4_lut (.A(n2505[14]), .B(n2525[14]), .C(n31944), 
         .D(n31848), .Z(n5223[3])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15802_2_lut_2_lut_4_lut.init = 16'h3500;
    LUT4 mux_1832_i3_3_lut_rep_641 (.A(n2505[2]), .B(n2525[2]), .C(n31944), 
         .Z(n31846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i3_3_lut_rep_641.init = 16'hcaca;
    PFUMX mux_845_i10 (.BLUT(n1742[9]), .ALUT(n1215[9]), .C0(n30167), 
          .Z(pc_23__N_911[9]));
    LUT4 i1_2_lut_adj_453 (.A(\pc[1] ), .B(\instr_addr_23__N_318[0] ), .Z(n28260)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(157[53:124])
    defparam i1_2_lut_adj_453.init = 16'hdddd;
    PFUMX mux_845_i9 (.BLUT(n1742[8]), .ALUT(n1215[8]), .C0(n30167), .Z(pc_23__N_911[8]));
    PFUMX mux_845_i8 (.BLUT(n1742[7]), .ALUT(n1215[7]), .C0(n30166), .Z(pc_23__N_911[7]));
    PFUMX mux_845_i7 (.BLUT(n1742[6]), .ALUT(n1215[6]), .C0(n30166), .Z(pc_23__N_911[6]));
    LUT4 data_ready_I_0_4_lut (.A(mem_data_ready), .B(n18518), .C(data_ready), 
         .D(n31958), .Z(data_ready_ext)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(231[27:66])
    defparam data_ready_I_0_4_lut.init = 16'h3022;
    LUT4 i1_3_lut_adj_454 (.A(next_pc_offset[3]), .B(n4_adj_3138), .C(\instr_write_offset[3] ), 
         .Z(n27056)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;
    defparam i1_3_lut_adj_454.init = 16'h9696;
    PFUMX mux_845_i6 (.BLUT(n1742[5]), .ALUT(n1215[5]), .C0(n30166), .Z(pc_23__N_911[5]));
    PFUMX mux_845_i5 (.BLUT(n1742[4]), .ALUT(n1215[4]), .C0(n30166), .Z(pc_23__N_911[4]));
    PFUMX mux_845_i4 (.BLUT(n1742[3]), .ALUT(n1215[3]), .C0(n30165), .Z(pc_23__N_911[3]));
    LUT4 instr_6__I_0_126_i6_2_lut_rep_611_4_lut (.A(n2505[2]), .B(n2525[2]), 
         .C(n31944), .D(n31852), .Z(n31816)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_6__I_0_126_i6_2_lut_rep_611_4_lut.init = 16'hff35;
    PFUMX mux_845_i3 (.BLUT(n1742[2]), .ALUT(n1215[2]), .C0(n30165), .Z(pc_23__N_911[2]));
    LUT4 i23894_2_lut_rep_610_4_lut (.A(n2505[2]), .B(n2525[2]), .C(n31944), 
         .D(n31847), .Z(n31815)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i23894_2_lut_rep_610_4_lut.init = 16'hca00;
    PFUMX mux_845_i2 (.BLUT(n1742[1]), .ALUT(n1215[1]), .C0(n30165), .Z(pc_23__N_911[1]));
    LUT4 i1_2_lut_adj_455 (.A(addr_c[26]), .B(addr[27]), .Z(n18518)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_adj_455.init = 16'h8888;
    LUT4 i26315_2_lut_4_lut (.A(n2505[2]), .B(n2525[2]), .C(n31944), .D(n31847), 
         .Z(n28871)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i26315_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_4_lut_adj_456 (.A(n28412), .B(n28400), .C(addr[27]), .D(n31997), 
         .Z(n10467)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_456.init = 16'hffef;
    LUT4 i1_4_lut_adj_457 (.A(n28410), .B(\addr[19] ), .C(\addr[24] ), 
         .D(\addr[16] ), .Z(n28412)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_457.init = 16'hfffe;
    LUT4 i1_4_lut_adj_458 (.A(n28398), .B(\addr[12] ), .C(\addr[22] ), 
         .D(\addr[18] ), .Z(n28400)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_458.init = 16'hfffe;
    LUT4 i1_4_lut_adj_459 (.A(\addr[21] ), .B(\addr[13] ), .C(\addr[23] ), 
         .D(\addr[11] ), .Z(n28410)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_459.init = 16'hfffe;
    LUT4 i1_4_lut_adj_460 (.A(\addr[20] ), .B(\addr[17] ), .C(\addr[14] ), 
         .D(\addr[15] ), .Z(n28398)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_4_lut_adj_460.init = 16'hfffe;
    LUT4 i1_4_lut_adj_461 (.A(load_done_N_1741), .B(clk_c_enable_36), .C(n9710), 
         .D(n32026), .Z(address_ready)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(332[19:66])
    defparam i1_4_lut_adj_461.init = 16'h4000;
    PFUMX mux_845_i1 (.BLUT(n1742[0]), .ALUT(n1215[0]), .C0(n30165), .Z(pc_23__N_911[0]));
    LUT4 i1_2_lut_4_lut_adj_462 (.A(n2505[2]), .B(n2525[2]), .C(n31944), 
         .D(n33488), .Z(n28032)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_462.init = 16'hca00;
    LUT4 n14_bdd_2_lut_27983_2_lut_4_lut (.A(n2505[2]), .B(n2525[2]), .C(n31944), 
         .D(n31867), .Z(n30609)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam n14_bdd_2_lut_27983_2_lut_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_631_4_lut (.A(n2505[2]), .B(n2525[2]), .C(n31944), 
         .D(n31852), .Z(n31820)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_631_4_lut.init = 16'hffca;
    LUT4 mux_1832_i5_3_lut_rep_642 (.A(n2505[4]), .B(n2525[4]), .C(n31944), 
         .Z(n31847)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i5_3_lut_rep_642.init = 16'hcaca;
    LUT4 i23948_2_lut_rep_828 (.A(qv_data_write_n[1]), .B(qv_data_write_n[0]), 
         .Z(n32033)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23948_2_lut_rep_828.init = 16'h8888;
    LUT4 i1_2_lut_4_lut_adj_463 (.A(n2505[4]), .B(n2525[4]), .C(n31944), 
         .D(n31851), .Z(n26202)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_463.init = 16'h3500;
    LUT4 i1_2_lut_rep_600_4_lut (.A(n2505[4]), .B(n2525[4]), .C(n31944), 
         .D(n33488), .Z(n31805)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_600_4_lut.init = 16'hca00;
    LUT4 mux_1832_i12_3_lut_rep_643 (.A(n2505[11]), .B(n2525[11]), .C(n31944), 
         .Z(n31848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i12_3_lut_rep_643.init = 16'hcaca;
    LUT4 i1_2_lut_rep_666_3_lut (.A(qv_data_write_n[1]), .B(qv_data_write_n[0]), 
         .C(is_timer_addr), .Z(n31871)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_rep_666_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_635_3_lut_4_lut (.A(qv_data_write_n[1]), .B(qv_data_write_n[0]), 
         .C(\addr[2] ), .D(is_timer_addr), .Z(n31840)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;
    defparam i1_2_lut_rep_635_3_lut_4_lut.init = 16'h0700;
    LUT4 i27701_2_lut_rep_618_4_lut (.A(n2505[11]), .B(n2525[11]), .C(n31944), 
         .D(n31849), .Z(n31823)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i27701_2_lut_rep_618_4_lut.init = 16'h35ff;
    LUT4 mux_1832_i11_3_lut_rep_644 (.A(n2505[10]), .B(n2525[10]), .C(n31944), 
         .Z(n31849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i11_3_lut_rep_644.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_464 (.A(qv_data_write_n[1]), .B(qv_data_write_n[0]), 
         .C(data_ready_sync), .Z(n28444)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_464.init = 16'hf8f8;
    LUT4 i15381_2_lut_rep_829 (.A(\addr[4] ), .B(\addr[5] ), .Z(n32034)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15381_2_lut_rep_829.init = 16'heeee;
    LUT4 i102_2_lut_rep_731_3_lut_4_lut (.A(\addr[4] ), .B(\addr[5] ), .C(\addr[3] ), 
         .D(n32035), .Z(n31936)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i102_2_lut_rep_731_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_rep_830 (.A(addr[0]), .B(\addr[1] ), .Z(n32035)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_830.init = 16'heeee;
    LUT4 i1_2_lut_rep_757_3_lut (.A(addr[0]), .B(\addr[1] ), .C(\addr[5] ), 
         .Z(n31962)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_757_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_720_3_lut_4_lut (.A(addr[0]), .B(\addr[1] ), .C(\addr[4] ), 
         .D(\addr[5] ), .Z(n31925)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_720_3_lut_4_lut.init = 16'hefff;
    LUT4 i1_2_lut_rep_722_3_lut_4_lut (.A(addr[0]), .B(\addr[1] ), .C(\addr[4] ), 
         .D(\addr[5] ), .Z(n31927)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_rep_722_3_lut_4_lut.init = 16'hfeff;
    PFUMX mux_2123_i8 (.BLUT(n3340[7]), .ALUT(n5121[7]), .C0(n4281), .Z(n3458[7]));
    LUT4 i1_3_lut_rep_759_4_lut (.A(addr[0]), .B(\addr[1] ), .C(\addr[6] ), 
         .D(n26282), .Z(n31964)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_3_lut_rep_759_4_lut.init = 16'hfffe;
    LUT4 i27917_2_lut_rep_762_3_lut_4_lut (.A(addr[0]), .B(\addr[1] ), .C(\addr[5] ), 
         .D(\addr[4] ), .Z(n31967)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i27917_2_lut_rep_762_3_lut_4_lut.init = 16'h0001;
    PFUMX mux_2123_i6 (.BLUT(n3340[5]), .ALUT(n5121[5]), .C0(n4281), .Z(n3458[5]));
    LUT4 mux_1879_i4_4_lut (.A(n31807), .B(instr[18]), .C(n2810), .D(n31838), 
         .Z(n2630[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam mux_1879_i4_4_lut.init = 16'hca0a;
    LUT4 n14_bdd_2_lut_4_lut (.A(n2505[10]), .B(n2525[10]), .C(n31944), 
         .D(n31850), .Z(n30610)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam n14_bdd_2_lut_4_lut.init = 16'h3500;
    LUT4 i15599_2_lut_2_lut_4_lut (.A(n2505[10]), .B(n2525[10]), .C(n31944), 
         .D(n31735), .Z(n1720[3])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15599_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 i1_3_lut_adj_465 (.A(n31742), .B(rst_reg_n), .C(n31737), .Z(clk_c_enable_448)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(35[19:36])
    defparam i1_3_lut_adj_465.init = 16'hc8c8;
    LUT4 mux_1153_i1_3_lut (.A(n5[0]), .B(n31164), .C(n2138), .Z(n1764[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_1153_i1_3_lut.init = 16'hcaca;
    LUT4 i15576_2_lut_2_lut_4_lut (.A(n2505[10]), .B(n2525[10]), .C(n31944), 
         .D(n31860), .Z(n1725[3])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15576_2_lut_2_lut_4_lut.init = 16'hcaff;
    LUT4 i1_4_lut_adj_466 (.A(clk_c_enable_448), .B(n31742), .C(n27804), 
         .D(n31738), .Z(n2138)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_466.init = 16'ha888;
    LUT4 i1_4_lut_adj_467 (.A(n31744), .B(n24_adj_3162), .C(n9894), .D(n28898), 
         .Z(n27804)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_467.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_adj_468 (.A(n2505[10]), .B(n2525[10]), .C(n31944), 
         .D(n33488), .Z(n27726)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_468.init = 16'hca00;
    LUT4 mux_1832_i7_3_lut_rep_645 (.A(n2505[6]), .B(n2525[6]), .C(n31944), 
         .Z(n31850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i7_3_lut_rep_645.init = 16'hcaca;
    LUT4 i1_4_lut_adj_469 (.A(n824), .B(n31743), .C(address_ready), .D(is_load), 
         .Z(clk_c_enable_117)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_469.init = 16'hfeff;
    LUT4 i1_4_lut_adj_470 (.A(n824), .B(n31743), .C(is_load), .D(mem_op[0]), 
         .Z(n26972)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_4_lut_adj_470.init = 16'hffef;
    LUT4 mux_2101_i3_4_lut (.A(n29033), .B(n31863), .C(n4281), .D(n31764), 
         .Z(n3340[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2101_i3_4_lut.init = 16'hca0a;
    LUT4 i15449_2_lut_rep_619_4_lut (.A(n2505[6]), .B(n2525[6]), .C(n31944), 
         .D(n31851), .Z(n31824)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15449_2_lut_rep_619_4_lut.init = 16'hca00;
    LUT4 i243_2_lut (.A(data_ready_ext), .B(load_started), .Z(n824)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(297[17:47])
    defparam i243_2_lut.init = 16'h8888;
    LUT4 i15404_2_lut_4_lut (.A(n2505[6]), .B(n2525[6]), .C(n31944), .D(n31868), 
         .Z(n2982[4])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15404_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_2101_i4_4_lut (.A(n2152), .B(n31849), .C(n4281), .D(n31764), 
         .Z(n3340[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2101_i4_4_lut.init = 16'hca0a;
    LUT4 instr_6__I_0_127_i7_2_lut_rep_616_4_lut (.A(n2505[6]), .B(n2525[6]), 
         .C(n31944), .D(n31851), .Z(n31821)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_6__I_0_127_i7_2_lut_rep_616_4_lut.init = 16'hcaff;
    LUT4 i1_2_lut_rep_627_4_lut (.A(n2505[6]), .B(n2525[6]), .C(n31944), 
         .D(n31851), .Z(n7)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_627_4_lut.init = 16'hffca;
    LUT4 mux_1832_i6_3_lut_rep_646 (.A(n2505[5]), .B(n2525[5]), .C(n31944), 
         .Z(n31851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i6_3_lut_rep_646.init = 16'hcaca;
    LUT4 mux_1879_i1_4_lut (.A(n2602[0]), .B(n31868), .C(n2810), .D(n31838), 
         .Z(n2630[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam mux_1879_i1_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_rep_595_4_lut (.A(n2505[5]), .B(n2525[5]), .C(n31944), 
         .D(rst_reg_n), .Z(n31800)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_595_4_lut.init = 16'hca00;
    LUT4 i15412_3_lut (.A(n2804), .B(n2808), .C(n31864), .Z(n2621[0])) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(210[22] 212[16])
    defparam i15412_3_lut.init = 16'hc8c8;
    LUT4 mux_2119_i15_3_lut_4_lut (.A(n26), .B(n31722), .C(n3381[11]), 
         .D(n5223[13]), .Z(n3422[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_2119_i15_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_1832_i4_3_lut_rep_647 (.A(n2505[3]), .B(n2525[3]), .C(n31944), 
         .Z(n31852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i4_3_lut_rep_647.init = 16'hcaca;
    LUT4 mux_1822_i6_3_lut (.A(n21[5]), .B(n27[5]), .C(n2504), .Z(n2505[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i6_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_471 (.A(n2505[3]), .B(n2525[3]), .C(n31944), 
         .D(rst_reg_n), .Z(n28060)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_471.init = 16'hca00;
    LUT4 i27694_4_lut (.A(n31748), .B(rst_reg_n), .C(debug_ret), .D(n27680), 
         .Z(clk_c_enable_343)) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;
    defparam i27694_4_lut.init = 16'h3733;
    LUT4 i15397_2_lut_4_lut (.A(n2505[3]), .B(n2525[3]), .C(n31944), .D(n31868), 
         .Z(n2982[7])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15397_2_lut_4_lut.init = 16'hffca;
    LUT4 mux_1832_i13_3_lut_rep_648 (.A(n2505[12]), .B(n2525[12]), .C(n31944), 
         .Z(n31853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i13_3_lut_rep_648.init = 16'hcaca;
    LUT4 mux_1826_i6_3_lut (.A(n31[5]), .B(n6[5]), .C(n2524), .Z(n2525[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i6_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_472 (.A(n2505[12]), .B(n2525[12]), .C(n31944), 
         .D(additional_mem_ops_2__N_1132[0]), .Z(n4_adj_3163)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_472.init = 16'h00ca;
    LUT4 i1_2_lut_4_lut_adj_473 (.A(n2505[12]), .B(n2525[12]), .C(n31944), 
         .D(n31867), .Z(n28366)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_473.init = 16'hca00;
    LUT4 equal_25_i3_2_lut_4_lut (.A(n2505[12]), .B(n2525[12]), .C(n31944), 
         .D(n31867), .Z(n3)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam equal_25_i3_2_lut_4_lut.init = 16'hff35;
    LUT4 i15703_4_lut (.A(n31849), .B(n31845), .C(n31851), .D(n31860), 
         .Z(n3304[3])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15703_4_lut.init = 16'hc088;
    LUT4 i15704_4_lut (.A(n31848), .B(n31845), .C(n31850), .D(n31860), 
         .Z(n3304[4])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15704_4_lut.init = 16'hc088;
    LUT4 i1_2_lut_rep_524_4_lut (.A(n31744), .B(n31738), .C(n9894), .D(n31742), 
         .Z(clk_c_enable_30)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_524_4_lut.init = 16'h0004;
    LUT4 i1_4_lut_adj_474 (.A(n31748), .B(n28152), .C(n28156), .D(n8), 
         .Z(clk_c_enable_370)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_474.init = 16'hfafe;
    L6MUX21 shift_right_317_i272 (.D0(n29193), .D1(n10899), .SD(n29318), 
            .Z(debug_branch_N_840[31])) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i15705_4_lut (.A(n31846), .B(n31845), .C(n31853), .D(n31860), 
         .Z(n3304[5])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15705_4_lut.init = 16'hc088;
    PFUMX i27984 (.BLUT(n30610), .ALUT(n30609), .C0(n4269), .Z(n30611));
    LUT4 i15706_4_lut (.A(n31851), .B(n31845), .C(n31846), .D(n31860), 
         .Z(n3304[6])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15706_4_lut.init = 16'hc088;
    LUT4 i1_4_lut_adj_475 (.A(n32017), .B(n27214), .C(n32034), .D(n18518), 
         .Z(is_timer_addr)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_475.init = 16'h0400;
    LUT4 i1_4_lut_adj_476 (.A(\addr[3] ), .B(n28496), .C(n28498), .D(n28494), 
         .Z(n27214)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_476.init = 16'h4000;
    LUT4 i1_4_lut_adj_477 (.A(\addr[23] ), .B(n28486), .C(n28474), .D(addr_c[25]), 
         .Z(n28496)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_477.init = 16'h8000;
    LUT4 i1_4_lut_adj_478 (.A(\addr[12] ), .B(n28492), .C(n28480), .D(\addr[11] ), 
         .Z(n28498)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_478.init = 16'h8000;
    LUT4 i1_4_lut_adj_479 (.A(\addr[10] ), .B(\addr[20] ), .C(\addr[24] ), 
         .D(\addr[15] ), .Z(n28494)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_479.init = 16'h8000;
    LUT4 i1_2_lut_adj_480 (.A(\addr[9] ), .B(\addr[8] ), .Z(n28486)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_480.init = 16'h8888;
    LUT4 i1_2_lut_adj_481 (.A(\addr[16] ), .B(\addr[13] ), .Z(n28474)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_481.init = 16'h8888;
    LUT4 i1_4_lut_adj_482 (.A(\addr[17] ), .B(\addr[14] ), .C(\addr[19] ), 
         .D(\addr[21] ), .Z(n28492)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_482.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_483 (.A(n31744), .B(n31738), .C(n9894), .D(n26993), 
         .Z(clk_c_enable_358)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_483.init = 16'h0004;
    LUT4 n31199_bdd_3_lut_4_lut (.A(n31796), .B(n31852), .C(n31860), .D(n31198), 
         .Z(n31200)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam n31199_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_adj_484 (.A(\addr[22] ), .B(\addr[18] ), .Z(n28480)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_484.init = 16'h8888;
    LUT4 i1_2_lut_adj_485 (.A(\addr[2] ), .B(\addr[3] ), .Z(n26266)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_485.init = 16'hbbbb;
    PFUMX i29 (.BLUT(n29192), .ALUT(n29194), .C0(n31937), .Z(n10899));
    LUT4 mux_2096_i7_4_lut (.A(n2602[0]), .B(n31851), .C(n4271), .D(n31868), 
         .Z(n3271[6])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2096_i7_4_lut.init = 16'hfaca;
    LUT4 i15707_4_lut (.A(n31850), .B(n31845), .C(n31852), .D(n31860), 
         .Z(n3304[7])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15707_4_lut.init = 16'hc088;
    LUT4 mux_2138_i9_4_lut (.A(n3381[8]), .B(instr[28]), .C(n4285), .D(n31728), 
         .Z(n3505[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2138_i9_4_lut.init = 16'hca0a;
    LUT4 i21203_1_lut (.A(counter_hi[2]), .Z(c_2__N_1861[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i21203_1_lut.init = 16'h5555;
    LUT4 mux_2084_i4_4_lut (.A(n31851), .B(n27734), .C(n31719), .D(n31738), 
         .Z(n3195[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2084_i4_4_lut.init = 16'hca0a;
    LUT4 mux_2084_i7_4_lut (.A(n31864), .B(n27744), .C(n31719), .D(n31738), 
         .Z(n3195[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2084_i7_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_4_lut_adj_486 (.A(n29025), .B(n29043), .C(n31944), .D(n33488), 
         .Z(n28098)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_486.init = 16'hca00;
    LUT4 mux_1832_i2_3_lut_rep_655 (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .Z(n31860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i2_3_lut_rep_655.init = 16'hcaca;
    LUT4 i23859_2_lut_rep_580_3_lut_2_lut_4_lut (.A(n2505[1]), .B(n2525[1]), 
         .C(n31944), .D(n31869), .Z(n31785)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i23859_2_lut_rep_580_3_lut_2_lut_4_lut.init = 16'h35ca;
    LUT4 instr_1__bdd_2_lut_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .D(n31864), .Z(n31163)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam instr_1__bdd_2_lut_4_lut.init = 16'hffca;
    PFUMX i26532 (.BLUT(n29148), .ALUT(n227), .C0(counter_hi[4]), .Z(n29149));
    LUT4 i1_3_lut_rep_653_4_lut (.A(n32033), .B(n31905), .C(\addr[2] ), 
         .D(n31936), .Z(clk_c_enable_390)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_3_lut_rep_653_4_lut.init = 16'h0004;
    LUT4 i4439_2_lut_rep_837 (.A(\pc[1] ), .B(instr_len[1]), .Z(n32042)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i4439_2_lut_rep_837.init = 16'h6666;
    LUT4 i1_4_lut_4_lut_adj_487 (.A(\pc[1] ), .B(instr_len[1]), .C(debug_instr_valid), 
         .D(\instr_addr_23__N_318[0] ), .Z(n10112)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_4_lut_4_lut_adj_487.init = 16'h956a;
    LUT4 i1_2_lut_rep_604_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .D(n31869), .Z(n31809)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_604_4_lut.init = 16'h3500;
    L6MUX21 i27041 (.D0(n29656), .D1(n29657), .SD(counter_hi[3]), .Z(n29658));
    PFUMX i48 (.BLUT(n12_adj_3164), .ALUT(n30_adj_3165), .C0(n31860), 
          .Z(n43));
    LUT4 i26518_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), .C(counter_hi[2]), 
         .D(\next_pc_for_core[5] ), .Z(n29135)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i26518_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_2119_i8_3_lut (.A(n3271[7]), .B(n3304[7]), .C(n4279), .Z(n3422[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2119_i8_3_lut.init = 16'hcaca;
    LUT4 i4581_2_lut_rep_760_3_lut (.A(\pc[1] ), .B(instr_len[1]), .C(\instr_addr_23__N_318[0] ), 
         .Z(n31965)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i4581_2_lut_rep_760_3_lut.init = 16'hf9f9;
    LUT4 mux_347_i1_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), .C(debug_ret), 
         .D(return_addr[1]), .Z(n34[0])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam mux_347_i1_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i27120 (.D0(n29733), .D1(n29734), .SD(counter_hi[2]), .Z(n29737));
    LUT4 i15263_1_lut_rep_584_2_lut_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .D(n31869), .Z(n31789)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15263_1_lut_rep_584_2_lut_4_lut.init = 16'h35ff;
    LUT4 i1_3_lut_rep_563 (.A(is_timer_addr), .B(data_ready_ext), .C(data_ready_latch), 
         .Z(n31768)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(258[53:106])
    defparam i1_3_lut_rep_563.init = 16'hfefe;
    PFUMX i26520 (.BLUT(n29136), .ALUT(n226), .C0(n33484), .Z(n29137));
    LUT4 i5711_2_lut_4_lut (.A(is_timer_addr), .B(data_ready_ext), .C(data_ready_latch), 
         .D(load_done_N_1741), .Z(n8289)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(258[53:106])
    defparam i5711_2_lut_4_lut.init = 16'hfe00;
    LUT4 i2_2_lut_rep_626_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .D(n31869), .Z(n31831)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i2_2_lut_rep_626_4_lut.init = 16'h00ca;
    LUT4 i15544_3_lut_4_lut (.A(n31790), .B(n31845), .C(n31868), .D(n31867), 
         .Z(n29)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (D)))) */ ;
    defparam i15544_3_lut_4_lut.init = 16'h001f;
    LUT4 i15574_2_lut_2_lut_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .D(n31865), .Z(n1725[1])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15574_2_lut_2_lut_4_lut.init = 16'h3500;
    LUT4 i15575_2_lut_2_lut_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .D(n31863), .Z(n1725[2])) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15575_2_lut_2_lut_4_lut.init = 16'h3500;
    LUT4 gnd_bdd_2_lut_28463_2_lut_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .D(n31437), .Z(n31438)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam gnd_bdd_2_lut_28463_2_lut_4_lut.init = 16'h3500;
    L6MUX21 i27039 (.D0(n29652), .D1(n29653), .SD(counter_hi[2]), .Z(n29656));
    LUT4 i27926_2_lut_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), .D(n31868), 
         .Z(n29293)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i27926_2_lut_4_lut.init = 16'hcaff;
    L6MUX21 i27040 (.D0(n29654), .D1(n29655), .SD(counter_hi[2]), .Z(n29657));
    L6MUX21 i27046 (.D0(n29659), .D1(n29660), .SD(counter_hi[2]), .Z(n29663));
    LUT4 i4419_3_lut_4_lut (.A(rd_c[1]), .B(rd[0]), .C(rd_c[2]), .D(rd_c[3]), 
         .Z(n108[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(180[19:31])
    defparam i4419_3_lut_4_lut.init = 16'h7f80;
    LUT4 i1_3_lut_4_lut_adj_488 (.A(rd_c[1]), .B(rd[0]), .C(n32046), .D(rd_c[2]), 
         .Z(n28222)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)))+!A !(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(180[19:31])
    defparam i1_3_lut_4_lut_adj_488.init = 16'h7080;
    LUT4 i1_3_lut_rep_841 (.A(additional_mem_ops[1]), .B(additional_mem_ops[0]), 
         .C(additional_mem_ops[2]), .Z(n32046)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_3_lut_rep_841.init = 16'hfefe;
    PFUMX next_pc_for_core_23__I_0_i209 (.BLUT(n149), .ALUT(n225_adj_3166), 
          .C0(counter_hi[4]), .Z(n209)) /* synthesis LSE_LINE_FILE_ID=16, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=94, LSE_RLINE=130 */ ;
    LUT4 i1_2_lut_4_lut_adj_489 (.A(additional_mem_ops[1]), .B(additional_mem_ops[0]), 
         .C(additional_mem_ops[2]), .D(n33488), .Z(n28204)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(159[12] 214[8])
    defparam i1_2_lut_4_lut_adj_489.init = 16'hfe00;
    LUT4 i1_4_lut_adj_490 (.A(n2808), .B(n31722), .C(n31863), .D(n4_adj_3136), 
         .Z(n26829)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;
    defparam i1_4_lut_adj_490.init = 16'h20a0;
    LUT4 i15262_2_lut_rep_633_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .D(n31869), .Z(n31838)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15262_2_lut_rep_633_4_lut.init = 16'hca00;
    LUT4 i27770_2_lut_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), .D(n31869), 
         .Z(n29215)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i27770_2_lut_4_lut.init = 16'hffca;
    LUT4 i166_2_lut_rep_613_4_lut (.A(n2505[1]), .B(n2525[1]), .C(n31944), 
         .D(n31869), .Z(n31818)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i166_2_lut_rep_613_4_lut.init = 16'h3500;
    LUT4 i1_4_lut_adj_491 (.A(addr_out[3]), .B(n31898), .C(addr_offset[3]), 
         .D(addr_offset[2]), .Z(n27068)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(121[15:26])
    defparam i1_4_lut_adj_491.init = 16'h965a;
    PFUMX i27117 (.BLUT(\mem_data_from_read[7] ), .ALUT(\data_from_read[7] ), 
          .C0(n30171), .Z(n29734));
    LUT4 mux_1538_i5_3_lut_rep_656 (.A(n29023), .B(n29041), .C(n31944), 
         .Z(n31861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1538_i5_3_lut_rep_656.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_492 (.A(n29023), .B(n29041), .C(n31944), .D(n33488), 
         .Z(n28110)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_492.init = 16'hca00;
    LUT4 i15268_3_lut (.A(n32046), .B(rst_reg_n), .C(n31740), .Z(data_continue_N_963)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i15268_3_lut.init = 16'ha8a8;
    LUT4 no_write_in_progress_I_42_4_lut (.A(n28444), .B(addr_out[27]), 
         .C(n31903), .D(data_ready_ext), .Z(no_write_in_progress_N_471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(279[18] 289[12])
    defparam no_write_in_progress_I_42_4_lut.init = 16'hcfca;
    LUT4 i1_3_lut_adj_493 (.A(n31744), .B(n31742), .C(n9894), .Z(n27846)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_493.init = 16'hfefe;
    PFUMX i27116 (.BLUT(\mem_data_from_read[3] ), .ALUT(\data_from_read[3] ), 
          .C0(n30170), .Z(n29733));
    LUT4 i21208_2_lut_rep_844 (.A(counter_hi[3]), .B(counter_hi[2]), .Z(n32049)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i21208_2_lut_rep_844.init = 16'h8888;
    LUT4 i15260_4_lut (.A(instr_fetch_running_N_943), .B(rst_reg_n), .C(was_early_branch), 
         .D(n31748), .Z(n6411)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(385[12] 432[8])
    defparam i15260_4_lut.init = 16'hc088;
    LUT4 i15665_2_lut_3_lut_4_lut_3_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(counter_hi[4]), .Z(csr_read_3__N_1443[0])) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i15665_2_lut_3_lut_4_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 i1_3_lut_4_lut_adj_494 (.A(n33486), .B(counter_hi[2]), .C(debug_instr_valid), 
         .D(n33484), .Z(n27018)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i1_3_lut_4_lut_adj_494.init = 16'hf7ff;
    LUT4 i21212_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(counter_hi[4]), 
         .Z(n36[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i21212_2_lut_3_lut.init = 16'h7878;
    LUT4 i13_3_lut_4_lut_rep_835_3_lut (.A(counter_hi[3]), .B(counter_hi[2]), 
         .C(counter_hi[4]), .Z(n32040)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i13_3_lut_4_lut_rep_835_3_lut.init = 16'h8181;
    PFUMX i26945 (.BLUT(n29558), .ALUT(n29559), .C0(counter_hi[3]), .Z(n29562));
    LUT4 i4370_2_lut_rep_845 (.A(rs2[0]), .B(mem_op_increment_reg), .Z(n32050)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i4370_2_lut_rep_845.init = 16'h8888;
    LUT4 i4378_2_lut_rep_770_3_lut (.A(rs2[0]), .B(mem_op_increment_reg), 
         .C(rs2[1]), .Z(n31975)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i4378_2_lut_rep_770_3_lut.init = 16'h8080;
    LUT4 i4385_2_lut_3_lut_4_lut (.A(rs2[0]), .B(mem_op_increment_reg), 
         .C(rs2[2]), .D(rs2[1]), .Z(n6668)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(179[20:56])
    defparam i4385_2_lut_3_lut_4_lut.init = 16'h8000;
    PFUMX i27035 (.BLUT(\mem_data_from_read[0] ), .ALUT(\data_from_read[0] ), 
          .C0(n30170), .Z(n29652));
    PFUMX i26946 (.BLUT(n29560), .ALUT(n29561), .C0(counter_hi[3]), .Z(n29563));
    PFUMX i27036 (.BLUT(\mem_data_from_read[4] ), .ALUT(\data_from_read[4] ), 
          .C0(n31958), .Z(n29653));
    PFUMX i27037 (.BLUT(\mem_data_from_read[8] ), .ALUT(\data_from_read[8] ), 
          .C0(n30171), .Z(n29654));
    PFUMX i26952 (.BLUT(n29565), .ALUT(n29566), .C0(counter_hi[3]), .Z(n29569));
    LUT4 pc_23__I_0_450_i269_3_lut (.A(n209_adj_3151), .B(data_rs1[0]), 
         .C(alu_a_in_3__N_1552), .Z(debug_branch_N_442[28])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam pc_23__I_0_450_i269_3_lut.init = 16'hacac;
    LUT4 mux_2119_i5_3_lut (.A(n3271[4]), .B(n3304[4]), .C(n4279), .Z(n3422[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2119_i5_3_lut.init = 16'hcaca;
    PFUMX i27038 (.BLUT(\mem_data_from_read[12] ), .ALUT(\data_from_read[12] ), 
          .C0(n30171), .Z(n29655));
    LUT4 mux_1832_i10_3_lut_rep_658 (.A(n2505[9]), .B(n2525[9]), .C(n31944), 
         .Z(n31863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i10_3_lut_rep_658.init = 16'hcaca;
    LUT4 i1_2_lut_rep_632_4_lut (.A(n2505[9]), .B(n2525[9]), .C(n31944), 
         .D(n31864), .Z(n31837)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_632_4_lut.init = 16'hffca;
    LUT4 i15598_2_lut_2_lut_4_lut (.A(n2505[9]), .B(n2525[9]), .C(n31944), 
         .D(n31735), .Z(n1720[2])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15598_2_lut_2_lut_4_lut.init = 16'h00ca;
    PFUMX i27042 (.BLUT(\mem_data_from_read[1] ), .ALUT(\data_from_read[1] ), 
          .C0(n31958), .Z(n29659));
    PFUMX i27043 (.BLUT(\mem_data_from_read[5] ), .ALUT(\data_from_read[5] ), 
          .C0(n30171), .Z(n29660));
    LUT4 mux_1832_i9_3_lut_rep_660 (.A(n2505[8]), .B(n2525[8]), .C(n31944), 
         .Z(n31865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i9_3_lut_rep_660.init = 16'hcaca;
    LUT4 pc_23__I_0_450_i157_3_lut (.A(\pc[8] ), .B(\pc[12] ), .C(counter_hi[2]), 
         .Z(n157_adj_3152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(350[15:27])
    defparam pc_23__I_0_450_i157_3_lut.init = 16'hcaca;
    LUT4 i27752_2_lut_3_lut_4_lut (.A(n31741), .B(n31748), .C(rst_reg_n), 
         .D(n27846), .Z(clk_c_enable_214)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i27752_2_lut_3_lut_4_lut.init = 16'h0fef;
    PFUMX i38 (.BLUT(n17_adj_3142), .ALUT(n22_adj_3167), .C0(n31868), 
          .Z(n24_adj_3162));
    LUT4 i15597_2_lut_2_lut_4_lut (.A(n2505[8]), .B(n2525[8]), .C(n31944), 
         .D(n31735), .Z(n1720[1])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15597_2_lut_2_lut_4_lut.init = 16'h00ca;
    LUT4 i15601_2_lut_4_lut (.A(n2505[8]), .B(n2525[8]), .C(n31944), .D(n2804), 
         .Z(n2597[1])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15601_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_3_lut_rep_532_4_lut (.A(n31741), .B(n31748), .C(n9894), .D(n31744), 
         .Z(n31737)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(186[22:86])
    defparam i1_3_lut_rep_532_4_lut.init = 16'h000e;
    PFUMX i26953 (.BLUT(n29567), .ALUT(n29568), .C0(counter_hi[3]), .Z(n29570));
    LUT4 mux_2138_i11_4_lut (.A(n2982[13]), .B(instr[30]), .C(n4285), 
         .D(n31728), .Z(n3505[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2138_i11_4_lut.init = 16'hca0a;
    LUT4 mux_1832_i14_3_lut_rep_662 (.A(n2505[13]), .B(n2525[13]), .C(n31944), 
         .Z(n31867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i14_3_lut_rep_662.init = 16'hcaca;
    LUT4 i15787_2_lut_4_lut (.A(n2505[13]), .B(n2525[13]), .C(n31944), 
         .D(additional_mem_ops_2__N_1132[0]), .Z(mem_op_2__N_1114[1])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15787_2_lut_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_rep_599_4_lut (.A(n2505[13]), .B(n2525[13]), .C(n31944), 
         .D(n31869), .Z(n31804)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_599_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_rep_849 (.A(\instr_len[2] ), .B(\pc[2] ), .Z(n32054)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_2_lut_rep_849.init = 16'h6666;
    LUT4 mux_2138_i13_3_lut (.A(n3271[13]), .B(n3422[12]), .C(n29428), 
         .Z(n3505[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2138_i13_3_lut.init = 16'hcaca;
    LUT4 i15228_2_lut_rep_601_4_lut (.A(n2505[13]), .B(n2525[13]), .C(n31944), 
         .D(n31869), .Z(n31806)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i15228_2_lut_rep_601_4_lut.init = 16'hffca;
    LUT4 i224_2_lut_rep_614_3_lut_4_lut (.A(n32033), .B(n31905), .C(n31932), 
         .D(n31922), .Z(n31819)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i224_2_lut_rep_614_3_lut_4_lut.init = 16'h0004;
    PFUMX i26959 (.BLUT(n29572), .ALUT(n29573), .C0(counter_hi[3]), .Z(n29576));
    PFUMX i54 (.BLUT(n37), .ALUT(n32_adj_3168), .C0(n29293), .Z(n35));
    LUT4 i1_2_lut_3_lut_adj_495 (.A(\instr_len[2] ), .B(\pc[2] ), .C(instr_addr_23__N_318[1]), 
         .Z(n28284)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1_2_lut_3_lut_adj_495.init = 16'h9696;
    LUT4 i1_4_lut_adj_496 (.A(n824), .B(n31743), .C(is_load), .D(mem_op[1]), 
         .Z(n26971)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_4_lut_adj_496.init = 16'hffef;
    LUT4 mux_2138_i14_3_lut (.A(n3271[13]), .B(n3422[13]), .C(n29428), 
         .Z(n3505[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2138_i14_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_629_4_lut (.A(n2505[13]), .B(n2525[13]), .C(n31944), 
         .D(n31868), .Z(n31834)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_629_4_lut.init = 16'h00ca;
    LUT4 mux_2138_i15_3_lut (.A(n3271[13]), .B(n3422[14]), .C(n29428), 
         .Z(n3505[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2138_i15_3_lut.init = 16'hcaca;
    PFUMX i42 (.BLUT(n10), .ALUT(n29), .C0(n31869), .Z(n23));
    LUT4 i1842_3_lut_rep_739_4_lut_4_lut (.A(\instr_len[2] ), .B(\pc[2] ), 
         .C(debug_instr_valid), .D(n32055), .Z(n31944)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C (D))+!B !(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i1842_3_lut_rep_739_4_lut_4_lut.init = 16'h9c6c;
    LUT4 mux_1832_i16_3_lut_rep_663 (.A(n2505[15]), .B(n2525[15]), .C(n31944), 
         .Z(n31868)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i16_3_lut_rep_663.init = 16'hcaca;
    PFUMX i26960 (.BLUT(n29574), .ALUT(n29575), .C0(counter_hi[3]), .Z(n29577));
    LUT4 i4441_2_lut_rep_850 (.A(\pc[1] ), .B(instr_len[1]), .Z(n32055)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i4441_2_lut_rep_850.init = 16'h8888;
    LUT4 i2_2_lut_rep_773_3_lut_4_lut (.A(\pc[1] ), .B(instr_len[1]), .C(\pc[2] ), 
         .D(\instr_len[2] ), .Z(n31978)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(155[33:70])
    defparam i2_2_lut_rep_773_3_lut_4_lut.init = 16'h8778;
    PFUMX i26543 (.BLUT(\mem_data_from_read[24] ), .ALUT(\mem_data_from_read[28] ), 
          .C0(counter_hi[2]), .Z(n29160));
    PFUMX i26549 (.BLUT(\mem_data_from_read[25] ), .ALUT(\mem_data_from_read[29] ), 
          .C0(counter_hi[2]), .Z(n29166));
    LUT4 data_from_read_11__bdd_3_lut_then_3_lut (.A(n31879), .B(n19), .C(n31885), 
         .Z(n32065)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam data_from_read_11__bdd_3_lut_then_3_lut.init = 16'hcece;
    LUT4 data_from_read_11__bdd_3_lut_else_3_lut (.A(n31879), .B(n19), .C(\peri_data_out[11] ), 
         .D(n4), .Z(n32064)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam data_from_read_11__bdd_3_lut_else_3_lut.init = 16'heeec;
    PFUMX i26981 (.BLUT(n29594), .ALUT(n29595), .C0(counter_hi[3]), .Z(n29598));
    LUT4 i1_2_lut_rep_617_4_lut (.A(n2505[15]), .B(n2525[15]), .C(n31944), 
         .D(n31869), .Z(n31822)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_617_4_lut.init = 16'h00ca;
    LUT4 i1_2_lut_2_lut_4_lut (.A(n2505[15]), .B(n2525[15]), .C(n31944), 
         .D(n31869), .Z(n12_adj_3164)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_2_lut_4_lut.init = 16'h3500;
    LUT4 i27650_2_lut_rep_607_4_lut (.A(n2505[15]), .B(n2525[15]), .C(n31944), 
         .D(n31869), .Z(n31812)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+(D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i27650_2_lut_rep_607_4_lut.init = 16'h0035;
    LUT4 i1_2_lut_rep_628_4_lut (.A(n2505[15]), .B(n2525[15]), .C(n31944), 
         .D(n31869), .Z(n31833)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_rep_628_4_lut.init = 16'hca00;
    LUT4 i1_2_lut_4_lut_adj_497 (.A(n2505[15]), .B(n2525[15]), .C(n31944), 
         .D(n33488), .Z(n27688)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i1_2_lut_4_lut_adj_497.init = 16'hca00;
    PFUMX i26573 (.BLUT(\mem_data_from_read[26] ), .ALUT(\mem_data_from_read[30] ), 
          .C0(counter_hi[2]), .Z(n29190));
    LUT4 mux_2138_i16_3_lut (.A(n3271[13]), .B(n3422[15]), .C(n29428), 
         .Z(n3505[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2138_i16_3_lut.init = 16'hcaca;
    LUT4 mux_1832_i1_3_lut_rep_664 (.A(n2505[0]), .B(n2525[0]), .C(n31944), 
         .Z(n31869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1832_i1_3_lut_rep_664.init = 16'hcaca;
    LUT4 i4977_1_lut_rep_630_3_lut (.A(n2505[0]), .B(n2525[0]), .C(n31944), 
         .Z(n31835)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam i4977_1_lut_rep_630_3_lut.init = 16'h3535;
    PFUMX i26576 (.BLUT(\mem_data_from_read[27] ), .ALUT(\mem_data_from_read[31] ), 
          .C0(counter_hi[2]), .Z(n29193));
    LUT4 i1_3_lut_3_lut_adj_498 (.A(n31742), .B(n4322[0]), .C(n4322[1]), 
         .Z(n4_adj_3169)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i1_3_lut_3_lut_adj_498.init = 16'hfdfd;
    LUT4 i27659_4_lut (.A(n31748), .B(n31744), .C(n9894), .D(is_ret_de), 
         .Z(debug_instr_valid_N_436)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i27659_4_lut.init = 16'h0001;
    PFUMX i28152 (.BLUT(n33493), .ALUT(n30950), .C0(n31718), .Z(n3505[17]));
    PFUMX i38_adj_499 (.BLUT(n24_adj_3140), .ALUT(n17), .C0(n31860), .Z(n22_adj_3135));
    LUT4 i1_3_lut_adj_500 (.A(n4322[1]), .B(n4322[0]), .C(n31742), .Z(additional_mem_ops_2__N_749[1])) /* synthesis lut_function=(A (B+!(C))+!A !(B+!(C))) */ ;
    defparam i1_3_lut_adj_500.init = 16'h9a9a;
    LUT4 i27834_4_lut (.A(counter_hi[2]), .B(n31966), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(clk_c_enable_173)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(307[12] 313[8])
    defparam i27834_4_lut.init = 16'h0080;
    LUT4 i1_3_lut_adj_501 (.A(is_jal_de), .B(rst_reg_n), .C(is_ret_de), 
         .Z(n28150)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut_adj_501.init = 16'hc8c8;
    LUT4 i15455_2_lut (.A(n30611), .B(n4277), .Z(n3381[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam i15455_2_lut.init = 16'h8888;
    LUT4 n3301_bdd_4_lut (.A(n31714), .B(n4277), .C(n26656), .D(n31850), 
         .Z(n30707)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (C))) */ ;
    defparam n3301_bdd_4_lut.init = 16'he2c0;
    LUT4 i16_4_lut_adj_502 (.A(n4285), .B(clk_c_enable_30), .C(rst_reg_n), 
         .D(n26899), .Z(clk_c_enable_221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i16_4_lut_adj_502.init = 16'hcfca;
    LUT4 i1_4_lut_adj_503 (.A(n31744), .B(n31738), .C(n31742), .D(n28008), 
         .Z(n26899)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_503.init = 16'h0400;
    LUT4 i1_4_lut_adj_504 (.A(n26), .B(n28006), .C(n35), .D(n22), .Z(n28008)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_504.init = 16'hccc8;
    LUT4 mux_2147_i7_3_lut (.A(n3505[6]), .B(n3458[6]), .C(n4285), .Z(n3546[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i7_3_lut.init = 16'hcaca;
    LUT4 mux_2147_i6_3_lut (.A(n3505[5]), .B(n3458[5]), .C(n4285), .Z(n3546[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i6_3_lut.init = 16'hcaca;
    LUT4 mux_2147_i4_3_lut (.A(n3505[3]), .B(n3458[3]), .C(n4285), .Z(n3546[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i4_3_lut.init = 16'hcaca;
    LUT4 mux_2147_i2_3_lut (.A(n3505[1]), .B(n31121), .C(n4285), .Z(n3546[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2147_i2_3_lut.init = 16'hcaca;
    PFUMX i26982 (.BLUT(n29596), .ALUT(n29597), .C0(counter_hi[3]), .Z(n29599));
    LUT4 i1_2_lut_3_lut_4_lut_adj_505 (.A(n31860), .B(n31806), .C(n31800), 
         .D(n31845), .Z(n27738)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_505.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_506 (.A(n31860), .B(n31806), .C(n27726), 
         .D(n31845), .Z(n27728)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_506.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_507 (.A(instr_addr_23__N_318[1]), .B(n31910), 
         .C(n1), .D(\pc[2] ), .Z(n27606)) /* synthesis lut_function=(A (B (C+(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i1_2_lut_3_lut_4_lut_adj_507.init = 16'hf9f6;
    LUT4 mux_346_i2_3_lut_4_lut (.A(instr_addr_23__N_318[1]), .B(n31910), 
         .C(debug_ret), .D(return_addr[2]), .Z(n1764_adj_3181[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam mux_346_i2_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_1822_i7_3_lut (.A(n21[6]), .B(n27[6]), .C(n2504), .Z(n2505[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1826_i7_3_lut (.A(n31[6]), .B(n6[6]), .C(n2524), .Z(n2525[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i7_3_lut.init = 16'hcaca;
    LUT4 mux_1822_i11_3_lut (.A(n21[10]), .B(n27[10]), .C(n2504), .Z(n2505[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i11_3_lut.init = 16'hcaca;
    LUT4 mux_2096_i9_3_lut_4_lut (.A(n31853), .B(n31808), .C(n4279), .D(n2602[2]), 
         .Z(n3271[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2096_i9_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_1826_i11_3_lut (.A(n31[10]), .B(n6[10]), .C(n2524), .Z(n2525[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i11_3_lut.init = 16'hcaca;
    LUT4 n30949_bdd_3_lut_4_lut (.A(n31853), .B(n31808), .C(n4279), .D(n30949), 
         .Z(n30950)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n30949_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2096_i17_3_lut_4_lut (.A(n31853), .B(n31808), .C(n4279), 
         .D(n2982[16]), .Z(n3271[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2096_i17_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_1822_i12_3_lut (.A(n21[11]), .B(n27[11]), .C(n2504), .Z(n2505[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i12_3_lut.init = 16'hcaca;
    LUT4 n30836_bdd_3_lut_28546_4_lut (.A(n31853), .B(n31808), .C(n4279), 
         .D(n30836), .Z(n30837)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n30836_bdd_3_lut_28546_4_lut.init = 16'h8f80;
    LUT4 mux_1826_i12_3_lut (.A(n31[11]), .B(n6[11]), .C(n2524), .Z(n2525[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i12_3_lut.init = 16'hcaca;
    LUT4 pc_3__bdd_3_lut_28046 (.A(\pc[7] ), .B(\pc[15] ), .C(counter_hi[3]), 
         .Z(n30742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_3__bdd_3_lut_28046.init = 16'hcaca;
    LUT4 mux_2096_i14_3_lut_4_lut (.A(n31853), .B(n31808), .C(n4279), 
         .D(n2982[13]), .Z(n3271[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2096_i14_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_1822_i5_3_lut (.A(n21[4]), .B(n27[4]), .C(n2504), .Z(n2505[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i5_3_lut.init = 16'hcaca;
    LUT4 mux_1826_i5_3_lut (.A(n31[4]), .B(n6[4]), .C(n2524), .Z(n2525[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i5_3_lut.init = 16'hcaca;
    LUT4 i27673_4_lut (.A(n31748), .B(debug_ret), .C(n31942), .D(n27978), 
         .Z(clk_c_enable_287)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i27673_4_lut.init = 16'h0010;
    PFUMX i29_adj_508 (.BLUT(n20_adj_3144), .ALUT(n13_adj_3146), .C0(n31845), 
          .Z(n16_adj_3171));
    LUT4 mux_1822_i3_3_lut (.A(n21[2]), .B(n27[2]), .C(n2504), .Z(n2505[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i3_3_lut.init = 16'hcaca;
    LUT4 mux_1826_i3_3_lut (.A(n31[2]), .B(n6[2]), .C(n2524), .Z(n2525[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i3_3_lut.init = 16'hcaca;
    LUT4 i43_3_lut_4_lut (.A(n31812), .B(n31817), .C(n31860), .D(n23), 
         .Z(n26_adj_3172)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam i43_3_lut_4_lut.init = 16'h2f20;
    PFUMX i29_adj_509 (.BLUT(n9_c), .ALUT(n12_c), .C0(debug_instr_valid), 
          .Z(n16));
    LUT4 mux_1532_i11_3_lut (.A(n6[10]), .B(n21[10]), .C(n2524), .Z(n2163[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i11_3_lut.init = 16'hcaca;
    LUT4 mux_1528_i11_rep_105_3_lut (.A(n27[10]), .B(n31[10]), .C(n2504), 
         .Z(n29051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i11_rep_105_3_lut.init = 16'hcaca;
    LUT4 mux_2101_i16_3_lut_4_lut (.A(instr[31]), .B(n31838), .C(n31733), 
         .D(n5081[8]), .Z(n3340[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2101_i16_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_2101_i13_3_lut_4_lut (.A(instr[31]), .B(n31838), .C(n31733), 
         .D(n5081[5]), .Z(n3340[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2101_i13_3_lut_4_lut.init = 16'hf808;
    LUT4 n13_bdd_3_lut_28389 (.A(\mem_data_from_read[18] ), .B(\mem_data_from_read[22] ), 
         .C(counter_hi[2]), .Z(n31315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n13_bdd_3_lut_28389.init = 16'hcaca;
    LUT4 pc_3__bdd_3_lut_28703 (.A(\pc[3] ), .B(\pc[11] ), .C(counter_hi[3]), 
         .Z(n30743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_3__bdd_3_lut_28703.init = 16'hcaca;
    LUT4 mux_1532_i8_rep_101_3_lut (.A(\instr_data[3][7] ), .B(n21[7]), 
         .C(n2524), .Z(n29047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i8_rep_101_3_lut.init = 16'hcaca;
    LUT4 mux_2101_i15_3_lut_4_lut (.A(instr[31]), .B(n31838), .C(n31733), 
         .D(n5081[7]), .Z(n3340[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2101_i15_3_lut_4_lut.init = 16'hf808;
    LUT4 n31317_bdd_3_lut (.A(n32282), .B(n29759), .C(counter_hi[3]), 
         .Z(n31318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31317_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_1532_i7_rep_99_3_lut (.A(n6[6]), .B(n21[6]), .C(n2524), .Z(n29045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i7_rep_99_3_lut.init = 16'hcaca;
    LUT4 mux_2101_i14_3_lut_4_lut (.A(instr[31]), .B(n31838), .C(n31733), 
         .D(n5081[6]), .Z(n3340[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2101_i14_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_1528_i7_rep_87_3_lut (.A(n27[6]), .B(n31[6]), .C(n2504), 
         .Z(n29033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i7_rep_87_3_lut.init = 16'hcaca;
    LUT4 mux_1822_i15_3_lut (.A(n21[14]), .B(n27[14]), .C(n2504), .Z(n2505[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1822_i15_3_lut.init = 16'hcaca;
    LUT4 is_store_I_0_469_2_lut_rep_698 (.A(is_store), .B(address_ready), 
         .Z(n31903)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(275[22:47])
    defparam is_store_I_0_469_2_lut_rep_698.init = 16'h8888;
    LUT4 mux_1532_i6_rep_97_3_lut (.A(n6[5]), .B(n21[5]), .C(n2524), .Z(n29043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i6_rep_97_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_510 (.A(is_store), .B(address_ready), 
         .C(mem_op[1]), .D(rst_reg_n), .Z(data_write_n_1__N_369[1])) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(275[22:47])
    defparam i1_2_lut_3_lut_4_lut_adj_510.init = 16'hf7ff;
    LUT4 mux_1528_i6_rep_79_3_lut (.A(n27[5]), .B(n31[5]), .C(n2504), 
         .Z(n29025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i6_rep_79_3_lut.init = 16'hcaca;
    LUT4 mux_1532_i5_rep_95_3_lut (.A(n6[4]), .B(n21[4]), .C(n2524), .Z(n29041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i5_rep_95_3_lut.init = 16'hcaca;
    LUT4 mux_1528_i5_rep_77_3_lut (.A(n27[4]), .B(n31[4]), .C(n2504), 
         .Z(n29023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i5_rep_77_3_lut.init = 16'hcaca;
    LUT4 mux_1826_i15_3_lut (.A(n31[14]), .B(n6[14]), .C(n2524), .Z(n2525[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1826_i15_3_lut.init = 16'hcaca;
    LUT4 n3352_bdd_3_lut_28061_4_lut (.A(instr[31]), .B(n31838), .C(n31733), 
         .D(n30764), .Z(n30765)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3352_bdd_3_lut_28061_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_3_lut_4_lut_adj_511 (.A(is_store), .B(address_ready), 
         .C(mem_op[0]), .D(rst_reg_n), .Z(data_write_n_1__N_369[0])) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(275[22:47])
    defparam i1_2_lut_3_lut_4_lut_adj_511.init = 16'hf7ff;
    LUT4 n3352_bdd_3_lut_28066_4_lut (.A(instr[31]), .B(n31838), .C(n31733), 
         .D(n30772), .Z(n30773)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3352_bdd_3_lut_28066_4_lut.init = 16'hf808;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n31934), .B(n10467), .C(gpio_out_sel[7]), 
         .D(\addr[5] ), .Z(n14)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'hf3f2;
    LUT4 i1_2_lut_4_lut_4_lut_adj_512 (.A(n31934), .B(n10467), .C(gpio_out_sel[6]), 
         .D(\addr[5] ), .Z(n14_adj_12)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_512.init = 16'hf3f2;
    LUT4 i23812_2_lut_4_lut_4_lut (.A(n31934), .B(n10467), .C(\addr[4] ), 
         .D(\addr[5] ), .Z(n26310)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+!(D)))) */ ;
    defparam i23812_2_lut_4_lut_4_lut.init = 16'hfcfd;
    LUT4 i27665_4_lut (.A(debug_instr_valid), .B(is_store), .C(no_write_in_progress), 
         .D(is_load), .Z(stall_core)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(149[50:61])
    defparam i27665_4_lut.init = 16'ha0a2;
    LUT4 i15458_2_lut_4_lut_4_lut (.A(n31934), .B(n10467), .C(n31961), 
         .D(\addr[4] ), .Z(n5171)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C (D))))) */ ;
    defparam i15458_2_lut_4_lut_4_lut.init = 16'h3020;
    LUT4 mux_3131_i21_3_lut_4_lut (.A(instr[31]), .B(n31838), .C(n4285), 
         .D(n3505[17]), .Z(n5121[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3131_i21_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_2119_i1_4_lut (.A(n27694), .B(n27850), .C(n4279), .D(n31755), 
         .Z(n29006)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2119_i1_4_lut.init = 16'hca0a;
    LUT4 i16103_4_lut_4_lut (.A(n31934), .B(n10467), .C(n32027), .D(n28686), 
         .Z(n18680)) /* synthesis lut_function=(!(A (B)+!A (B+!(C (D))))) */ ;
    defparam i16103_4_lut_4_lut.init = 16'h3222;
    LUT4 n3352_bdd_3_lut_28057_4_lut (.A(instr[31]), .B(n31838), .C(n4281), 
         .D(n30760), .Z(n30761)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3352_bdd_3_lut_28057_4_lut.init = 16'hf808;
    LUT4 mux_3126_i5_4_lut_4_lut (.A(instr[31]), .B(n31838), .C(n31764), 
         .D(n4281), .Z(n5081[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3126_i5_4_lut_4_lut.init = 16'ha088;
    LUT4 mux_3126_i10_3_lut_4_lut (.A(instr[31]), .B(n31838), .C(n31733), 
         .D(n29057), .Z(n5081[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3126_i10_3_lut_4_lut.init = 16'hf808;
    LUT4 n3352_bdd_3_lut_28600_4_lut (.A(instr[31]), .B(n31838), .C(n31733), 
         .D(n31684), .Z(n31685)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam n3352_bdd_3_lut_28600_4_lut.init = 16'hf808;
    FD1S3IX counter_hi_3563__i3_rep_860 (.D(n36[1]), .CK(clk_c), .CD(n31980), 
            .Q(n33486));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3563__i3_rep_860.GSR = "DISABLED";
    LUT4 mux_1532_i15_3_lut (.A(n6[14]), .B(n21[14]), .C(n2524), .Z(n2163[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i15_3_lut.init = 16'hcaca;
    LUT4 mux_1528_i15_rep_110_3_lut (.A(n27[14]), .B(n31[14]), .C(n2504), 
         .Z(n29056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i15_rep_110_3_lut.init = 16'hcaca;
    LUT4 n30744_bdd_3_lut (.A(n30744), .B(n30741), .C(n33484), .Z(debug_branch_N_442[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30744_bdd_3_lut.init = 16'hcaca;
    LUT4 pc_2__bdd_3_lut_28050 (.A(\pc[6] ), .B(\pc[14] ), .C(counter_hi[3]), 
         .Z(n30747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_2__bdd_3_lut_28050.init = 16'hcaca;
    LUT4 pc_2__bdd_3_lut_28699 (.A(\pc[2] ), .B(\pc[10] ), .C(counter_hi[3]), 
         .Z(n30748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam pc_2__bdd_3_lut_28699.init = 16'hcaca;
    LUT4 i4820_2_lut_3_lut (.A(n31942), .B(\instr_addr_23__N_318[0] ), .C(instr_addr_23__N_318[1]), 
         .Z(n7103)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam i4820_2_lut_3_lut.init = 16'h8080;
    LUT4 next_instr_write_offset_3__I_0_i2_2_lut_rep_661_3_lut_4_lut (.A(n31942), 
         .B(\instr_addr_23__N_318[0] ), .C(\pc[2] ), .D(instr_addr_23__N_318[1]), 
         .Z(n31866)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam next_instr_write_offset_3__I_0_i2_2_lut_rep_661_3_lut_4_lut.init = 16'h8778;
    LUT4 i1_2_lut_rep_513_3_lut_4_lut (.A(rst_reg_n), .B(clk_c_enable_30), 
         .C(n26), .D(n31838), .Z(n31718)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_513_3_lut_4_lut.init = 16'h0080;
    LUT4 mux_1528_i3_rep_117_3_lut (.A(n27[2]), .B(n31[2]), .C(n2504), 
         .Z(n29063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i3_rep_117_3_lut.init = 16'hcaca;
    LUT4 next_instr_write_offset_3__I_0_i1_2_lut_3_lut (.A(n31942), .B(\instr_addr_23__N_318[0] ), 
         .C(\pc[1] ), .Z(n1)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam next_instr_write_offset_3__I_0_i1_2_lut_3_lut.init = 16'h9696;
    LUT4 mux_346_i1_3_lut_4_lut (.A(n31942), .B(\instr_addr_23__N_318[0] ), 
         .C(debug_ret), .D(return_addr[1]), .Z(n1764_adj_3181[0])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(380[42:147])
    defparam mux_346_i1_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_2119_i16_3_lut_4_lut (.A(n26), .B(n31722), .C(n3381[11]), 
         .D(n5223[14]), .Z(n3422[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (C)) */ ;
    defparam mux_2119_i16_3_lut_4_lut.init = 16'hf870;
    LUT4 mux_1532_i3_3_lut (.A(n6[2]), .B(n21[2]), .C(n2524), .Z(n2163[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i3_3_lut.init = 16'hcaca;
    LUT4 n5587_bdd_3_lut_28435 (.A(counter_hi[2]), .B(instr_data[9]), .C(instr_data[13]), 
         .Z(n31405)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5587_bdd_3_lut_28435.init = 16'he4e4;
    LUT4 n5587_bdd_3_lut_28442 (.A(counter_hi[2]), .B(\qspi_data_buf[9] ), 
         .C(\qspi_data_buf[13] ), .Z(n31406)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5587_bdd_3_lut_28442.init = 16'he4e4;
    LUT4 n26646_bdd_4_lut_28231_4_lut (.A(n31742), .B(n31853), .C(n31784), 
         .D(n27694), .Z(n30947)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam n26646_bdd_4_lut_28231_4_lut.init = 16'hd8cc;
    LUT4 mux_1528_i2_3_lut (.A(n27[1]), .B(n31[1]), .C(n2504), .Z(n2143[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1528_i2_3_lut.init = 16'hcaca;
    LUT4 n30749_bdd_3_lut (.A(n30749), .B(n30746), .C(n33484), .Z(debug_branch_N_442[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30749_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_513 (.A(n33488), .B(clk_c_enable_30), 
         .C(n16_adj_3171), .D(n31838), .Z(n4279)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_513.init = 16'h0080;
    LUT4 mux_2119_i11_3_lut_3_lut_4_lut (.A(n26), .B(n31722), .C(n3271[10]), 
         .D(n3381[11]), .Z(n3422[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_2119_i11_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1532_i2_3_lut (.A(n6[1]), .B(n21[1]), .C(n2524), .Z(n2163[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1532_i2_3_lut.init = 16'hcaca;
    LUT4 i27749_4_lut (.A(n31748), .B(rst_reg_n), .C(debug_ret), .D(n27776), 
         .Z(clk_c_enable_289)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i27749_4_lut.init = 16'h3337;
    LUT4 i1_4_lut_4_lut_adj_514 (.A(n31742), .B(n31791), .C(n22), .D(n9894), 
         .Z(n27576)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i1_4_lut_4_lut_adj_514.init = 16'h0010;
    PFUMX i28099 (.BLUT(n30838), .ALUT(n30837), .C0(n31718), .Z(n30839));
    LUT4 i27877_4_lut (.A(n31748), .B(debug_ret), .C(n31942), .D(n27966), 
         .Z(clk_c_enable_303)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i27877_4_lut.init = 16'h0010;
    LUT4 i27871_4_lut (.A(n31748), .B(rst_reg_n), .C(debug_ret), .D(n27772), 
         .Z(clk_c_enable_305)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i27871_4_lut.init = 16'h3337;
    LUT4 mux_2119_i17_3_lut_3_lut_4_lut (.A(n26), .B(n31722), .C(n5223[15]), 
         .D(n3381[11]), .Z(n3422[16])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_2119_i17_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 i27874_4_lut (.A(n31748), .B(debug_ret), .C(n31942), .D(n27972), 
         .Z(clk_c_enable_319)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i27874_4_lut.init = 16'h0010;
    LUT4 mux_3160_i15_3_lut (.A(n31853), .B(n31851), .C(n31845), .Z(n5223[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3160_i15_3_lut.init = 16'hcaca;
    LUT4 i27868_4_lut (.A(n31748), .B(rst_reg_n), .C(debug_ret), .D(n27780), 
         .Z(clk_c_enable_321)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i27868_4_lut.init = 16'h3337;
    LUT4 n5587_bdd_3_lut_28447 (.A(counter_hi[2]), .B(\qspi_data_buf[11] ), 
         .C(\qspi_data_buf[15] ), .Z(n31416)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5587_bdd_3_lut_28447.init = 16'he4e4;
    LUT4 i1_3_lut_4_lut_adj_515 (.A(n31949), .B(rst_reg_n), .C(data_ready_latch), 
         .D(address_ready), .Z(clk_c_enable_375)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_515.init = 16'hff7f;
    LUT4 i1_3_lut_4_lut_adj_516 (.A(n31949), .B(rst_reg_n), .C(data_ready_latch), 
         .D(data_ready_ext), .Z(n27110)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_516.init = 16'h0800;
    LUT4 n3520_bdd_3_lut_28060 (.A(n3505[17]), .B(n30761), .C(n4285), 
         .Z(n30762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3520_bdd_3_lut_28060.init = 16'hcaca;
    LUT4 i1_3_lut_adj_517 (.A(n35), .B(n26_adj_3172), .C(n27956), .Z(n27960)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_517.init = 16'h8080;
    LUT4 i1_4_lut_adj_518 (.A(n31748), .B(debug_ret), .C(n31942), .D(n27998), 
         .Z(clk_c_enable_342)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(410[18] 430[16])
    defparam i1_4_lut_adj_518.init = 16'h1000;
    LUT4 n5587_bdd_3_lut_28443 (.A(counter_hi[2]), .B(instr_data[11]), .C(instr_data[15]), 
         .Z(n31415)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5587_bdd_3_lut_28443.init = 16'he4e4;
    LUT4 n5587_bdd_3_lut (.A(counter_hi[2]), .B(\qspi_data_buf[10] ), .C(\qspi_data_buf[14] ), 
         .Z(n31424)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5587_bdd_3_lut.init = 16'he4e4;
    LUT4 n5587_bdd_3_lut_28448 (.A(counter_hi[2]), .B(instr_data[10]), .C(instr_data[14]), 
         .Z(n31423)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n5587_bdd_3_lut_28448.init = 16'he4e4;
    LUT4 i1_2_lut_3_lut_4_lut_adj_519 (.A(n32027), .B(n31962), .C(n31899), 
         .D(\addr[4] ), .Z(clk_c_enable_273)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_519.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_520 (.A(rst_reg_n), .B(clk_c_enable_30), 
         .C(n26_adj_3172), .D(n31838), .Z(n4269)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_520.init = 16'h0080;
    LUT4 n31792_bdd_4_lut_28720 (.A(n31792), .B(data_txn_len[0]), .C(instr_data[14]), 
         .D(instr_data[6]), .Z(n32279)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam n31792_bdd_4_lut_28720.init = 16'hfd20;
    LUT4 mux_3160_i14_3_lut (.A(n31853), .B(n31847), .C(n31845), .Z(n5223[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3160_i14_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_521 (.A(n32027), .B(n31962), .C(n31899), 
         .D(\addr[4] ), .Z(clk_c_enable_357)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_521.init = 16'h0020;
    LUT4 mux_3160_i13_3_lut (.A(n31853), .B(n31852), .C(n31845), .Z(n5223[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3160_i13_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_522 (.A(\addr[4] ), .B(n31962), .C(n31899), 
         .D(n26266), .Z(clk_c_enable_349)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_4_lut_adj_522.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_523 (.A(\addr[4] ), .B(n31962), .C(n31899), 
         .D(n32003), .Z(clk_c_enable_259)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(260[12] 268[8])
    defparam i1_2_lut_3_lut_4_lut_adj_523.init = 16'h2000;
    LUT4 mux_3160_i12_3_lut (.A(n31853), .B(n31846), .C(n31845), .Z(n5223[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3160_i12_3_lut.init = 16'hcaca;
    LUT4 mux_2096_i11_4_lut (.A(n31865), .B(n31778), .C(n4279), .D(n31845), 
         .Z(n3271[10])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_2096_i11_4_lut.init = 16'hc0ca;
    LUT4 mux_1538_i15_3_lut (.A(n29056), .B(n2163[14]), .C(n31944), .Z(instr[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[36:78])
    defparam mux_1538_i15_3_lut.init = 16'hcaca;
    LUT4 n17863_bdd_3_lut_28591 (.A(n2163[14]), .B(n29056), .C(n31944), 
         .Z(n30759)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n17863_bdd_3_lut_28591.init = 16'hacac;
    LUT4 i1_2_lut_3_lut_4_lut_adj_524 (.A(n31962), .B(\addr[4] ), .C(n31899), 
         .D(n32003), .Z(clk_c_enable_360)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_524.init = 16'h1000;
    LUT4 n4275_bdd_3_lut_28076 (.A(n4263), .B(instr[31]), .C(instr[19]), 
         .Z(n30764)) /* synthesis lut_function=(A (B)+!A (C)) */ ;
    defparam n4275_bdd_3_lut_28076.init = 16'hd8d8;
    LUT4 i1_2_lut_3_lut_4_lut_adj_525 (.A(rst_reg_n), .B(clk_c_enable_30), 
         .C(n19_c), .D(n31838), .Z(n4271)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_525.init = 16'h0080;
    LUT4 n15_bdd_4_lut (.A(n31845), .B(n31868), .C(n31790), .D(n31869), 
         .Z(n31472)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;
    defparam n15_bdd_4_lut.init = 16'hc800;
    PFUMX mux_1538_i4 (.BLUT(n2143[3]), .ALUT(n2163[3]), .C0(n31944), 
          .Z(instr[19]));
    PFUMX mux_1538_i9 (.BLUT(n2143[8]), .ALUT(n2163[8]), .C0(n31944), 
          .Z(instr[24]));
    PFUMX mux_1538_i10 (.BLUT(n2143[9]), .ALUT(n2163[9]), .C0(n31944), 
          .Z(instr[25]));
    LUT4 i1_2_lut_rep_699_3_lut (.A(n31964), .B(\addr[9] ), .C(n10467), 
         .Z(n31904)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_699_3_lut.init = 16'hfefe;
    PFUMX mux_1538_i12 (.BLUT(n2143[11]), .ALUT(n2163[11]), .C0(n31944), 
          .Z(instr[27]));
    LUT4 i1_4_lut_adj_526 (.A(n31853), .B(n33488), .C(n31849), .D(n31867), 
         .Z(n27892)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_526.init = 16'hc088;
    LUT4 connect_peripheral_3__I_1_i4_3_lut_rep_674_3_lut_4_lut (.A(n31964), 
         .B(\addr[9] ), .C(\addr[5] ), .D(n10467), .Z(n31879)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam connect_peripheral_3__I_1_i4_3_lut_rep_674_3_lut_4_lut.init = 16'h00fe;
    LUT4 i1_4_lut_adj_527 (.A(n31850), .B(n33488), .C(n31848), .D(n31867), 
         .Z(n27868)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_527.init = 16'hc088;
    LUT4 connect_peripheral_3__I_1_i3_3_lut_rep_680_3_lut_4_lut (.A(n31964), 
         .B(\addr[9] ), .C(\addr[4] ), .D(n10467), .Z(n31885)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam connect_peripheral_3__I_1_i3_3_lut_rep_680_3_lut_4_lut.init = 16'h00fe;
    PFUMX mux_1538_i13 (.BLUT(n2143[12]), .ALUT(n2163[12]), .C0(n31944), 
          .Z(instr[28]));
    LUT4 i27929_2_lut_3_lut_4_lut (.A(n31964), .B(\addr[9] ), .C(\addr[4] ), 
         .D(n10467), .Z(n4)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i27929_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i6038_3_lut_3_lut_4_lut (.A(n31964), .B(\addr[9] ), .C(n32027), 
         .D(n10467), .Z(n19)) /* synthesis lut_function=(A (D)+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i6038_3_lut_3_lut_4_lut.init = 16'hff01;
    PFUMX mux_1538_i14 (.BLUT(n2143[13]), .ALUT(n2163[13]), .C0(n31944), 
          .Z(instr[29]));
    LUT4 mux_3160_i16_3_lut (.A(n31853), .B(n31850), .C(n31845), .Z(n5223[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(178[18] 213[12])
    defparam mux_3160_i16_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_528 (.A(n31804), .B(n31830), .C(n31803), .D(n31860), 
         .Z(n4_adj_3136)) /* synthesis lut_function=(!((B (C (D))+!B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_528.init = 16'h0a88;
    PFUMX i28085 (.BLUT(n30804), .ALUT(n30803), .C0(counter_hi[2]), .Z(n30805));
    LUT4 i1_4_lut_adj_529 (.A(clk_c_enable_325), .B(n31838), .C(n31831), 
         .D(n31802), .Z(n2810)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_529.init = 16'ha888;
    LUT4 i1_4_lut_adj_530 (.A(clk_c_enable_325), .B(n31838), .C(n20), 
         .D(n25), .Z(n2812)) /* synthesis lut_function=(A (B+!(C+(D)))) */ ;
    defparam i1_4_lut_adj_530.init = 16'h888a;
    LUT4 i1_4_lut_adj_531 (.A(n31868), .B(n31853), .C(n31763), .D(n31762), 
         .Z(n26119)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_531.init = 16'h22a0;
    LUT4 n3520_bdd_3_lut_28064 (.A(n3505[17]), .B(n30766), .C(n4285), 
         .Z(n30767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3520_bdd_3_lut_28064.init = 16'hcaca;
    LUT4 i1_2_lut_adj_532 (.A(n26_adj_3172), .B(n27956), .Z(n27922)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_532.init = 16'h8888;
    PFUMX i28592 (.BLUT(n31685), .ALUT(n31682), .C0(n4281), .Z(n31686));
    LUT4 i1_4_lut_adj_533 (.A(n31853), .B(n33488), .C(n31863), .D(n31867), 
         .Z(n27880)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_533.init = 16'hc088;
    LUT4 i21205_2_lut (.A(counter_hi[3]), .B(counter_hi[2]), .Z(n36[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam i21205_2_lut.init = 16'h6666;
    LUT4 i21226_4_lut (.A(n31734), .B(n28282), .C(addr_offset[3]), .D(instr_complete_N_1647), 
         .Z(n33[1])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(183[18] 213[12])
    defparam i21226_4_lut.init = 16'h6ca0;
    FD1S3IX counter_hi_3563__i4_rep_858 (.D(n36[2]), .CK(clk_c), .CD(n31980), 
            .Q(n33484));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(241[27:41])
    defparam counter_hi_3563__i4_rep_858.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_534 (.A(n31853), .B(n33488), .C(n31865), .D(n31867), 
         .Z(n27928)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_534.init = 16'hc088;
    LUT4 i1_3_lut_4_lut_adj_535 (.A(n31838), .B(rst_reg_n), .C(n4_adj_3136), 
         .D(n9894), .Z(n27810)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_535.init = 16'h0040;
    LUT4 i1_4_lut_adj_536 (.A(n31853), .B(n33488), .C(n31864), .D(n31867), 
         .Z(n27904)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_536.init = 16'hc088;
    LUT4 n4263_bdd_3_lut_28065 (.A(n2163[2]), .B(n31944), .C(n29063), 
         .Z(n30771)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n4263_bdd_3_lut_28065.init = 16'hb8b8;
    LUT4 i1_3_lut_4_lut_adj_537 (.A(n31838), .B(n33488), .C(n28864), .D(n9894), 
         .Z(n28128)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_537.init = 16'h0004;
    LUT4 n30771_bdd_3_lut (.A(n30771), .B(instr[31]), .C(n4263), .Z(n30772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30771_bdd_3_lut.init = 16'hcaca;
    L6MUX21 i28723 (.D0(n32281), .D1(n32278), .SD(n30170), .Z(n32282));
    PFUMX i28721 (.BLUT(n32280), .ALUT(n32279), .C0(counter_hi[2]), .Z(n32281));
    PFUMX i28622 (.BLUT(n32078), .ALUT(n32079), .C0(n31944), .Z(instr[31]));
    PFUMX i28619 (.BLUT(n32074), .ALUT(n32075), .C0(n31944), .Z(n32076));
    PFUMX i28617 (.BLUT(n32070), .ALUT(n32071), .C0(counter_hi[2]), .Z(n32072));
    LUT4 n3520_bdd_3_lut_28069 (.A(n3505[17]), .B(n30774), .C(n4285), 
         .Z(n30775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3520_bdd_3_lut_28069.init = 16'hcaca;
    tinyQV_time i_timer (.timer_interrupt(timer_interrupt), .clk_c(clk_c), 
            .clk_c_enable_36(clk_c_enable_36), .mtimecmp({Open_73, Open_74, 
            Open_75, Open_76, Open_77, Open_78, Open_79, Open_80, 
            Open_81, Open_82, Open_83, Open_84, Open_85, Open_86, 
            Open_87, Open_88, Open_89, Open_90, Open_91, Open_92, 
            Open_93, Open_94, Open_95, Open_96, mtimecmp[7:6], Open_97, 
            Open_98, Open_99, Open_100, Open_101, Open_102}), .\mtimecmp[5] (mtimecmp[5]), 
            .\mtimecmp[4] (mtimecmp[4]), .n31980(n31980), .mtimecmp_2__N_1939(mtimecmp_2__N_1939), 
            .mtimecmp_3__N_1935(mtimecmp_3__N_1935), .mtimecmp_1__N_1941(mtimecmp_1__N_1941), 
            .mtimecmp_0__N_1943(mtimecmp_0__N_1943), .time_pulse_r(time_pulse_r), 
            .clk_c_enable_249(clk_c_enable_249), .n31913(n31913), .\addr[2] (\addr[2] ), 
            .timer_data({timer_data}), .\mtime_out[0] (mtime_out[0]), .n10573(n10573), 
            .cy(cy), .rst_reg_n(rst_reg_n), .instr_fetch_stopped(instr_fetch_stopped), 
            .instr_fetch_running_N_945(instr_fetch_running_N_945), .n28156(n28156), 
            .address_ready(address_ready), .is_store(is_store), .clk_c_enable_109(clk_c_enable_109), 
            .\instr_data[1] (instr_data[1]), .\instr_data_0__15__N_638[49] (instr_data_0__15__N_638[49]), 
            .n31876(n31876), .n31957(n31957), .n31946(n31946), .clk_c_enable_449(clk_c_enable_449), 
            .no_write_in_progress(no_write_in_progress), .clk_c_enable_157(clk_c_enable_157), 
            .n33488(n33488), .n31966(n31966), .\cycle_count_wide[3] (cycle_count_wide[3]), 
            .n31870(n31870), .clk_c_enable_233(clk_c_enable_233), .n31893(n31893), 
            .is_double_fault_r(is_double_fault_r), .mstatus_mte(mstatus_mte), 
            .n31841(n31841), .clk_c_enable_107(clk_c_enable_107), .\reg_access[3][2] (\reg_access[3] [2]), 
            .clk_c_enable_177(clk_c_enable_177), .n32033(n32033), .is_timer_addr(is_timer_addr), 
            .n8(n8), .n28028(n28028), .n31748(n31748), .n26290(n26290), 
            .mstatus_mie_N_1709(mstatus_mie_N_1709), .n31878(n31878), .mstatus_mie_N_1707(mstatus_mie_N_1707), 
            .n15604(n15604), .clk_c_enable_161(clk_c_enable_161), .n31742(n31742), 
            .n31737(n31737), .clk_c_enable_347(clk_c_enable_347), .\instr_data[0] (instr_data[0]), 
            .\instr_data_0__15__N_638[0] (instr_data_0__15__N_638[0]), .n31884(n31884), 
            .n31872(n31872), .n31889(n31889), .data_out_slice({\data_out_slice[3] , 
            data_out_slice[2:0]}), .n31840(n31840)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(450[17] 461[6])
    tinyqv_decoder i_decoder (.n31850(n31850), .n31441(n31441), .n31860(n31860), 
            .n31402(n31402), .n31774(n31774), .n31869(n31869), .n31814(n31814), 
            .n31847(n31847), .n31821(n31821), .n31820(n31820), .\instr[26] (instr[26]), 
            .n31837(n31837), .n31849(n31849), .n31865(n31865), .n31845(n31845), 
            .n10904(n10904), .n31848(n31848), .n31763(n31763), .n31867(n31867), 
            .n32(n32_adj_3168), .\mem_op_2__N_1114[1] (mem_op_2__N_1114[1]), 
            .n31772(n31772), .n31773(n31773), .n31833(n31833), .n31868(n31868), 
            .n31823(n31823), .n31853(n31853), .n31194(n31194), .n4269(n4269), 
            .n31852(n31852), .n31851(n31851), .n3265(n3234[1]), .n31846(n31846), 
            .n31813(n31813), .n31799(n31799), .n31817(n31817), .n3006(n2982[8]), 
            .n31784(n31784), .n31764(n31764), .n31838(n31838), .\mem_op_de[1] (mem_op_de[1]), 
            .n31786(n31786), .n31766(n31766), .n31758(n31758), .n31796(n31796), 
            .n17976(n17976), .n31790(n31790), .n7(n7), .n10(n10), .n24(n24_adj_3160), 
            .\alu_op_3__N_1170[2] (alu_op_3__N_1170[2]), .n28366(n28366), 
            .\additional_mem_ops_2__N_1132[0] (additional_mem_ops_2__N_1132[0]), 
            .n31795(n31795), .n31864(n31864), .n8302(n8302), .n31471(n31471), 
            .n41(n41), .n32_adj_3(n32), .n30(n30_adj_3165), .n4(n4_adj_3163), 
            .n31762(n31762), .n31816(n31816), .is_auipc_de(is_auipc_de), 
            .n29004(n29004), .n31863(n31863), .n31769(n31769), .n31798(n31798), 
            .n22(n22_adj_3167), .\instr[27] (instr[27]), .n3365(n3340[7]), 
            .n33488(n33488), .n27746(n27746), .n28332(n28332), .n31791(n31791), 
            .n9894(n9894), .n28006(n28006), .n17998(n17998), .n31861(n31861), 
            .n31733(n31733), .n27246(n27246), .n31944(n31944), .n4281(n4281), 
            .n29375(n29375), .\instr[16] (instr[16]), .n2610(n2607[1]), 
            .\instr[25] (instr[25]), .n3367(n3340[5]), .n2169(n2163[10]), 
            .n29048(n29048), .mem_op_increment_reg_de(mem_op_increment_reg_de), 
            .n4263(n4263), .n31732(n31732), .n28898(n28898), .n10068(n10068), 
            .n4_adj_4(n4_adj_3169), .n13248(n13248), .\instr[30] (instr[30]), 
            .n3(n3), .n28871(n28871), .n26113(n26113), .rst_reg_n(rst_reg_n), 
            .n27850(n27850), .is_alu_imm_de(is_alu_imm_de), .n31831(n31831), 
            .is_jalr_N_1370(is_jalr_N_1370), .\instr[31] (instr[31]), .n5137(n5121[15]), 
            .n5140(n5121[12]), .\instr[29] (instr[29]), .n5123(n5121[29]), 
            .\instr[24] (instr[24]), .n5128(n5121[24]), .n5127(n5121[25]), 
            .n30771(n30771), .n30770(n30770), .n31728(n31728), .\instr[28] (instr[28]), 
            .n5124(n5121[28]), .n30759(n30759), .n30760(n30760), .\instr[19] (instr[19]), 
            .n30763(n30763), .n29041(n29041), .n29018(n29018), .n29049(n29049), 
            .n5125(n5121[27]), .n5136(n5121[16]), .n29043(n29043), .n29020(n29020), 
            .n29045(n29045), .n29026(n29026), .n29047(n29047), .n29028(n29028), 
            .\instr[17] (instr[17]), .n31682(n31682), .n5139(n5121[13]), 
            .n5138(n5121[14]), .n31818(n31818), .n15(n15_adj_3143), .alu_op_de({alu_op_de}), 
            .n30_adj_5(n30), .n31835(n31835), .n31436(n31436), .is_alu_reg_de(is_alu_reg_de), 
            .n31824(n31824), .n31822(n31822), .is_store_de(is_store_de), 
            .is_lui_N_1365(is_lui_N_1365), .is_lui_de(is_lui_de), .n157(n155[2]), 
            .n31815(n31815), .n3001(n2982[13]), .n8(n8_adj_3147), .n29215(n29215), 
            .is_load_de(is_load_de), .n15_adj_6(n15_adj_3139), .n30_adj_7(n30_adj_3145), 
            .is_jal_de(is_jal_de), .is_jalr_de(is_jalr_de), .clk_c_enable_325(clk_c_enable_325), 
            .n4285(n4285), .n26(n26), .n29385(n29385), .n22_adj_8(n22), 
            .n31760(n31760), .n31714(n31714), .n5147(n5121[5]), .n5152(n5121[0]), 
            .n5148(n5121[4]), .n5145(n5121[7]), .n31830(n31830), .n31809(n31809), 
            .is_branch_de(is_branch_de), .n2998(n2982[16]), .n26202(n26202), 
            .n27956(n27956), .n28032(n28032), .n28864(n28864), .n28040(n28040), 
            .n27790(n27790), .n27928(n27928), .n26_adj_9(n26_adj_3172), 
            .n27934(n27934), .n27688(n27688), .n19(n19_c), .n27694(n27694), 
            .n28060(n28060), .n28068(n28068), .n31805(n31805), .n28054(n28054), 
            .n12(n12_adj_3176), .n2810(n2810), .n2604(n2602[2]), .n2632(n2630[2]), 
            .n27892(n27892), .n27898(n27898), .n27880(n27880), .n27886(n27886), 
            .n27904(n27904), .n27910(n27910), .n31785(n31785), .\mem_op_de[2] (mem_op_de[2]), 
            .n27832(n27832), .n27838(n27838), .n19_adj_10(n19_adj_3141), 
            .n26478(n26478), .n27868(n27868), .n27874(n27874), .n27818(n27818), 
            .n27824(n27824), .is_system_de(is_system_de)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    tinyqv_core i_core (.clk_c(clk_c), .n31841(n31841), .n31980(n31980), 
            .clk_c_enable_234(clk_c_enable_234), .counter_hi({counter_hi}), 
            .n92({n92}), .n18324(n18324), .instr_complete_N_1647(instr_complete_N_1647), 
            .clk_c_enable_449(clk_c_enable_449), .\ui_in_sync[0] (\ui_in_sync[0] ), 
            .mstatus_mte(mstatus_mte), .\imm[10] (\imm[10] ), .n31744(n31744), 
            .n31738(n31738), .n27838(n27838), .n31742(n31742), .n26648(n26648), 
            .\imm[1] (\imm[1] ), .n27934(n27934), .n26764(n26764), .n27874(n27874), 
            .n26794(n26794), .data_rs1({Open_103, Open_104, Open_105, 
            data_rs1[0]}), .n27810(n27810), .n2804(n2804), .n27886(n27886), 
            .n26788(n26788), .n28020(n28020), .n2498(n2498), .n27960(n27960), 
            .n3402(n3381[11]), .n28068(n28068), .n26807(n26807), .n28080(n28080), 
            .n26889(n26889), .n27672(n27672), .n31758(n31758), .n31733(n31733), 
            .n27862(n27862), .n2592(n2589[1]), .n9894(n9894), .n27728(n27728), 
            .n27734(n27734), .\next_pc_for_core[7] (\next_pc_for_core[7] ), 
            .\next_pc_for_core[3] (\next_pc_for_core[3] ), .n27910(n27910), 
            .n26776(n26776), .\next_pc_for_core[23] (\next_pc_for_core[23] ), 
            .\next_pc_for_core[19] (\next_pc_for_core[19] ), .n28116(n28116), 
            .n26871(n26871), .n27946(n27946), .n31735(n31735), .\next_pc_for_core[15] (\next_pc_for_core[15] ), 
            .\next_pc_for_core[11] (\next_pc_for_core[11] ), .n27922(n27922), 
            .n26770(n26770), .\alu_op[0] (alu_op[0]), .\alu_op[3] (alu_op[3]), 
            .\alu_op[1] (alu_op[1]), .\alu_op_in[2] (alu_op_in[2]), .n29006(n29006), 
            .n28881(n28881), .n27738(n27738), .n27744(n27744), .n27898(n27898), 
            .n26782(n26782), .n30947(n30947), .n31853(n31853), .n30949(n30949), 
            .n27790(n27790), .n12(n12_adj_3176), .n27796(n27796), .n28128(n28128), 
            .n26827(n26827), .n28140(n28140), .n26905(n26905), .n28054(n28054), 
            .n26814(n26814), .n31894(n31894), .n31875(n31875), .n1160(n1160), 
            .load_done(load_done), .clk_c_enable_249(clk_c_enable_249), 
            .n8289(n8289), .\imm[2] (\imm[2] ), .\imm[6] (\imm[6] ), .clk_c_enable_233(clk_c_enable_233), 
            .n27576(n27576), .n31720(n31720), .n26800(n26800), .n31838(n31838), 
            .is_jalr_N_1370(is_jalr_N_1370), .n27724(n27724), .n28040(n28040), 
            .n26821(n26821), .stall_core(stall_core), .clk_c_enable_36(clk_c_enable_36), 
            .n28204(n28204), .n26993(n26993), .is_double_fault_r(is_double_fault_r), 
            .n31893(n31893), .n31878(n31878), .n28092(n28092), .n26883(n26883), 
            .n28104(n28104), .n26877(n26877), .n27824(n27824), .n26656(n26656), 
            .\imm[0] (imm[0]), .cycle({cycle_c[1], cycle[0]}), .n10486(n10486), 
            .\alu_b_in[3] (\alu_b_in[3] ), .n31949(n31949), .n31946(n31946), 
            .n4325(n4322[0]), .\additional_mem_ops_2__N_749[0] (additional_mem_ops_2__N_749[0]), 
            .n27018(n27018), .n31741(n31741), .n32040(n32040), .is_load(is_load), 
            .n844(n844), .n26290(n26290), .clk_c_enable_527(clk_c_enable_527), 
            .n32046(n32046), .interrupt_core(interrupt_core), .n31876(n31876), 
            .n5014({n5014}), .n1766(n1764_adj_3181[1]), .\instr_write_offset_3__N_934[1] (instr_write_offset_3__N_934[1]), 
            .\debug_branch_N_450[1] (debug_branch_N_450[1]), .n1767(n1764_adj_3181[0]), 
            .\instr_write_offset_3__N_934[0] (instr_write_offset_3__N_934[0]), 
            .n15(n15_adj_3148), .n31743(n31743), .n1768({n34}), .pc_2__N_932({pc_2__N_932}), 
            .n29665(n29665), .n31311(n31311), .debug_rd({debug_rd}), .instr_fetch_running(instr_fetch_running), 
            .was_early_branch(was_early_branch), .n31745(n31745), .n31957(n31957), 
            .\ui_in_sync[1] (\ui_in_sync[1] ), .debug_rd_3__N_1575(debug_rd_3__N_1575), 
            .n31915(n31915), .n31892(n31892), .load_done_N_1741(load_done_N_1741), 
            .\data_rs2[0] (data_rs2[0]), .\data_rs2[2] (data_rs2[2]), .n84(n84), 
            .\data_rs2[1] (data_rs2[1]), .\next_fsm_state_3__N_3015[3] (\next_fsm_state_3__N_3015[3] ), 
            .rd({rd_c[3:1], rd[0]}), .fsm_state({fsm_state}), .debug_instr_valid(debug_instr_valid), 
            .is_lui(is_lui), .is_jal(is_jal), .n31948(n31948), .n31966(n31966), 
            .clk_c_enable_169(clk_c_enable_169), .is_branch(is_branch), 
            .is_jalr(is_jalr), .is_auipc(is_auipc), .is_system(is_system), 
            .n33486(n33486), .n33484(n33484), .clk_c_enable_165(clk_c_enable_165), 
            .\imm[5] (\imm[5] ), .\imm[3] (\imm[3] ), .n32015(n32015), 
            .mem_op({mem_op}), .n31987(n31987), .n26175(n26175), .n31955(n31955), 
            .accum({accum}), .d_3__N_1868({d_3__N_1868}), .n31929(n31929), 
            .timer_interrupt(timer_interrupt), .clk_c_enable_181(clk_c_enable_181), 
            .\mul_out[1] (\mul_out[1] ), .clk_c_enable_184(clk_c_enable_184), 
            .n32185(n32185), .\timer_data[0] (timer_data[0]), .is_timer_addr(is_timer_addr), 
            .\mul_out[2] (\mul_out[2] ), .data_out_3__N_1385(data_out_3__N_1385), 
            .n29318(n29318), .n31319(n31319), .\timer_data[2] (timer_data[2]), 
            .\mul_out[3] (\mul_out[3] ), .n31999(n31999), .\debug_branch_N_450[3] (debug_branch_N_450[3]), 
            .load_top_bit(load_top_bit), .n5677({n5677}), .\imm[7] (\imm[7] ), 
            .n9033(n9033), .\imm[11] (\imm[11] ), .is_alu_imm(is_alu_imm), 
            .is_alu_reg(is_alu_reg), .debug_rd_3__N_413(debug_rd_3__N_413), 
            .\cycle_count_wide[3] (cycle_count_wide[3]), .n5626(n5624[2]), 
            .n32049(n32049), .\imm[9] (\imm[9] ), .\imm[8] (\imm[8] ), 
            .\addr_out[26] (addr_out[26]), .\imm[4] (\imm[4] ), .\addr_out[25] (addr_out[25]), 
            .\addr_out[24] (addr_out[24]), .\addr_out[27] (addr_out[27]), 
            .mstatus_mie_N_1709(mstatus_mie_N_1709), .mstatus_mie_N_1707(mstatus_mie_N_1707), 
            .n26997(n26997), .n28222(n28222), .n26995(n26995), .n109(n108[3]), 
            .n26996(n26996), .n31963(n31963), .n31932(n31932), .next_bit(next_bit), 
            .n28800(n28800), .n31389(n31389), .\data_out_slice[0] (data_out_slice[0]), 
            .is_store(is_store), .n9710(n9710), .n29739(n29739), .n13(n13), 
            .n29194(n29194), .n29137(n29137), .n29330(n29330), .\debug_branch_N_450[0] (debug_branch_N_450[0]), 
            .n32044(n32044), .n32039(n32039), .n29190(n29190), .n29149(n29149), 
            .\debug_branch_N_446[28] (debug_branch_N_446[28]), .n238(n234[0]), 
            .n29240(n29240), .n31768(n31768), .data_ready_sync(data_ready_sync), 
            .data_ready_core(data_ready_core), .\next_pc_for_core[20] (\next_pc_for_core[20] ), 
            .\next_pc_for_core[16] (\next_pc_for_core[16] ), .n225(n225_adj_3166), 
            .\pc[23] (\pc[23] ), .\pc[19] (\pc[19] ), .n30741(n30741), 
            .\pc[21] (\pc[21] ), .\pc[17] (\pc[17] ), .n30802(n30802), 
            .\next_pc_for_core[22] (\next_pc_for_core[22] ), .\next_pc_for_core[18] (\next_pc_for_core[18] ), 
            .n227(n227), .\pc[20] (\pc[20] ), .\pc[16] (\pc[16] ), .n225_adj_1(n225), 
            .\pc[22] (\pc[22] ), .\pc[18] (\pc[18] ), .n30746(n30746), 
            .\next_pc_for_core[21] (\next_pc_for_core[21] ), .\next_pc_for_core[17] (\next_pc_for_core[17] ), 
            .n226(n226), .\debug_branch_N_442[31] (debug_branch_N_442[31]), 
            .alu_a_in_3__N_1552(alu_a_in_3__N_1552), .\debug_branch_N_442[30] (debug_branch_N_442[30]), 
            .\debug_rd_3__N_405[30] (debug_rd_3__N_405[30]), .alu_b_in_3__N_1504(alu_b_in_3__N_1504), 
            .\debug_rd_3__N_405[29] (debug_rd_3__N_405[29]), .n157(n157_adj_3152), 
            .\debug_branch_N_442[28] (debug_branch_N_442[28]), .n29220(n29220), 
            .\debug_rd_3__N_405[28] (debug_rd_3__N_405[28]), .\debug_branch_N_442[29] (debug_branch_N_442[29]), 
            .n29147(n29147), .\debug_branch_N_446[30] (debug_branch_N_446[30]), 
            .n29333(n29333), .n29135(n29135), .\debug_branch_N_446[29] (debug_branch_N_446[29]), 
            .n15604(n15604), .\data_out_slice[2] (data_out_slice[2]), .\data_out_slice[1] (data_out_slice[1]), 
            .n31972(n31972), .n31914(n31914), .\timer_data[1] (timer_data[1]), 
            .\mem_data_from_read[17] (\mem_data_from_read[17] ), .\mem_data_from_read[21] (\mem_data_from_read[21] ), 
            .n31310(n31310), .\addr_offset[2] (addr_offset[2]), .n701(n699[0]), 
            .n29012(n29012), .n29162(n29162), .\debug_rd_3__N_405[31] (\debug_rd_3__N_405[31] ), 
            .rst_reg_n(rst_reg_n), .cy(cy), .time_pulse_r(time_pulse_r), 
            .n10573(n10573), .n31889(n31889), .n9538(n9538), .\mtime_out[0] (mtime_out[0]), 
            .n31913(n31913), .n31872(n31872), .\addr_out[23] (addr_out[23]), 
            .\addr_out[0] (addr_out[0]), .\addr_out[1] (addr_out[1]), .n31898(n31898), 
            .\addr_out[22] (addr_out[22]), .\addr_out[21] (addr_out[21]), 
            .\addr_out[20] (addr_out[20]), .\addr_out[19] (addr_out[19]), 
            .\addr_out[18] (addr_out[18]), .\addr_out[17] (addr_out[17]), 
            .\addr_out[16] (addr_out[16]), .\addr_out[15] (addr_out[15]), 
            .\addr_out[14] (addr_out[14]), .\addr_out[13] (addr_out[13]), 
            .\addr_out[12] (addr_out[12]), .\addr_out[11] (addr_out[11]), 
            .\addr_out[10] (addr_out[10]), .\addr_out[9] (addr_out[9]), 
            .\addr_out[8] (addr_out[8]), .\addr_out[7] (addr_out[7]), .\addr_out[6] (addr_out[6]), 
            .\addr_out[5] (addr_out[5]), .\addr_out[4] (addr_out[4]), .\addr_out[3] (addr_out[3]), 
            .n33493(n33493), .instr_complete_N_1651(instr_complete_N_1651), 
            .n5661(n5659[2]), .n28282(n28282), .\next_pc_offset[3] (next_pc_offset[3]), 
            .n27604(n27604), .n31888(n31888), .n18086(n18086), .\debug_branch_N_446[31] (debug_branch_N_446[31]), 
            .\csr_read_3__N_1443[0] (csr_read_3__N_1443[0]), .\csr_read_3__N_1447[2] (\csr_read_3__N_1447[2] ), 
            .GND_net(GND_net), .VCC_net(VCC_net), .\next_accum[5] (\next_accum[5] ), 
            .\next_accum[6] (\next_accum[6] ), .\next_accum[7] (\next_accum[7] ), 
            .\next_accum[8] (\next_accum[8] ), .\next_accum[9] (\next_accum[9] ), 
            .\next_accum[10] (\next_accum[10] ), .\next_accum[11] (\next_accum[11] ), 
            .\next_accum[12] (\next_accum[12] ), .\next_accum[13] (\next_accum[13] ), 
            .\next_accum[14] (\next_accum[14] ), .\next_accum[15] (\next_accum[15] ), 
            .\next_accum[16] (\next_accum[16] ), .\next_accum[17] (\next_accum[17] ), 
            .\next_accum[18] (\next_accum[18] ), .\next_accum[19] (\next_accum[19] ), 
            .\next_accum[4] (\next_accum[4] ), .rs2({rs2}), .n12_adj_2(n12), 
            .n11(n11), .n9(n9), .n8(n8_adj_13), .rs1({rs1_c[3:1], rs1[0]}), 
            .return_addr({return_addr}), .\registers[5][7] (\registers[5][7] ), 
            .\registers[6][7] (\registers[6][7] ), .\registers[7][7] (\registers[7][7] ), 
            .n27480(n27480), .n31747(n31747), .no_write_in_progress(no_write_in_progress), 
            .n28150(n28150), .n27762(n27762), .n28182(n28182), .n29747(n29747), 
            .n4(n4_adj_14), .\reg_access[3][2] (\reg_access[3] [2]), .n30165(n30165), 
            .n30166(n30166), .n30169(n30169), .n31748(n31748), .n30167(n30167), 
            .n30168(n30168), .n31870(n31870)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(322[72] 368[6])
    
endmodule
//
// Verilog Description of module tinyQV_time
//

module tinyQV_time (timer_interrupt, clk_c, clk_c_enable_36, mtimecmp, 
            \mtimecmp[5] , \mtimecmp[4] , n31980, mtimecmp_2__N_1939, 
            mtimecmp_3__N_1935, mtimecmp_1__N_1941, mtimecmp_0__N_1943, 
            time_pulse_r, clk_c_enable_249, n31913, \addr[2] , timer_data, 
            \mtime_out[0] , n10573, cy, rst_reg_n, instr_fetch_stopped, 
            instr_fetch_running_N_945, n28156, address_ready, is_store, 
            clk_c_enable_109, \instr_data[1] , \instr_data_0__15__N_638[49] , 
            n31876, n31957, n31946, clk_c_enable_449, no_write_in_progress, 
            clk_c_enable_157, n33488, n31966, \cycle_count_wide[3] , 
            n31870, clk_c_enable_233, n31893, is_double_fault_r, mstatus_mte, 
            n31841, clk_c_enable_107, \reg_access[3][2] , clk_c_enable_177, 
            n32033, is_timer_addr, n8, n28028, n31748, n26290, mstatus_mie_N_1709, 
            n31878, mstatus_mie_N_1707, n15604, clk_c_enable_161, n31742, 
            n31737, clk_c_enable_347, \instr_data[0] , \instr_data_0__15__N_638[0] , 
            n31884, n31872, n31889, data_out_slice, n31840) /* synthesis syn_module_defined=1 */ ;
    output timer_interrupt;
    input clk_c;
    input clk_c_enable_36;
    output [31:0]mtimecmp;
    output \mtimecmp[5] ;
    output \mtimecmp[4] ;
    output n31980;
    input mtimecmp_2__N_1939;
    input mtimecmp_3__N_1935;
    input mtimecmp_1__N_1941;
    input mtimecmp_0__N_1943;
    output time_pulse_r;
    input clk_c_enable_249;
    output n31913;
    input \addr[2] ;
    output [3:0]timer_data;
    output \mtime_out[0] ;
    input n10573;
    output cy;
    input rst_reg_n;
    input instr_fetch_stopped;
    input instr_fetch_running_N_945;
    output n28156;
    input address_ready;
    input is_store;
    output clk_c_enable_109;
    input \instr_data[1] ;
    output \instr_data_0__15__N_638[49] ;
    input n31876;
    input n31957;
    input n31946;
    output clk_c_enable_449;
    input no_write_in_progress;
    output clk_c_enable_157;
    input n33488;
    output n31966;
    input \cycle_count_wide[3] ;
    input n31870;
    output clk_c_enable_233;
    input n31893;
    input is_double_fault_r;
    input mstatus_mte;
    output n31841;
    output clk_c_enable_107;
    input \reg_access[3][2] ;
    output clk_c_enable_177;
    input n32033;
    input is_timer_addr;
    input n8;
    input n28028;
    input n31748;
    output n26290;
    input mstatus_mie_N_1709;
    input n31878;
    output mstatus_mie_N_1707;
    input n15604;
    output clk_c_enable_161;
    input n31742;
    input n31737;
    output clk_c_enable_347;
    input \instr_data[0] ;
    output \instr_data_0__15__N_638[0] ;
    output n31884;
    input n31872;
    input n31889;
    input [3:0]data_out_slice;
    input n31840;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire timer_interrupt_N_1954;
    wire [3:0]mtime_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(29[16:25])
    
    wire n4, n32085, n32084;
    wire [31:0]mtimecmp_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(30[16:24])
    
    wire cy_c;
    wire [4:0]comparison;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[16:26])
    
    wire n6, n2;
    
    FD1P3AX timer_interrupt_94 (.D(timer_interrupt_N_1954), .SP(clk_c_enable_36), 
            .CK(clk_c), .Q(timer_interrupt)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(78[12] 80[8])
    defparam timer_interrupt_94.GSR = "DISABLED";
    LUT4 i15451_4_lut_then_4_lut (.A(mtime_out[3]), .B(n4), .C(mtimecmp[6]), 
         .D(mtimecmp[7]), .Z(n32085)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (C+(D)))) */ ;
    defparam i15451_4_lut_then_4_lut.init = 16'h8241;
    LUT4 i15451_4_lut_else_4_lut (.A(mtime_out[3]), .B(n4), .C(mtimecmp[6]), 
         .D(mtimecmp[7]), .Z(n32084)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A (B (C+(D))+!B !(C (D))))) */ ;
    defparam i15451_4_lut_else_4_lut.init = 16'h1824;
    FD1S3AX mtimecmp_30__62 (.D(mtimecmp_c[2]), .CK(clk_c), .Q(mtimecmp_c[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_30__62.GSR = "DISABLED";
    FD1S3AX mtimecmp_29__63 (.D(mtimecmp_c[1]), .CK(clk_c), .Q(mtimecmp_c[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_29__63.GSR = "DISABLED";
    FD1S3AX mtimecmp_28__64 (.D(mtimecmp_c[0]), .CK(clk_c), .Q(mtimecmp_c[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_28__64.GSR = "DISABLED";
    FD1S3AX mtimecmp_27__65 (.D(mtimecmp_c[31]), .CK(clk_c), .Q(mtimecmp_c[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_27__65.GSR = "DISABLED";
    FD1S3AX mtimecmp_26__66 (.D(mtimecmp_c[30]), .CK(clk_c), .Q(mtimecmp_c[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_26__66.GSR = "DISABLED";
    FD1S3AX mtimecmp_25__67 (.D(mtimecmp_c[29]), .CK(clk_c), .Q(mtimecmp_c[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_25__67.GSR = "DISABLED";
    FD1S3AX mtimecmp_24__68 (.D(mtimecmp_c[28]), .CK(clk_c), .Q(mtimecmp_c[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_24__68.GSR = "DISABLED";
    FD1S3AX mtimecmp_23__69 (.D(mtimecmp_c[27]), .CK(clk_c), .Q(mtimecmp_c[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_23__69.GSR = "DISABLED";
    FD1S3AX mtimecmp_22__70 (.D(mtimecmp_c[26]), .CK(clk_c), .Q(mtimecmp_c[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_22__70.GSR = "DISABLED";
    FD1S3AX mtimecmp_21__71 (.D(mtimecmp_c[25]), .CK(clk_c), .Q(mtimecmp_c[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_21__71.GSR = "DISABLED";
    FD1S3AX mtimecmp_20__72 (.D(mtimecmp_c[24]), .CK(clk_c), .Q(mtimecmp_c[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_20__72.GSR = "DISABLED";
    FD1S3AX mtimecmp_19__73 (.D(mtimecmp_c[23]), .CK(clk_c), .Q(mtimecmp_c[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_19__73.GSR = "DISABLED";
    FD1S3AX mtimecmp_18__74 (.D(mtimecmp_c[22]), .CK(clk_c), .Q(mtimecmp_c[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_18__74.GSR = "DISABLED";
    FD1S3AX mtimecmp_17__75 (.D(mtimecmp_c[21]), .CK(clk_c), .Q(mtimecmp_c[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_17__75.GSR = "DISABLED";
    FD1S3AX mtimecmp_16__76 (.D(mtimecmp_c[20]), .CK(clk_c), .Q(mtimecmp_c[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_16__76.GSR = "DISABLED";
    FD1S3AX mtimecmp_15__77 (.D(mtimecmp_c[19]), .CK(clk_c), .Q(mtimecmp_c[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_15__77.GSR = "DISABLED";
    FD1S3AX mtimecmp_14__78 (.D(mtimecmp_c[18]), .CK(clk_c), .Q(mtimecmp_c[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_14__78.GSR = "DISABLED";
    FD1S3AX mtimecmp_13__79 (.D(mtimecmp_c[17]), .CK(clk_c), .Q(mtimecmp_c[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_13__79.GSR = "DISABLED";
    FD1S3AX mtimecmp_12__80 (.D(mtimecmp_c[16]), .CK(clk_c), .Q(mtimecmp_c[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_12__80.GSR = "DISABLED";
    FD1S3AX mtimecmp_11__81 (.D(mtimecmp_c[15]), .CK(clk_c), .Q(mtimecmp_c[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_11__81.GSR = "DISABLED";
    FD1S3AX mtimecmp_10__82 (.D(mtimecmp_c[14]), .CK(clk_c), .Q(mtimecmp_c[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_10__82.GSR = "DISABLED";
    FD1S3AX mtimecmp_9__83 (.D(mtimecmp_c[13]), .CK(clk_c), .Q(mtimecmp_c[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_9__83.GSR = "DISABLED";
    FD1S3AX mtimecmp_8__84 (.D(mtimecmp_c[12]), .CK(clk_c), .Q(mtimecmp_c[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_8__84.GSR = "DISABLED";
    FD1S3AX mtimecmp_7__85 (.D(mtimecmp_c[11]), .CK(clk_c), .Q(mtimecmp[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_7__85.GSR = "DISABLED";
    FD1S3AX mtimecmp_6__86 (.D(mtimecmp_c[10]), .CK(clk_c), .Q(mtimecmp[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_6__86.GSR = "DISABLED";
    FD1S3AX mtimecmp_5__87 (.D(mtimecmp_c[9]), .CK(clk_c), .Q(\mtimecmp[5] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_5__87.GSR = "DISABLED";
    FD1S3AX mtimecmp_4__88 (.D(mtimecmp_c[8]), .CK(clk_c), .Q(\mtimecmp[4] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_4__88.GSR = "DISABLED";
    FD1S3JX cy_93 (.D(comparison[4]), .CK(clk_c), .PD(clk_c_enable_36), 
            .Q(cy_c)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(74[12] 76[8])
    defparam cy_93.GSR = "DISABLED";
    FD1S3AX mtimecmp_31__61 (.D(mtimecmp_c[3]), .CK(clk_c), .Q(mtimecmp_c[31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(60[12:53])
    defparam mtimecmp_31__61.GSR = "DISABLED";
    FD1S3IX mtimecmp_2__90 (.D(mtimecmp_2__N_1939), .CK(clk_c), .CD(n31980), 
            .Q(mtimecmp_c[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_2__90.GSR = "DISABLED";
    FD1S3IX mtimecmp_3__89 (.D(mtimecmp_3__N_1935), .CK(clk_c), .CD(n31980), 
            .Q(mtimecmp_c[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_3__89.GSR = "DISABLED";
    FD1S3IX mtimecmp_1__91 (.D(mtimecmp_1__N_1941), .CK(clk_c), .CD(n31980), 
            .Q(mtimecmp_c[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_1__91.GSR = "DISABLED";
    FD1S3IX mtimecmp_0__92 (.D(mtimecmp_0__N_1943), .CK(clk_c), .CD(n31980), 
            .Q(mtimecmp_c[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(62[12] 69[8])
    defparam mtimecmp_0__92.GSR = "DISABLED";
    FD1S3IX time_pulse_r_95 (.D(n31913), .CK(clk_c), .CD(clk_c_enable_249), 
            .Q(time_pulse_r)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=450, LSE_RLINE=461 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(82[12] 85[8])
    defparam time_pulse_r_95.GSR = "DISABLED";
    LUT4 mtime_out_3__I_0_96_i4_3_lut (.A(mtime_out[3]), .B(mtimecmp[7]), 
         .C(\addr[2] ), .Z(timer_data[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i4_3_lut.init = 16'hcaca;
    LUT4 mtime_out_3__I_0_96_i1_3_lut (.A(\mtime_out[0] ), .B(\mtimecmp[4] ), 
         .C(\addr[2] ), .Z(timer_data[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i1_3_lut.init = 16'hcaca;
    LUT4 mtime_out_3__I_0_96_i2_3_lut (.A(mtime_out[1]), .B(\mtimecmp[5] ), 
         .C(\addr[2] ), .Z(timer_data[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i2_3_lut.init = 16'hcaca;
    LUT4 mtime_out_3__I_0_96_i3_3_lut (.A(mtime_out[2]), .B(mtimecmp[6]), 
         .C(\addr[2] ), .Z(timer_data[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(87[23:64])
    defparam mtime_out_3__I_0_96_i3_3_lut.init = 16'hcaca;
    LUT4 i4617_3_lut (.A(mtime_out[2]), .B(mtimecmp[6]), .C(n4), .Z(n6)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i4617_3_lut.init = 16'hb2b2;
    LUT4 i4610_3_lut (.A(mtime_out[1]), .B(\mtimecmp[5] ), .C(n2), .Z(n4)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i4610_3_lut.init = 16'hb2b2;
    LUT4 i4603_3_lut (.A(\mtime_out[0] ), .B(\mtimecmp[4] ), .C(cy_c), 
         .Z(n2)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i4603_3_lut.init = 16'hb2b2;
    LUT4 i4624_3_lut (.A(mtime_out[3]), .B(mtimecmp[7]), .C(n6), .Z(comparison[4])) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(72[29:71])
    defparam i4624_3_lut.init = 16'hb2b2;
    LUT4 time_pulse_I_0_2_lut_rep_708 (.A(n10573), .B(time_pulse_r), .Z(n31913)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(37[14:39])
    defparam time_pulse_I_0_2_lut_rep_708.init = 16'hdddd;
    PFUMX i28626 (.BLUT(n32084), .ALUT(n32085), .C0(mtime_out[2]), .Z(timer_interrupt_N_1954));
    tinyqv_counter i_mtime (.clk_c(clk_c), .n31980(n31980), .cy(cy), .mtime_out({mtime_out[3:1], 
            \mtime_out[0] }), .rst_reg_n(rst_reg_n), .instr_fetch_stopped(instr_fetch_stopped), 
            .instr_fetch_running_N_945(instr_fetch_running_N_945), .n28156(n28156), 
            .clk_c_enable_36(clk_c_enable_36), .address_ready(address_ready), 
            .is_store(is_store), .clk_c_enable_109(clk_c_enable_109), .\instr_data[1] (\instr_data[1] ), 
            .\instr_data_0__15__N_638[49] (\instr_data_0__15__N_638[49] ), 
            .n31876(n31876), .n31957(n31957), .n31946(n31946), .clk_c_enable_449(clk_c_enable_449), 
            .no_write_in_progress(no_write_in_progress), .clk_c_enable_157(clk_c_enable_157), 
            .n33488(n33488), .n31966(n31966), .\cycle_count_wide[3] (\cycle_count_wide[3] ), 
            .n31870(n31870), .clk_c_enable_233(clk_c_enable_233), .n31893(n31893), 
            .is_double_fault_r(is_double_fault_r), .mstatus_mte(mstatus_mte), 
            .n31841(n31841), .clk_c_enable_107(clk_c_enable_107), .\reg_access[3][2] (\reg_access[3][2] ), 
            .clk_c_enable_177(clk_c_enable_177), .\addr[2] (\addr[2] ), 
            .n32033(n32033), .is_timer_addr(is_timer_addr), .n8(n8), .n28028(n28028), 
            .n31748(n31748), .n26290(n26290), .mstatus_mie_N_1709(mstatus_mie_N_1709), 
            .n31878(n31878), .mstatus_mie_N_1707(mstatus_mie_N_1707), .n15604(n15604), 
            .clk_c_enable_161(clk_c_enable_161), .n31742(n31742), .n31737(n31737), 
            .clk_c_enable_347(clk_c_enable_347), .\instr_data[0] (\instr_data[0] ), 
            .\instr_data_0__15__N_638[0] (\instr_data_0__15__N_638[0] ), .n31884(n31884), 
            .n31872(n31872), .n31889(n31889), .data_out_slice({data_out_slice}), 
            .n31840(n31840)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/time.v(34[20] 42[6])
    
endmodule
//
// Verilog Description of module tinyqv_counter
//

module tinyqv_counter (clk_c, n31980, cy, mtime_out, rst_reg_n, instr_fetch_stopped, 
            instr_fetch_running_N_945, n28156, clk_c_enable_36, address_ready, 
            is_store, clk_c_enable_109, \instr_data[1] , \instr_data_0__15__N_638[49] , 
            n31876, n31957, n31946, clk_c_enable_449, no_write_in_progress, 
            clk_c_enable_157, n33488, n31966, \cycle_count_wide[3] , 
            n31870, clk_c_enable_233, n31893, is_double_fault_r, mstatus_mte, 
            n31841, clk_c_enable_107, \reg_access[3][2] , clk_c_enable_177, 
            \addr[2] , n32033, is_timer_addr, n8, n28028, n31748, 
            n26290, mstatus_mie_N_1709, n31878, mstatus_mie_N_1707, 
            n15604, clk_c_enable_161, n31742, n31737, clk_c_enable_347, 
            \instr_data[0] , \instr_data_0__15__N_638[0] , n31884, n31872, 
            n31889, data_out_slice, n31840) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    output n31980;
    output cy;
    output [3:0]mtime_out;
    input rst_reg_n;
    input instr_fetch_stopped;
    input instr_fetch_running_N_945;
    output n28156;
    input clk_c_enable_36;
    input address_ready;
    input is_store;
    output clk_c_enable_109;
    input \instr_data[1] ;
    output \instr_data_0__15__N_638[49] ;
    input n31876;
    input n31957;
    input n31946;
    output clk_c_enable_449;
    input no_write_in_progress;
    output clk_c_enable_157;
    input n33488;
    output n31966;
    input \cycle_count_wide[3] ;
    input n31870;
    output clk_c_enable_233;
    input n31893;
    input is_double_fault_r;
    input mstatus_mte;
    output n31841;
    output clk_c_enable_107;
    input \reg_access[3][2] ;
    output clk_c_enable_177;
    input \addr[2] ;
    input n32033;
    input is_timer_addr;
    input n8;
    input n28028;
    input n31748;
    output n26290;
    input mstatus_mie_N_1709;
    input n31878;
    output mstatus_mie_N_1707;
    input n15604;
    output clk_c_enable_161;
    input n31742;
    input n31737;
    output clk_c_enable_347;
    input \instr_data[0] ;
    output \instr_data_0__15__N_638[0] ;
    output n31884;
    input n31872;
    input n31889;
    input [3:0]data_out_slice;
    input n31840;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    wire [4:0]increment_result;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[16:32])
    
    wire n8835;
    wire [4:0]increment_result_3__N_1925;
    
    wire n31839, n31801;
    
    FD1S3IX register_2__48 (.D(increment_result[2]), .CK(clk_c), .CD(n31980), 
            .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result[1]), .CK(clk_c), .CD(n31980), 
            .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(increment_result[0]), .CK(clk_c), .CD(n31980), 
            .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3IX cy_51 (.D(increment_result_3__N_1925[4]), .CK(clk_c), .CD(n8835), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(register[10])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(register[9])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(register[8])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(mtime_out[3])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(register[10]), .CK(clk_c), .Q(mtime_out[2])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(register[9]), .CK(clk_c), .Q(mtime_out[1])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(register[8]), .CK(clk_c), .Q(mtime_out[0])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result[3]), .CK(clk_c), .CD(n31980), 
            .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=15, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=34, LSE_RLINE=42 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 rstn_I_0_1_lut_rep_775 (.A(rst_reg_n), .Z(n31980)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam rstn_I_0_1_lut_rep_775.init = 16'h5555;
    LUT4 i1_3_lut_3_lut (.A(rst_reg_n), .B(instr_fetch_stopped), .C(instr_fetch_running_N_945), 
         .Z(n28156)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(clk_c_enable_36), 
         .C(address_ready), .D(is_store), .Z(clk_c_enable_109)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hfddd;
    LUT4 i15292_2_lut_2_lut (.A(rst_reg_n), .B(\instr_data[1] ), .Z(\instr_data_0__15__N_638[49] )) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i15292_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_397 (.A(rst_reg_n), .B(n31876), 
         .C(n31957), .D(n31946), .Z(clk_c_enable_449)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_397.init = 16'h2000;
    LUT4 i16129_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(clk_c_enable_36), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_157)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i16129_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i3818_3_lut_rep_761_3_lut (.A(n33488), .B(no_write_in_progress), 
         .C(is_store), .Z(n31966)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3818_3_lut_rep_761_3_lut.init = 16'hd5d5;
    LUT4 i3845_4_lut_4_lut (.A(n33488), .B(\cycle_count_wide[3] ), .C(n31870), 
         .D(clk_c_enable_36), .Z(clk_c_enable_233)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3845_4_lut_4_lut.init = 16'hd555;
    LUT4 rstn_N_1579_I_0_2_lut_rep_636_4_lut_4_lut (.A(n33488), .B(n31893), 
         .C(is_double_fault_r), .D(mstatus_mte), .Z(n31841)) /* synthesis lut_function=((B (C+!(D))+!B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam rstn_N_1579_I_0_2_lut_rep_636_4_lut_4_lut.init = 16'hf5fd;
    LUT4 i3815_2_lut_2_lut (.A(rst_reg_n), .B(address_ready), .Z(clk_c_enable_107)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i3815_2_lut_2_lut.init = 16'hdddd;
    LUT4 i27832_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(\reg_access[3][2] ), 
         .C(no_write_in_progress), .D(is_store), .Z(clk_c_enable_177)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i27832_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i6240_2_lut_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(\addr[2] ), .C(n32033), 
         .D(is_timer_addr), .Z(n8835)) /* synthesis lut_function=(!(A (B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i6240_2_lut_3_lut_4_lut_4_lut.init = 16'h5755;
    LUT4 i1_4_lut_4_lut (.A(rst_reg_n), .B(n8), .C(n28028), .D(n31748), 
         .Z(n26290)) /* synthesis lut_function=((B (D)+!B (C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_4_lut_4_lut.init = 16'hff75;
    LUT4 i15345_3_lut_4_lut_4_lut (.A(rst_reg_n), .B(mstatus_mie_N_1709), 
         .C(n31878), .D(n31876), .Z(mstatus_mie_N_1707)) /* synthesis lut_function=((B ((D)+!C)+!B (D))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i15345_3_lut_4_lut_4_lut.init = 16'hff5d;
    LUT4 i27845_2_lut_4_lut_4_lut (.A(rst_reg_n), .B(n15604), .C(no_write_in_progress), 
         .D(is_store), .Z(clk_c_enable_161)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i27845_2_lut_4_lut_4_lut.init = 16'hc444;
    LUT4 i1_2_lut_3_lut_3_lut (.A(rst_reg_n), .B(n31742), .C(n31737), 
         .Z(clk_c_enable_347)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h7575;
    LUT4 i15259_2_lut_2_lut (.A(rst_reg_n), .B(\instr_data[0] ), .Z(\instr_data_0__15__N_638[0] )) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i15259_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_679_3_lut_3_lut (.A(n33488), .B(address_ready), .C(is_store), 
         .Z(n31884)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(221[13:18])
    defparam i1_2_lut_rep_679_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i4868_2_lut_3_lut_4_lut (.A(mtime_out[1]), .B(n31872), .C(mtime_out[3]), 
         .D(mtime_out[2]), .Z(increment_result_3__N_1925[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4868_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4854_2_lut_rep_634_3_lut (.A(mtime_out[0]), .B(n31889), .C(mtime_out[1]), 
         .Z(n31839)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4854_2_lut_rep_634_3_lut.init = 16'h8080;
    LUT4 i4861_2_lut_rep_596_3_lut_4_lut (.A(mtime_out[0]), .B(n31889), 
         .C(mtime_out[2]), .D(mtime_out[1]), .Z(n31801)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4861_2_lut_rep_596_3_lut_4_lut.init = 16'h8000;
    LUT4 increment_result_3__I_168_i3_4_lut (.A(mtime_out[2]), .B(data_out_slice[2]), 
         .C(n31840), .D(n31839), .Z(increment_result[2])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i3_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_168_i2_4_lut (.A(mtime_out[1]), .B(data_out_slice[1]), 
         .C(n31840), .D(n31872), .Z(increment_result[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i2_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_168_i1_4_lut (.A(mtime_out[0]), .B(data_out_slice[0]), 
         .C(n31840), .D(n31889), .Z(increment_result[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i1_4_lut.init = 16'hc5ca;
    LUT4 increment_result_3__I_168_i4_4_lut (.A(mtime_out[3]), .B(data_out_slice[3]), 
         .C(n31840), .D(n31801), .Z(increment_result[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[35:119])
    defparam increment_result_3__I_168_i4_4_lut.init = 16'hc5ca;
    
endmodule
//
// Verilog Description of module tinyqv_decoder
//

module tinyqv_decoder (n31850, n31441, n31860, n31402, n31774, n31869, 
            n31814, n31847, n31821, n31820, \instr[26] , n31837, 
            n31849, n31865, n31845, n10904, n31848, n31763, n31867, 
            n32, \mem_op_2__N_1114[1] , n31772, n31773, n31833, n31868, 
            n31823, n31853, n31194, n4269, n31852, n31851, n3265, 
            n31846, n31813, n31799, n31817, n3006, n31784, n31764, 
            n31838, \mem_op_de[1] , n31786, n31766, n31758, n31796, 
            n17976, n31790, n7, n10, n24, \alu_op_3__N_1170[2] , 
            n28366, \additional_mem_ops_2__N_1132[0] , n31795, n31864, 
            n8302, n31471, n41, n32_adj_3, n30, n4, n31762, n31816, 
            is_auipc_de, n29004, n31863, n31769, n31798, n22, \instr[27] , 
            n3365, n33488, n27746, n28332, n31791, n9894, n28006, 
            n17998, n31861, n31733, n27246, n31944, n4281, n29375, 
            \instr[16] , n2610, \instr[25] , n3367, n2169, n29048, 
            mem_op_increment_reg_de, n4263, n31732, n28898, n10068, 
            n4_adj_4, n13248, \instr[30] , n3, n28871, n26113, rst_reg_n, 
            n27850, is_alu_imm_de, n31831, is_jalr_N_1370, \instr[31] , 
            n5137, n5140, \instr[29] , n5123, \instr[24] , n5128, 
            n5127, n30771, n30770, n31728, \instr[28] , n5124, n30759, 
            n30760, \instr[19] , n30763, n29041, n29018, n29049, 
            n5125, n5136, n29043, n29020, n29045, n29026, n29047, 
            n29028, \instr[17] , n31682, n5139, n5138, n31818, n15, 
            alu_op_de, n30_adj_5, n31835, n31436, is_alu_reg_de, n31824, 
            n31822, is_store_de, is_lui_N_1365, is_lui_de, n157, n31815, 
            n3001, n8, n29215, is_load_de, n15_adj_6, n30_adj_7, 
            is_jal_de, is_jalr_de, clk_c_enable_325, n4285, n26, n29385, 
            n22_adj_8, n31760, n31714, n5147, n5152, n5148, n5145, 
            n31830, n31809, is_branch_de, n2998, n26202, n27956, 
            n28032, n28864, n28040, n27790, n27928, n26_adj_9, n27934, 
            n27688, n19, n27694, n28060, n28068, n31805, n28054, 
            n12, n2810, n2604, n2632, n27892, n27898, n27880, 
            n27886, n27904, n27910, n31785, \mem_op_de[2] , n27832, 
            n27838, n19_adj_10, n26478, n27868, n27874, n27818, 
            n27824, is_system_de) /* synthesis syn_module_defined=1 */ ;
    input n31850;
    input n31441;
    input n31860;
    input n31402;
    output n31774;
    input n31869;
    input n31814;
    input n31847;
    input n31821;
    input n31820;
    input \instr[26] ;
    input n31837;
    input n31849;
    input n31865;
    input n31845;
    output n10904;
    input n31848;
    output n31763;
    input n31867;
    output n32;
    input \mem_op_2__N_1114[1] ;
    output n31772;
    output n31773;
    input n31833;
    input n31868;
    input n31823;
    input n31853;
    output n31194;
    input n4269;
    input n31852;
    input n31851;
    output n3265;
    input n31846;
    output n31813;
    input n31799;
    input n31817;
    output n3006;
    output n31784;
    output n31764;
    input n31838;
    output \mem_op_de[1] ;
    output n31786;
    output n31766;
    output n31758;
    output n31796;
    output n17976;
    output n31790;
    input n7;
    output n10;
    output n24;
    input \alu_op_3__N_1170[2] ;
    input n28366;
    output \additional_mem_ops_2__N_1132[0] ;
    input n31795;
    input n31864;
    output n8302;
    output n31471;
    input n41;
    input n32_adj_3;
    output n30;
    input n4;
    output n31762;
    input n31816;
    output is_auipc_de;
    output n29004;
    input n31863;
    output n31769;
    output n31798;
    output n22;
    input \instr[27] ;
    output n3365;
    input n33488;
    output n27746;
    output n28332;
    output n31791;
    input n9894;
    output n28006;
    output n17998;
    input n31861;
    input n31733;
    output n27246;
    input n31944;
    input n4281;
    output n29375;
    input \instr[16] ;
    output n2610;
    input \instr[25] ;
    output n3367;
    input n2169;
    output n29048;
    output mem_op_increment_reg_de;
    output n4263;
    output n31732;
    output n28898;
    output n10068;
    input n4_adj_4;
    output n13248;
    input \instr[30] ;
    input n3;
    input n28871;
    output n26113;
    input rst_reg_n;
    output n27850;
    output is_alu_imm_de;
    input n31831;
    output is_jalr_N_1370;
    input \instr[31] ;
    output n5137;
    output n5140;
    input \instr[29] ;
    output n5123;
    input \instr[24] ;
    output n5128;
    output n5127;
    input n30771;
    output n30770;
    output n31728;
    input \instr[28] ;
    output n5124;
    input n30759;
    output n30760;
    input \instr[19] ;
    output n30763;
    input n29041;
    output n29018;
    output n29049;
    output n5125;
    output n5136;
    input n29043;
    output n29020;
    input n29045;
    output n29026;
    input n29047;
    output n29028;
    input \instr[17] ;
    output n31682;
    output n5139;
    output n5138;
    input n31818;
    output n15;
    output [3:0]alu_op_de;
    input n30_adj_5;
    input n31835;
    output n31436;
    output is_alu_reg_de;
    input n31824;
    input n31822;
    output is_store_de;
    input is_lui_N_1365;
    output is_lui_de;
    output n157;
    input n31815;
    output n3001;
    input n8;
    input n29215;
    output is_load_de;
    input n15_adj_6;
    input n30_adj_7;
    output is_jal_de;
    output is_jalr_de;
    input clk_c_enable_325;
    input n4285;
    input n26;
    output n29385;
    input n22_adj_8;
    input n31760;
    output n31714;
    output n5147;
    output n5152;
    output n5148;
    output n5145;
    input n31830;
    input n31809;
    output is_branch_de;
    output n2998;
    input n26202;
    output n27956;
    input n28032;
    input n28864;
    output n28040;
    output n27790;
    input n27928;
    input n26_adj_9;
    output n27934;
    input n27688;
    input n19;
    output n27694;
    input n28060;
    output n28068;
    input n31805;
    output n28054;
    output n12;
    input n2810;
    input n2604;
    output n2632;
    input n27892;
    output n27898;
    input n27880;
    output n27886;
    input n27904;
    output n27910;
    input n31785;
    output \mem_op_de[2] ;
    input n27832;
    output n27838;
    output n19_adj_10;
    output n26478;
    input n27868;
    output n27874;
    input n27818;
    output n27824;
    output is_system_de;
    
    
    wire n31487, n31486, n8899, n31442, n31443, n31401, n31403, 
        n31794, n19_c, n18578, n31771, n31781, n3_c;
    wire [3:0]alu_op_3__N_1337;
    
    wire n15_c, n27, alu_op_3__N_1181, n31779, n31782, n30_c, n7_c, 
        n31783, imm_31__N_1169, n9568, n9569, n28434;
    wire [3:0]n328;
    
    wire n15_adj_3117, n31793, n28464, n27216, n27129, mem_op_2__N_1384, 
        n31780, n8287;
    wire [3:0]alu_op_3__N_1107;
    
    wire n30653, n28458;
    wire [3:0]n155;
    
    wire n9023, n31765, n25010;
    wire [3:0]alu_op_3__N_1170;
    
    wire n9019, n31776, n28356, n31797, is_jal_N_1374, n26114, n29544;
    wire [2:0]additional_mem_ops_2__N_1129;
    
    wire n31757, n30657, n30656, n30655, n8300, n30654, n15_adj_3125, 
        n15_adj_3126, n18630;
    
    PFUMX i28481 (.BLUT(n31487), .ALUT(n31486), .C0(n31850), .Z(n8899));
    PFUMX i28459 (.BLUT(n31442), .ALUT(n31441), .C0(n31860), .Z(n31443));
    PFUMX i28433 (.BLUT(n31402), .ALUT(n31401), .C0(n31774), .Z(n31403));
    LUT4 i16006_4_lut_4_lut (.A(n31869), .B(n31814), .C(n31794), .D(n19_c), 
         .Z(n18578)) /* synthesis lut_function=(A (C)+!A !(B+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i16006_4_lut_4_lut.init = 16'hb1a0;
    LUT4 i25_2_lut_rep_566_4_lut (.A(n31847), .B(n31821), .C(n31820), 
         .D(\instr[26] ), .Z(n31771)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(67[27:51])
    defparam i25_2_lut_rep_566_4_lut.init = 16'h0200;
    LUT4 i8286_3_lut_4_lut (.A(n31837), .B(n31849), .C(n31865), .D(n31845), 
         .Z(n10904)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i8286_3_lut_4_lut.init = 16'h10f0;
    LUT4 i27790_2_lut_rep_558_4_lut (.A(n31849), .B(n31837), .C(n31848), 
         .D(n31865), .Z(n31763)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i27790_2_lut_rep_558_4_lut.init = 16'h0001;
    LUT4 i53_4_lut_4_lut (.A(n31867), .B(n31860), .C(n31781), .D(n31869), 
         .Z(n32)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i53_4_lut_4_lut.init = 16'hd1c0;
    LUT4 instr_1__I_0_133_Mux_1_i3_4_lut_4_lut_4_lut (.A(n31867), .B(\mem_op_2__N_1114[1] ), 
         .C(n31772), .D(n31773), .Z(n3_c)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam instr_1__I_0_133_Mux_1_i3_4_lut_4_lut_4_lut.init = 16'h505c;
    LUT4 i15842_4_lut_4_lut (.A(n31867), .B(n31845), .C(n31833), .D(alu_op_3__N_1337[2]), 
         .Z(n15_c)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i15842_4_lut_4_lut.init = 16'hd0c0;
    LUT4 instr_13__bdd_3_lut_28405_4_lut_4_lut (.A(n31867), .B(n31868), 
         .C(n31823), .D(n31853), .Z(n31194)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam instr_13__bdd_3_lut_28405_4_lut_4_lut.init = 16'h0400;
    LUT4 mux_2091_i2_4_lut_4_lut (.A(n31867), .B(n4269), .C(n31852), .D(n31851), 
         .Z(n3265)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam mux_2091_i2_4_lut_4_lut.init = 16'h7340;
    LUT4 i42_4_lut_4_lut (.A(n31867), .B(n31845), .C(n31869), .D(n31860), 
         .Z(n27)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i42_4_lut_4_lut.init = 16'h404a;
    LUT4 instr_6__I_0_142_i10_2_lut_3_lut (.A(n31852), .B(n31846), .C(n31813), 
         .Z(alu_op_3__N_1181)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam instr_6__I_0_142_i10_2_lut_3_lut.init = 16'h0808;
    LUT4 i1_3_lut_rep_608 (.A(n31850), .B(n31851), .C(n31847), .Z(n31813)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_rep_608.init = 16'hf7f7;
    LUT4 instr_6__I_0_157_i9_2_lut_rep_574_4_lut (.A(n31850), .B(n31851), 
         .C(n31847), .D(n31820), .Z(n31779)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam instr_6__I_0_157_i9_2_lut_rep_574_4_lut.init = 16'hfff7;
    LUT4 i1_3_lut_rep_577_4_lut (.A(n31845), .B(n31868), .C(n31867), .D(n31869), 
         .Z(n31782)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i1_3_lut_rep_577_4_lut.init = 16'hfbff;
    LUT4 i15841_2_lut_3_lut_4_lut (.A(n31845), .B(n31868), .C(n31867), 
         .D(n31869), .Z(n30_c)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i15841_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 instr_1__I_0_139_i7_4_lut (.A(n31799), .B(n31848), .C(n31868), 
         .D(n31817), .Z(n7_c)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam instr_1__I_0_139_i7_4_lut.init = 16'h0a3a;
    LUT4 mux_2063_i9_3_lut_4_lut_4_lut (.A(n31847), .B(n31846), .C(n31868), 
         .D(n31852), .Z(n3006)) /* synthesis lut_function=(A (B+((D)+!C))+!A (C (D))) */ ;
    defparam mux_2063_i9_3_lut_4_lut_4_lut.init = 16'hfa8a;
    LUT4 i27712_2_lut_rep_579_3_lut (.A(n31847), .B(n31846), .C(n31852), 
         .Z(n31784)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i27712_2_lut_rep_579_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_578_3_lut (.A(n31846), .B(n31852), .C(n31847), .Z(n31783)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(65[27:51])
    defparam i1_2_lut_rep_578_3_lut.init = 16'hdfdf;
    LUT4 i1_2_lut_rep_559_3_lut_4_lut (.A(n31846), .B(n31852), .C(n31850), 
         .D(n31847), .Z(n31764)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(65[27:51])
    defparam i1_2_lut_rep_559_3_lut_4_lut.init = 16'hfdff;
    LUT4 instr_6__I_0_127_i10_2_lut_3_lut_4_lut (.A(n31846), .B(n31852), 
         .C(n31821), .D(n31847), .Z(imm_31__N_1169)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(65[27:51])
    defparam instr_6__I_0_127_i10_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i6968_3_lut_4_lut_4_lut_4_lut_4_lut_4_lut (.A(n31867), .B(n31845), 
         .C(n31868), .D(n31838), .Z(n9568)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A ((D)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i6968_3_lut_4_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h00ce;
    LUT4 i27843_2_lut_rep_576_3_lut_4_lut (.A(n31867), .B(n31845), .C(n31868), 
         .D(n31869), .Z(n31781)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i27843_2_lut_rep_576_3_lut_4_lut.init = 16'h0001;
    LUT4 i15849_2_lut_3_lut (.A(n31869), .B(n31860), .C(n9569), .Z(\mem_op_de[1] )) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/cpu.v(73[20] 98[6])
    defparam i15849_2_lut_3_lut.init = 16'hd0d0;
    LUT4 i1_2_lut_rep_581_3_lut (.A(n31846), .B(n31852), .C(n31847), .Z(n31786)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam i1_2_lut_rep_581_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n31846), .B(n31852), .C(n8899), .D(n31813), 
         .Z(n28434)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i27653_3_lut_rep_589_4_lut (.A(n31846), .B(n31852), .C(n31821), 
         .D(n31847), .Z(n31794)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam i27653_3_lut_rep_589_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_561_3_lut_4_lut (.A(n31846), .B(n31852), .C(n31821), 
         .D(n31847), .Z(n31766)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam i1_2_lut_rep_561_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_553_3_lut_4_lut_4_lut (.A(n31851), .B(n31850), .C(n31783), 
         .D(n31786), .Z(n31758)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i1_2_lut_rep_553_3_lut_4_lut_4_lut.init = 16'hfcdc;
    LUT4 i1_2_lut_rep_591_3_lut_4_lut (.A(n31868), .B(n31869), .C(n31867), 
         .D(n31845), .Z(n31796)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i1_2_lut_rep_591_3_lut_4_lut.init = 16'h2000;
    LUT4 i15409_2_lut_3_lut_4_lut (.A(n31849), .B(n31848), .C(n31869), 
         .D(n31853), .Z(n17976)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i15409_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i15843_4_lut_4_lut_4_lut (.A(n31849), .B(n31848), .C(n328[1]), 
         .D(n31782), .Z(n15_adj_3117)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!B))) */ ;
    defparam i15843_4_lut_4_lut_4_lut.init = 16'h00c4;
    LUT4 i15305_2_lut_rep_588_3_lut (.A(n31849), .B(n31848), .C(n31853), 
         .Z(n31793)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i15305_2_lut_rep_588_3_lut.init = 16'hf7f7;
    LUT4 i601_2_lut_rep_585_3_lut (.A(n31849), .B(n31848), .C(n31853), 
         .Z(n31790)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i601_2_lut_rep_585_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_369 (.A(n31849), .B(n31848), .C(n7), 
         .D(n31853), .Z(alu_op_3__N_1337[2])) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_369.init = 16'hfff7;
    LUT4 i1_2_lut_3_lut (.A(n31851), .B(n31850), .C(n31860), .Z(n28464)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(218[25] 223[32])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 is_jalr_N_1372_bdd_2_lut_3_lut (.A(n31845), .B(n31868), .C(n31867), 
         .Z(n31442)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam is_jalr_N_1372_bdd_2_lut_3_lut.init = 16'h7070;
    LUT4 i2_2_lut_3_lut (.A(n31845), .B(n31868), .C(n31867), .Z(n10)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(n31845), .B(n31868), .C(n31867), 
         .D(n31838), .Z(n27216)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i37_3_lut_3_lut (.A(n31845), .B(n31868), .C(n31867), .Z(n24)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;
    defparam i37_3_lut_3_lut.init = 16'h7a7a;
    LUT4 i1_3_lut (.A(n8899), .B(\alu_op_3__N_1170[2] ), .C(n31869), .Z(n27129)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i597_4_lut (.A(n31850), .B(mem_op_2__N_1384), .C(n31780), .D(n28366), 
         .Z(\additional_mem_ops_2__N_1132[0] )) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(93[13] 98[16])
    defparam i597_4_lut.init = 16'h3733;
    LUT4 i15299_4_lut (.A(n31853), .B(n8899), .C(n31867), .D(n8287), 
         .Z(alu_op_3__N_1107[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(83[18] 85[91])
    defparam i15299_4_lut.init = 16'hc088;
    LUT4 is_alu_imm_N_1367_bdd_2_lut_28247_3_lut_4_lut (.A(n31850), .B(n31851), 
         .C(n31847), .D(n31820), .Z(n30653)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam is_alu_imm_N_1367_bdd_2_lut_28247_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_370 (.A(n31850), .B(n31851), .C(n31853), .Z(n28458)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam i1_2_lut_3_lut_adj_370.init = 16'hfefe;
    LUT4 i5724_4_lut_4_lut (.A(n31869), .B(n31795), .C(n31864), .D(\additional_mem_ops_2__N_1132[0] ), 
         .Z(n8302)) /* synthesis lut_function=(A (D)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i5724_4_lut_4_lut.init = 16'hea40;
    LUT4 n15_bdd_3_lut_3_lut (.A(n31869), .B(n31868), .C(n31845), .Z(n31471)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam n15_bdd_3_lut_3_lut.init = 16'h1414;
    LUT4 i6424_4_lut_4_lut (.A(n31869), .B(n155[3]), .C(n30_c), .D(n28434), 
         .Z(n9023)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i6424_4_lut_4_lut.init = 16'hd850;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n31869), .B(n41), .C(n32_adj_3), .D(n31867), 
         .Z(n30)) /* synthesis lut_function=(!(A+!(B+!((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h4454;
    LUT4 i1_4_lut (.A(n31765), .B(n4), .C(n31849), .D(n31774), .Z(n25010)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i1_4_lut.init = 16'h5044;
    LUT4 i6420_4_lut_4_lut (.A(n31869), .B(n8899), .C(n30_c), .D(alu_op_3__N_1170[1]), 
         .Z(n9019)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i6420_4_lut_4_lut.init = 16'hd850;
    LUT4 i26329_2_lut_rep_575_3_lut (.A(n31852), .B(n31846), .C(n31847), 
         .Z(n31780)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i26329_2_lut_rep_575_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_571_3_lut (.A(n31852), .B(n31846), .C(n31847), .Z(n31776)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_571_3_lut.init = 16'h1010;
    LUT4 i26331_2_lut_rep_557_3_lut_4_lut (.A(n31852), .B(n31846), .C(n7), 
         .D(n31847), .Z(n31762)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26331_2_lut_rep_557_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_371 (.A(n7), .B(n31816), .C(n31838), .D(n31847), 
         .Z(is_auipc_de)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_371.init = 16'h1000;
    LUT4 i26445_3_lut_4_lut (.A(n31852), .B(n31846), .C(n31845), .D(n7), 
         .Z(n29004)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26445_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut (.A(n31852), .B(n31846), .C(n31847), .D(n31853), 
         .Z(n28356)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_592_3_lut (.A(n31864), .B(n31863), .C(n31849), .Z(n31797)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_rep_592_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_564_3_lut_4_lut (.A(n31864), .B(n31863), .C(n31865), 
         .D(n31849), .Z(n31769)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_rep_564_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_3_lut_rep_593_4_lut (.A(n31864), .B(n31863), .C(n31848), .D(n31849), 
         .Z(n31798)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_3_lut_rep_593_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_4_lut_4_lut_adj_372 (.A(n31860), .B(n31867), .C(n31869), 
         .D(n31845), .Z(is_jal_N_1374)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_4_lut_4_lut_4_lut_adj_372.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_373 (.A(n31860), .B(n26114), .C(n31869), 
         .D(n31867), .Z(n22)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i1_4_lut_4_lut_4_lut_adj_373.init = 16'h005c;
    LUT4 i6904_3_lut_4_lut (.A(n31869), .B(n31860), .C(\instr[27] ), .D(n31865), 
         .Z(n3365)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i6904_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_adj_374 (.A(n31869), .B(n31860), .C(n33488), .Z(n27746)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_374.init = 16'h8080;
    LUT4 i1_3_lut_4_lut_adj_375 (.A(n31869), .B(n31860), .C(n27), .D(n31868), 
         .Z(n28332)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !((D)+!C)) */ ;
    defparam i1_3_lut_4_lut_adj_375.init = 16'h88f8;
    LUT4 i27766_2_lut_rep_586_3_lut (.A(n31869), .B(n31860), .C(n33488), 
         .Z(n31791)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i27766_2_lut_rep_586_3_lut.init = 16'h8f8f;
    LUT4 i1_2_lut_3_lut_4_lut_adj_376 (.A(n31869), .B(n31860), .C(n9894), 
         .D(n33488), .Z(n28006)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_376.init = 16'h0700;
    LUT4 i16027_2_lut_2_lut_3_lut_4_lut (.A(n31869), .B(n31860), .C(n31868), 
         .D(n31845), .Z(n17998)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;
    defparam i16027_2_lut_2_lut_3_lut_4_lut.init = 16'h7770;
    LUT4 i1_3_lut_3_lut_4_lut (.A(n31869), .B(n31860), .C(n31861), .D(n31733), 
         .Z(n27246)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i27902_3_lut_4_lut (.A(n31869), .B(n31860), .C(n31944), .D(n4281), 
         .Z(n29375)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;
    defparam i27902_3_lut_4_lut.init = 16'hff08;
    LUT4 i15577_2_lut_3_lut (.A(n31869), .B(n31860), .C(\instr[16] ), 
         .Z(n2610)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i15577_2_lut_3_lut.init = 16'h8080;
    LUT4 i6900_3_lut_4_lut (.A(n31869), .B(n31860), .C(\instr[25] ), .D(n31853), 
         .Z(n3367)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam i6900_3_lut_4_lut.init = 16'hf780;
    LUT4 i168_2_lut_rep_567_2_lut_3_lut (.A(n31869), .B(n31860), .C(n31845), 
         .Z(n31772)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i168_2_lut_rep_567_2_lut_3_lut.init = 16'h7070;
    LUT4 i167_2_lut_rep_569_2_lut_3_lut (.A(n31869), .B(n31860), .C(n31868), 
         .Z(n31774)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i167_2_lut_rep_569_2_lut_3_lut.init = 16'h7070;
    LUT4 mux_1538_i11_rep_102_3_lut_3_lut_4_lut (.A(n31869), .B(n31860), 
         .C(n2169), .D(n31864), .Z(n29048)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_1538_i11_rep_102_3_lut_3_lut_4_lut.init = 16'hf780;
    LUT4 i169_2_lut_rep_568_2_lut_3_lut (.A(n31869), .B(n31860), .C(n31867), 
         .Z(n31773)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i169_2_lut_rep_568_2_lut_3_lut.init = 16'h7070;
    LUT4 i15310_2_lut_2_lut_3_lut (.A(n31869), .B(n31860), .C(mem_op_2__N_1384), 
         .Z(mem_op_increment_reg_de)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i15310_2_lut_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i27781_2_lut_3_lut_3_lut_4_lut_3_lut (.A(n31869), .B(n31860), .C(n31868), 
         .Z(n29544)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i27781_2_lut_3_lut_3_lut_4_lut_3_lut.init = 16'h7474;
    LUT4 i6898_rep_527_4_lut (.A(n31869), .B(n31860), .C(n31733), .D(n4263), 
         .Z(n31732)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam i6898_rep_527_4_lut.init = 16'h08f8;
    LUT4 i26340_2_lut_3_lut (.A(n31869), .B(n31860), .C(n31845), .Z(n28898)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i26340_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i2_2_lut_3_lut_adj_377 (.A(n31869), .B(n31860), .C(n4281), .Z(n10068)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i2_2_lut_3_lut_adj_377.init = 16'hf8f8;
    LUT4 i5542_2_lut_rep_560_2_lut_3_lut_4_lut (.A(n31869), .B(n31860), 
         .C(n31845), .D(n31867), .Z(n31765)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;
    defparam i5542_2_lut_rep_560_2_lut_3_lut_4_lut.init = 16'h7770;
    LUT4 i5_3_lut_3_lut_4_lut (.A(n31869), .B(n31860), .C(additional_mem_ops_2__N_1129[2]), 
         .D(n4_adj_4), .Z(n13248)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;
    defparam i5_3_lut_3_lut_4_lut.init = 16'h708f;
    LUT4 mux_29_i2_4_lut (.A(n31845), .B(n31771), .C(n31779), .D(n31867), 
         .Z(alu_op_3__N_1170[1])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[18] 85[91])
    defparam mux_29_i2_4_lut.init = 16'hfaca;
    LUT4 i15572_4_lut (.A(\instr[30] ), .B(n31771), .C(n31851), .D(n3), 
         .Z(n155[3])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(85[18:91])
    defparam i15572_4_lut.init = 16'hecee;
    LUT4 i1_4_lut_adj_378 (.A(n28871), .B(n7), .C(n31852), .D(n31860), 
         .Z(n26113)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_378.init = 16'h0100;
    LUT4 i1_3_lut_rep_552_4_lut (.A(n7), .B(n31780), .C(n31868), .D(n31817), 
         .Z(n31757)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_rep_552_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_adj_379 (.A(n31865), .B(n31798), .C(n26113), .Z(n26114)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_3_lut_adj_379.init = 16'he0e0;
    LUT4 is_alu_imm_N_1367_bdd_3_lut_28248 (.A(n31845), .B(n31868), .C(n31867), 
         .Z(n30657)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam is_alu_imm_N_1367_bdd_3_lut_28248.init = 16'h0101;
    LUT4 i1_3_lut_4_lut_adj_380 (.A(n31865), .B(n31798), .C(rst_reg_n), 
         .D(n9894), .Z(n27850)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_3_lut_4_lut_adj_380.init = 16'h0010;
    LUT4 n30657_bdd_3_lut (.A(n30657), .B(n30656), .C(n31869), .Z(is_alu_imm_de)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30657_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_381 (.A(n31865), .B(n31798), .C(n31757), 
         .D(n31831), .Z(is_jalr_N_1370)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(278[29:45])
    defparam i1_2_lut_3_lut_4_lut_adj_381.init = 16'he000;
    LUT4 mux_3131_i16_3_lut_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n31868), .Z(n5137)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3131_i16_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_3131_i13_3_lut_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n31853), .Z(n5140)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3131_i13_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_3131_i30_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[29] ), 
         .D(\instr[31] ), .Z(n5123)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_3131_i30_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_3131_i25_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[24] ), 
         .D(\instr[31] ), .Z(n5128)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_3131_i25_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_3131_i26_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[25] ), 
         .D(\instr[31] ), .Z(n5127)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_3131_i26_3_lut_4_lut.init = 16'hfe10;
    LUT4 n30769_bdd_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n30771), .Z(n30770)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam n30769_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i7166_3_lut_rep_523_4_lut (.A(n31850), .B(n31783), .C(n4281), 
         .D(n31838), .Z(n31728)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i7166_3_lut_rep_523_4_lut.init = 16'hefe0;
    LUT4 mux_3131_i29_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[28] ), 
         .D(\instr[31] ), .Z(n5124)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_3131_i29_3_lut_4_lut.init = 16'hfe10;
    PFUMX i28003 (.BLUT(n30655), .ALUT(n30653), .C0(n31860), .Z(n30656));
    LUT4 n30759_bdd_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n30759), .Z(n30760)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam n30759_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n4275_bdd_3_lut_28056_4_lut (.A(n31850), .B(n31783), .C(\instr[19] ), 
         .D(\instr[31] ), .Z(n30763)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam n4275_bdd_3_lut_28056_4_lut.init = 16'hfe10;
    LUT4 mux_1538_i5_rep_72_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n29041), .Z(n29018)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1538_i5_rep_72_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1538_i11_rep_103_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n2169), .Z(n29049)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1538_i11_rep_103_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_3131_i28_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[27] ), 
         .D(\instr[31] ), .Z(n5125)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_3131_i28_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_3131_i17_3_lut_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(\instr[16] ), .Z(n5136)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3131_i17_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1538_i6_rep_74_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n29043), .Z(n29020)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1538_i6_rep_74_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1538_i7_rep_80_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n29045), .Z(n29026)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1538_i7_rep_80_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1538_i8_rep_82_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n29047), .Z(n29028)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_1538_i8_rep_82_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n31681_bdd_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(\instr[17] ), .Z(n31682)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam n31681_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_3131_i14_3_lut_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n31867), .Z(n5139)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3131_i14_3_lut_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_3131_i15_3_lut_3_lut_4_lut (.A(n31850), .B(n31783), .C(\instr[31] ), 
         .D(n31845), .Z(n5138)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_3131_i15_3_lut_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i6969 (.BLUT(n3_c), .ALUT(n9568), .C0(n29544), .Z(n9569));
    PFUMX instr_1__I_0_133_Mux_0_i15 (.BLUT(n25010), .ALUT(n27216), .C0(n31818), 
          .Z(n15)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    PFUMX i6421 (.BLUT(n15_adj_3117), .ALUT(n9019), .C0(n31860), .Z(alu_op_de[1]));
    PFUMX i5722 (.BLUT(alu_op_3__N_1107[0]), .ALUT(n30_adj_5), .C0(n31835), 
          .Z(n8300));
    LUT4 n31194_bdd_3_lut_4_lut (.A(n31865), .B(n31797), .C(n31867), .D(n31868), 
         .Z(n31436)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(282[33:52])
    defparam n31194_bdd_3_lut_4_lut.init = 16'h0020;
    LUT4 is_alu_imm_N_1367_bdd_3_lut_28005_4_lut (.A(n31865), .B(n31797), 
         .C(n31867), .D(n31845), .Z(n30654)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(282[33:52])
    defparam is_alu_imm_N_1367_bdd_3_lut_28005_4_lut.init = 16'h2f0f;
    PFUMX i6423 (.BLUT(n15_c), .ALUT(n27129), .C0(n31860), .Z(alu_op_de[2]));
    PFUMX i6425 (.BLUT(n15_adj_3125), .ALUT(n9023), .C0(n31860), .Z(alu_op_de[3]));
    PFUMX i16007 (.BLUT(n15_adj_3126), .ALUT(n18578), .C0(n31860), .Z(is_alu_reg_de));
    LUT4 i5723_4_lut (.A(alu_op_3__N_1337[0]), .B(n8300), .C(n31860), 
         .D(n31782), .Z(alu_op_de[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i5723_4_lut.init = 16'hc0ca;
    LUT4 i15304_4_lut (.A(n31824), .B(n31823), .C(n31784), .D(n31853), 
         .Z(alu_op_3__N_1337[0])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B+!(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(203[30] 224[24])
    defparam i15304_4_lut.init = 16'hcfee;
    LUT4 is_store_I_0_4_lut (.A(n18630), .B(n31766), .C(n31838), .D(n31822), 
         .Z(is_store_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam is_store_I_0_4_lut.init = 16'h3a30;
    LUT4 i16056_4_lut (.A(n31860), .B(n31845), .C(n31867), .D(n31848), 
         .Z(n18630)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i16056_4_lut.init = 16'hcdcc;
    PFUMX is_lui_I_0 (.BLUT(is_lui_N_1365), .ALUT(imm_31__N_1169), .C0(n31838), 
          .Z(is_lui_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 mux_28_i3_3_lut_4_lut (.A(\instr[26] ), .B(n31794), .C(\instr[27] ), 
         .D(n31845), .Z(n157)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(84[22:45])
    defparam mux_28_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i15840_4_lut_4_lut (.A(n31782), .B(n28458), .C(n31849), .D(n31848), 
         .Z(n15_adj_3125)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i15840_4_lut_4_lut.init = 16'h1050;
    LUT4 mux_2063_i10_rep_93_3_lut_4_lut (.A(n31852), .B(n31815), .C(n31868), 
         .D(n31853), .Z(n3001)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(205[25] 214[32])
    defparam mux_2063_i10_rep_93_3_lut_4_lut.init = 16'hefe0;
    PFUMX i21 (.BLUT(n7_c), .ALUT(n8), .C0(n29215), .Z(is_load_de));
    PFUMX instr_1__I_0_138_Mux_2_i31 (.BLUT(n15_adj_6), .ALUT(n30_adj_7), 
          .C0(n31860), .Z(additional_mem_ops_2__N_1129[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    PFUMX is_jal_I_0 (.BLUT(is_jal_N_1374), .ALUT(alu_op_3__N_1181), .C0(n31838), 
          .Z(is_jal_de)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=73, LSE_RLINE=98 */ ;
    LUT4 i5709_2_lut_3_lut_4_lut (.A(n31820), .B(n31813), .C(n31794), 
         .D(\instr[26] ), .Z(n8287)) /* synthesis lut_function=(A (C (D))+!A ((C (D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(69[27:51])
    defparam i5709_2_lut_3_lut_4_lut.init = 16'hf111;
    LUT4 i15955_2_lut_4_lut (.A(n31869), .B(n31814), .C(n31867), .D(n31793), 
         .Z(n15_adj_3126)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(121[13] 320[20])
    defparam i15955_2_lut_4_lut.init = 16'h0002;
    LUT4 is_jalr_I_0_4_lut (.A(is_jalr_N_1370), .B(n31816), .C(n31838), 
         .D(n31813), .Z(is_jalr_de)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam is_jalr_I_0_4_lut.init = 16'h0a3a;
    LUT4 i27895_2_lut_3_lut_4_lut (.A(n31838), .B(clk_c_enable_325), .C(n4285), 
         .D(n26), .Z(n29385)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i27895_2_lut_3_lut_4_lut.init = 16'hfbff;
    LUT4 i15439_2_lut_rep_509_3_lut_4_lut_4_lut (.A(n31838), .B(clk_c_enable_325), 
         .C(n22_adj_8), .D(n31760), .Z(n31714)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(62[13:32])
    defparam i15439_2_lut_rep_509_3_lut_4_lut_4_lut.init = 16'hffbf;
    LUT4 i15686_2_lut_3_lut_4_lut (.A(n31847), .B(n31816), .C(\instr[25] ), 
         .D(n31850), .Z(n5147)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i15686_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i15407_2_lut_3_lut_4_lut (.A(n31847), .B(n31816), .C(n31864), 
         .D(n31850), .Z(n5152)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i15407_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i15685_2_lut_3_lut_4_lut (.A(n31847), .B(n31816), .C(n31848), 
         .D(n31850), .Z(n5148)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i15685_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i15688_2_lut_3_lut_4_lut (.A(n31847), .B(n31816), .C(\instr[27] ), 
         .D(n31850), .Z(n5145)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(68[27:51])
    defparam i15688_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 is_branch_I_0_4_lut (.A(n31830), .B(n31779), .C(n31838), .D(n31809), 
         .Z(is_branch_de)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam is_branch_I_0_4_lut.init = 16'h3a30;
    LUT4 mux_2063_i17_3_lut_4_lut (.A(n31852), .B(n31815), .C(n31868), 
         .D(n31853), .Z(n2998)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_2063_i17_3_lut_4_lut.init = 16'h4f40;
    LUT4 i1_4_lut_adj_382 (.A(n31852), .B(n26202), .C(n31846), .D(n31850), 
         .Z(n4263)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_382.init = 16'h0400;
    LUT4 mux_61_i2_3_lut_4_lut (.A(n31852), .B(n31815), .C(n31853), .D(n31850), 
         .Z(n328[1])) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(206[29:35])
    defparam mux_61_i2_3_lut_4_lut.init = 16'hbfb0;
    LUT4 additional_mem_ops_2__N_1132_0__bdd_3_lut (.A(n31848), .B(n31849), 
         .C(n31850), .Z(n31401)) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam additional_mem_ops_2__N_1132_0__bdd_3_lut.init = 16'h1515;
    LUT4 i15600_2_lut_3_lut_4_lut (.A(n31847), .B(n31820), .C(n31867), 
         .D(n7), .Z(n19_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(63[27:51])
    defparam i15600_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_383 (.A(n31867), .B(n31821), .C(n31845), .D(n28356), 
         .Z(mem_op_2__N_1384)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut_adj_383.init = 16'hffdf;
    LUT4 i1_4_lut_4_lut (.A(n31838), .B(n33488), .C(n31853), .D(n9894), 
         .Z(n27956)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_384 (.A(n31838), .B(n28032), .C(n28864), .D(n9894), 
         .Z(n28040)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_384.init = 16'h0004;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n31838), .B(n31818), .C(n31831), .D(n31868), 
         .Z(n27790)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h1000;
    LUT4 i1_4_lut_4_lut_adj_385 (.A(n31838), .B(n27928), .C(n9894), .D(n26_adj_9), 
         .Z(n27934)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_385.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_386 (.A(n31838), .B(n27688), .C(n9894), .D(n19), 
         .Z(n27694)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_386.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_387 (.A(n31838), .B(n28060), .C(n28864), .D(n9894), 
         .Z(n28068)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_387.init = 16'h0004;
    LUT4 i1_4_lut_4_lut_adj_388 (.A(n31838), .B(n31805), .C(n28864), .D(n9894), 
         .Z(n28054)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_388.init = 16'h0004;
    LUT4 instr_3__bdd_4_lut (.A(n31852), .B(n31846), .C(n31851), .D(n31847), 
         .Z(n31487)) /* synthesis lut_function=(A+(B (C+!(D))+!B (D))) */ ;
    defparam instr_3__bdd_4_lut.init = 16'hfbee;
    LUT4 instr_3__bdd_3_lut (.A(n31846), .B(n31851), .C(n31847), .Z(n31486)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam instr_3__bdd_3_lut.init = 16'hf7f7;
    LUT4 i2_2_lut_3_lut_4_lut_4_lut (.A(n31838), .B(n31817), .C(n31786), 
         .D(n7), .Z(n12)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i2_2_lut_3_lut_4_lut_4_lut.init = 16'hfff4;
    LUT4 mux_1879_i3_4_lut_4_lut (.A(n31838), .B(n2810), .C(\instr[17] ), 
         .D(n2604), .Z(n2632)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;
    defparam mux_1879_i3_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i1_4_lut_4_lut_adj_389 (.A(n31838), .B(n27892), .C(n9894), .D(n26_adj_9), 
         .Z(n27898)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_389.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_390 (.A(n31838), .B(n27880), .C(n9894), .D(n26_adj_9), 
         .Z(n27886)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_390.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_391 (.A(n31838), .B(n27904), .C(n9894), .D(n26_adj_9), 
         .Z(n27910)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_391.init = 16'h0400;
    LUT4 i1_3_lut_4_lut_4_lut_adj_392 (.A(n31838), .B(n31403), .C(n31785), 
         .D(n31817), .Z(\mem_op_de[2] )) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C+(D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_392.init = 16'h080c;
    LUT4 i1_4_lut_4_lut_adj_393 (.A(n31838), .B(n27832), .C(n9894), .D(n26_adj_9), 
         .Z(n27838)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_393.init = 16'h0400;
    LUT4 i1_3_lut_4_lut_4_lut_adj_394 (.A(n31838), .B(n31818), .C(n31848), 
         .D(n31867), .Z(n19_adj_10)) /* synthesis lut_function=(A (B+(C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_394.init = 16'ha8fc;
    LUT4 i23975_2_lut_3_lut_4_lut_4_lut (.A(n31838), .B(n31867), .C(n31818), 
         .D(n31831), .Z(n26478)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i23975_2_lut_3_lut_4_lut_4_lut.init = 16'hfff4;
    LUT4 i1_4_lut_4_lut_adj_395 (.A(n31838), .B(n27868), .C(n9894), .D(n26_adj_9), 
         .Z(n27874)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_395.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_396 (.A(n31838), .B(n27818), .C(n9894), .D(n26_adj_9), 
         .Z(n27824)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_4_lut_adj_396.init = 16'h0400;
    LUT4 n30654_bdd_3_lut_4_lut_4_lut (.A(n31817), .B(n30654), .C(n31868), 
         .D(n31793), .Z(n30655)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam n30654_bdd_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i25_4_lut (.A(n31443), .B(n28464), .C(n31869), .D(n31776), 
         .Z(is_system_de)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/decode.v(103[18] 321[12])
    defparam i25_4_lut.init = 16'hca0a;
    
endmodule
//
// Verilog Description of module tinyqv_core
//

module tinyqv_core (clk_c, n31841, n31980, clk_c_enable_234, counter_hi, 
            n92, n18324, instr_complete_N_1647, clk_c_enable_449, \ui_in_sync[0] , 
            mstatus_mte, \imm[10] , n31744, n31738, n27838, n31742, 
            n26648, \imm[1] , n27934, n26764, n27874, n26794, data_rs1, 
            n27810, n2804, n27886, n26788, n28020, n2498, n27960, 
            n3402, n28068, n26807, n28080, n26889, n27672, n31758, 
            n31733, n27862, n2592, n9894, n27728, n27734, \next_pc_for_core[7] , 
            \next_pc_for_core[3] , n27910, n26776, \next_pc_for_core[23] , 
            \next_pc_for_core[19] , n28116, n26871, n27946, n31735, 
            \next_pc_for_core[15] , \next_pc_for_core[11] , n27922, n26770, 
            \alu_op[0] , \alu_op[3] , \alu_op[1] , \alu_op_in[2] , n29006, 
            n28881, n27738, n27744, n27898, n26782, n30947, n31853, 
            n30949, n27790, n12, n27796, n28128, n26827, n28140, 
            n26905, n28054, n26814, n31894, n31875, n1160, load_done, 
            clk_c_enable_249, n8289, \imm[2] , \imm[6] , clk_c_enable_233, 
            n27576, n31720, n26800, n31838, is_jalr_N_1370, n27724, 
            n28040, n26821, stall_core, clk_c_enable_36, n28204, n26993, 
            is_double_fault_r, n31893, n31878, n28092, n26883, n28104, 
            n26877, n27824, n26656, \imm[0] , cycle, n10486, \alu_b_in[3] , 
            n31949, n31946, n4325, \additional_mem_ops_2__N_749[0] , 
            n27018, n31741, n32040, is_load, n844, n26290, clk_c_enable_527, 
            n32046, interrupt_core, n31876, n5014, n1766, \instr_write_offset_3__N_934[1] , 
            \debug_branch_N_450[1] , n1767, \instr_write_offset_3__N_934[0] , 
            n15, n31743, n1768, pc_2__N_932, n29665, n31311, debug_rd, 
            instr_fetch_running, was_early_branch, n31745, n31957, \ui_in_sync[1] , 
            debug_rd_3__N_1575, n31915, n31892, load_done_N_1741, \data_rs2[0] , 
            \data_rs2[2] , n84, \data_rs2[1] , \next_fsm_state_3__N_3015[3] , 
            rd, fsm_state, debug_instr_valid, is_lui, is_jal, n31948, 
            n31966, clk_c_enable_169, is_branch, is_jalr, is_auipc, 
            is_system, n33486, n33484, clk_c_enable_165, \imm[5] , 
            \imm[3] , n32015, mem_op, n31987, n26175, n31955, accum, 
            d_3__N_1868, n31929, timer_interrupt, clk_c_enable_181, 
            \mul_out[1] , clk_c_enable_184, n32185, \timer_data[0] , 
            is_timer_addr, \mul_out[2] , data_out_3__N_1385, n29318, 
            n31319, \timer_data[2] , \mul_out[3] , n31999, \debug_branch_N_450[3] , 
            load_top_bit, n5677, \imm[7] , n9033, \imm[11] , is_alu_imm, 
            is_alu_reg, debug_rd_3__N_413, \cycle_count_wide[3] , n5626, 
            n32049, \imm[9] , \imm[8] , \addr_out[26] , \imm[4] , 
            \addr_out[25] , \addr_out[24] , \addr_out[27] , mstatus_mie_N_1709, 
            mstatus_mie_N_1707, n26997, n28222, n26995, n109, n26996, 
            n31963, n31932, next_bit, n28800, n31389, \data_out_slice[0] , 
            is_store, n9710, n29739, n13, n29194, n29137, n29330, 
            \debug_branch_N_450[0] , n32044, n32039, n29190, n29149, 
            \debug_branch_N_446[28] , n238, n29240, n31768, data_ready_sync, 
            data_ready_core, \next_pc_for_core[20] , \next_pc_for_core[16] , 
            n225, \pc[23] , \pc[19] , n30741, \pc[21] , \pc[17] , 
            n30802, \next_pc_for_core[22] , \next_pc_for_core[18] , n227, 
            \pc[20] , \pc[16] , n225_adj_1, \pc[22] , \pc[18] , n30746, 
            \next_pc_for_core[21] , \next_pc_for_core[17] , n226, \debug_branch_N_442[31] , 
            alu_a_in_3__N_1552, \debug_branch_N_442[30] , \debug_rd_3__N_405[30] , 
            alu_b_in_3__N_1504, \debug_rd_3__N_405[29] , n157, \debug_branch_N_442[28] , 
            n29220, \debug_rd_3__N_405[28] , \debug_branch_N_442[29] , 
            n29147, \debug_branch_N_446[30] , n29333, n29135, \debug_branch_N_446[29] , 
            n15604, \data_out_slice[2] , \data_out_slice[1] , n31972, 
            n31914, \timer_data[1] , \mem_data_from_read[17] , \mem_data_from_read[21] , 
            n31310, \addr_offset[2] , n701, n29012, n29162, \debug_rd_3__N_405[31] , 
            rst_reg_n, cy, time_pulse_r, n10573, n31889, n9538, 
            \mtime_out[0] , n31913, n31872, \addr_out[23] , \addr_out[0] , 
            \addr_out[1] , n31898, \addr_out[22] , \addr_out[21] , \addr_out[20] , 
            \addr_out[19] , \addr_out[18] , \addr_out[17] , \addr_out[16] , 
            \addr_out[15] , \addr_out[14] , \addr_out[13] , \addr_out[12] , 
            \addr_out[11] , \addr_out[10] , \addr_out[9] , \addr_out[8] , 
            \addr_out[7] , \addr_out[6] , \addr_out[5] , \addr_out[4] , 
            \addr_out[3] , n33493, instr_complete_N_1651, n5661, n28282, 
            \next_pc_offset[3] , n27604, n31888, n18086, \debug_branch_N_446[31] , 
            \csr_read_3__N_1443[0] , \csr_read_3__N_1447[2] , GND_net, 
            VCC_net, \next_accum[5] , \next_accum[6] , \next_accum[7] , 
            \next_accum[8] , \next_accum[9] , \next_accum[10] , \next_accum[11] , 
            \next_accum[12] , \next_accum[13] , \next_accum[14] , \next_accum[15] , 
            \next_accum[16] , \next_accum[17] , \next_accum[18] , \next_accum[19] , 
            \next_accum[4] , rs2, n12_adj_2, n11, n9, n8, rs1, 
            return_addr, \registers[5][7] , \registers[6][7] , \registers[7][7] , 
            n27480, n31747, no_write_in_progress, n28150, n27762, 
            n28182, n29747, n4, \reg_access[3][2] , n30165, n30166, 
            n30169, n31748, n30167, n30168, n31870) /* synthesis syn_module_defined=1 */ ;
    input clk_c;
    input n31841;
    input n31980;
    input clk_c_enable_234;
    input [4:2]counter_hi;
    input [3:0]n92;
    input n18324;
    output instr_complete_N_1647;
    input clk_c_enable_449;
    input \ui_in_sync[0] ;
    output mstatus_mte;
    input \imm[10] ;
    output n31744;
    output n31738;
    input n27838;
    output n31742;
    output n26648;
    input \imm[1] ;
    input n27934;
    output n26764;
    input n27874;
    output n26794;
    output [3:0]data_rs1;
    input n27810;
    output n2804;
    input n27886;
    output n26788;
    input n28020;
    output n2498;
    input n27960;
    output n3402;
    input n28068;
    output n26807;
    input n28080;
    output n26889;
    input n27672;
    input n31758;
    output n31733;
    input n27862;
    output n2592;
    input n9894;
    input n27728;
    output n27734;
    input \next_pc_for_core[7] ;
    input \next_pc_for_core[3] ;
    input n27910;
    output n26776;
    input \next_pc_for_core[23] ;
    input \next_pc_for_core[19] ;
    input n28116;
    output n26871;
    input n27946;
    output n31735;
    input \next_pc_for_core[15] ;
    input \next_pc_for_core[11] ;
    input n27922;
    output n26770;
    input \alu_op[0] ;
    input \alu_op[3] ;
    input \alu_op[1] ;
    input \alu_op_in[2] ;
    input n29006;
    output n28881;
    input n27738;
    output n27744;
    input n27898;
    output n26782;
    input n30947;
    input n31853;
    output n30949;
    input n27790;
    input n12;
    output n27796;
    input n28128;
    output n26827;
    input n28140;
    output n26905;
    input n28054;
    output n26814;
    input n31894;
    input n31875;
    output n1160;
    output load_done;
    output clk_c_enable_249;
    input n8289;
    input \imm[2] ;
    input \imm[6] ;
    input clk_c_enable_233;
    input n27576;
    input n31720;
    output n26800;
    input n31838;
    input is_jalr_N_1370;
    output n27724;
    input n28040;
    output n26821;
    input stall_core;
    output clk_c_enable_36;
    input n28204;
    output n26993;
    output is_double_fault_r;
    output n31893;
    output n31878;
    input n28092;
    output n26883;
    input n28104;
    output n26877;
    input n27824;
    output n26656;
    input \imm[0] ;
    output [1:0]cycle;
    output n10486;
    input \alu_b_in[3] ;
    output n31949;
    output n31946;
    input n4325;
    output \additional_mem_ops_2__N_749[0] ;
    input n27018;
    output n31741;
    input n32040;
    input is_load;
    output n844;
    input n26290;
    output clk_c_enable_527;
    input n32046;
    input interrupt_core;
    output n31876;
    input [1:0]n5014;
    input n1766;
    output \instr_write_offset_3__N_934[1] ;
    input \debug_branch_N_450[1] ;
    input n1767;
    output \instr_write_offset_3__N_934[0] ;
    input n15;
    output n31743;
    input [1:0]n1768;
    output [1:0]pc_2__N_932;
    input n29665;
    input n31311;
    output [3:0]debug_rd;
    input instr_fetch_running;
    input was_early_branch;
    output n31745;
    output n31957;
    input \ui_in_sync[1] ;
    input debug_rd_3__N_1575;
    input n31915;
    input n31892;
    output load_done_N_1741;
    output \data_rs2[0] ;
    output \data_rs2[2] ;
    input n84;
    output \data_rs2[1] ;
    input \next_fsm_state_3__N_3015[3] ;
    input [3:0]rd;
    input [3:0]fsm_state;
    input debug_instr_valid;
    input is_lui;
    input is_jal;
    input n31948;
    input n31966;
    output clk_c_enable_169;
    input is_branch;
    input is_jalr;
    input is_auipc;
    input is_system;
    input n33486;
    input n33484;
    output clk_c_enable_165;
    input \imm[5] ;
    input \imm[3] ;
    input n32015;
    input [2:0]mem_op;
    input n31987;
    output n26175;
    output n31955;
    output [15:0]accum;
    output [19:0]d_3__N_1868;
    output n31929;
    input timer_interrupt;
    output clk_c_enable_181;
    input \mul_out[1] ;
    output clk_c_enable_184;
    input n32185;
    input \timer_data[0] ;
    input is_timer_addr;
    input \mul_out[2] ;
    output data_out_3__N_1385;
    input n29318;
    input n31319;
    input \timer_data[2] ;
    input \mul_out[3] ;
    output n31999;
    input \debug_branch_N_450[3] ;
    output load_top_bit;
    output [3:0]n5677;
    input \imm[7] ;
    output n9033;
    input \imm[11] ;
    input is_alu_imm;
    input is_alu_reg;
    input debug_rd_3__N_413;
    output \cycle_count_wide[3] ;
    output n5626;
    input n32049;
    input \imm[9] ;
    input \imm[8] ;
    output \addr_out[26] ;
    input \imm[4] ;
    output \addr_out[25] ;
    output \addr_out[24] ;
    output \addr_out[27] ;
    output mstatus_mie_N_1709;
    input mstatus_mie_N_1707;
    output n26997;
    input n28222;
    output n26995;
    input n109;
    output n26996;
    output n31963;
    output n31932;
    input next_bit;
    output n28800;
    input n31389;
    output \data_out_slice[0] ;
    input is_store;
    output n9710;
    input n29739;
    input n13;
    output n29194;
    input n29137;
    input n29330;
    input \debug_branch_N_450[0] ;
    output n32044;
    output n32039;
    input n29190;
    input n29149;
    input \debug_branch_N_446[28] ;
    input n238;
    input n29240;
    input n31768;
    input data_ready_sync;
    output data_ready_core;
    input \next_pc_for_core[20] ;
    input \next_pc_for_core[16] ;
    output n225;
    input \pc[23] ;
    input \pc[19] ;
    output n30741;
    input \pc[21] ;
    input \pc[17] ;
    output n30802;
    input \next_pc_for_core[22] ;
    input \next_pc_for_core[18] ;
    output n227;
    input \pc[20] ;
    input \pc[16] ;
    output n225_adj_1;
    input \pc[22] ;
    input \pc[18] ;
    output n30746;
    input \next_pc_for_core[21] ;
    input \next_pc_for_core[17] ;
    output n226;
    input \debug_branch_N_442[31] ;
    output alu_a_in_3__N_1552;
    input \debug_branch_N_442[30] ;
    input \debug_rd_3__N_405[30] ;
    output alu_b_in_3__N_1504;
    input \debug_rd_3__N_405[29] ;
    input n157;
    input \debug_branch_N_442[28] ;
    input n29220;
    input \debug_rd_3__N_405[28] ;
    input \debug_branch_N_442[29] ;
    input n29147;
    input \debug_branch_N_446[30] ;
    input n29333;
    input n29135;
    input \debug_branch_N_446[29] ;
    output n15604;
    output \data_out_slice[2] ;
    output \data_out_slice[1] ;
    input n31972;
    input n31914;
    input \timer_data[1] ;
    input \mem_data_from_read[17] ;
    input \mem_data_from_read[21] ;
    output n31310;
    input \addr_offset[2] ;
    output n701;
    input n29012;
    input n29162;
    input \debug_rd_3__N_405[31] ;
    input rst_reg_n;
    input cy;
    input time_pulse_r;
    input n10573;
    output n31889;
    output n9538;
    input \mtime_out[0] ;
    input n31913;
    output n31872;
    output \addr_out[23] ;
    output \addr_out[0] ;
    output \addr_out[1] ;
    output n31898;
    output \addr_out[22] ;
    output \addr_out[21] ;
    output \addr_out[20] ;
    output \addr_out[19] ;
    output \addr_out[18] ;
    output \addr_out[17] ;
    output \addr_out[16] ;
    output \addr_out[15] ;
    output \addr_out[14] ;
    output \addr_out[13] ;
    output \addr_out[12] ;
    output \addr_out[11] ;
    output \addr_out[10] ;
    output \addr_out[9] ;
    output \addr_out[8] ;
    output \addr_out[7] ;
    output \addr_out[6] ;
    output \addr_out[5] ;
    output \addr_out[4] ;
    output \addr_out[3] ;
    output n33493;
    input instr_complete_N_1651;
    input n5661;
    output n28282;
    input \next_pc_offset[3] ;
    output n27604;
    input n31888;
    output n18086;
    input \debug_branch_N_446[31] ;
    input \csr_read_3__N_1443[0] ;
    output \csr_read_3__N_1447[2] ;
    input GND_net;
    input VCC_net;
    input \next_accum[5] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[4] ;
    input [3:0]rs2;
    output n12_adj_2;
    output n11;
    output n9;
    output n8;
    input [3:0]rs1;
    output [23:1]return_addr;
    output \registers[5][7] ;
    output \registers[6][7] ;
    output \registers[7][7] ;
    output n27480;
    output n31747;
    input no_write_in_progress;
    input n28150;
    output n27762;
    output n28182;
    output n29747;
    input n4;
    output \reg_access[3][2] ;
    output n30165;
    output n30166;
    output n30169;
    output n31748;
    output n30167;
    output n30168;
    output n31870;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [16:0]mie;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(323[16:19])
    
    wire clk_c_enable_274, n30581;
    wire [5:0]mcause;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(325[15:21])
    
    wire clk_c_enable_251;
    wire [5:0]n611;
    wire [17:16]mip_reg;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(321[17:24])
    wire [1:0]n979;
    wire [2:0]time_hi;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(292[15:22])
    wire [2:0]n1;
    
    wire n31988, cy_c, instr_retired, n31890;
    wire [5:0]shift_amt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[16:25])
    
    wire clk_c_enable_80;
    wire [4:0]shift_amt_adj_3116;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(124[15:24])
    
    wire clk_c_enable_77, cmp, cmp_out;
    wire [31:0]tmp_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(88[16:24])
    
    wire clk_c_enable_544;
    wire [23:0]mepc;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(68[16:20])
    
    wire clk_c_enable_543;
    wire [1:0]last_interrupt_req;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(417[15:33])
    
    wire cy_adj_3108, cy_out, clk_c_enable_137, mstatus_mte_N_1703, 
        n32095, n31588, n31589;
    wire [6:0]cycle_count_wide;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(279[16:32])
    
    wire cy_adj_3109, n31912, n31959, n31924;
    wire [4:0]increment_result_3__N_1911;
    
    wire n32094, n32093, n32098, n32097;
    wire [3:0]tmp_data_in_3__N_1582;
    
    wire n5737;
    wire [3:0]tmp_data_in_3__N_1514;
    
    wire n32329, n32326, n32327, n30969, n30968, n4874;
    wire [3:0]csr_read_3__N_1447;
    
    wire n26019, n28972, n30989, n30988;
    wire [3:0]time_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(299[16:26])
    
    wire n29171;
    wire [3:0]n5633;
    
    wire n26121;
    wire [3:0]n5665;
    
    wire n32004, n31981, instr_complete_N_1652, n32008, n30868, n30870;
    wire [3:0]alu_b_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[16:24])
    wire [3:0]alu_a_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[16:24])
    wire [3:0]n4913;
    
    wire n10727, n26148, n28518, n7754, n26149, n24774, n28520;
    wire [3:0]csr_read_3__N_1455;
    
    wire n31353, n31351, n31956, debug_reg_wen, n31917, n31943, 
        n29163;
    wire [2:0]n498;
    
    wire interrupt_pending_N_1671, n27534, n25168, n32024, n27089, 
        n32045, n32023, n27061, n27308, n6096, n31938, mstatus_mpie, 
        clk_c_enable_250, n6337, clk_c_enable_252, n25282, clk_c_enable_258, 
        n25292, n926, n927, n928, clk_c_enable_264, n25290, n893, 
        n894, n895, clk_c_enable_269, n25288, n860, n861, n31896, 
        n31926, n862, n25284, n793, n26597, n794, n31313, n29329;
    wire [3:0]debug_rd_3__N_1571;
    
    wire n652;
    wire [3:0]n653;
    
    wire n32005;
    wire [3:0]n191;
    wire [3:0]shift_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(132[16:25])
    
    wire n31746, n29550;
    wire [3:0]n196;
    wire [3:0]debug_rd_3__N_1559;
    wire [3:0]debug_rd_3__N_1563;
    wire [3:0]debug_rd_3__N_1396;
    
    wire n31312;
    wire [3:0]debug_rd_3__N_1392;
    wire [3:0]csr_read_3__N_1459;
    
    wire clk_c_enable_348, n31, n10548, n17438;
    wire [3:0]data_rs1_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(83[16:24])
    wire [3:0]debug_rd_3__N_1567;
    
    wire n30944, n28620, n31842, n14, n21, n28946, n27176, n18, 
        n30945;
    wire [1:0]n948;
    wire [1:0]n809;
    wire [1:0]n822;
    
    wire n30580;
    wire [3:0]alu_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(110[16:23])
    
    wire n30704, n30701, n31973;
    wire [3:0]tmp_data_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(242[15:26])
    wire [59:0]debug_branch_N_840;
    
    wire n30702, n30703, n28210, n32025, n28318, n10873, n18719, 
        n30987, n31947, n28558, n31854, clk_c_enable_536, n31983, 
        n27528, n26486, n28374, load_top_bit_next_N_1731, n27288, 
        n31945, n18685, clk_c_enable_545, n31172, n31173, instr_complete_N_1656, 
        instr_complete_N_1654, n29158, n5670, n46, debug_rd_3__N_1401, 
        n11557, n30667, n30665, n30668, n30695, n31826, n31827, 
        n31825, n29243, n31856, n31960, n31979;
    wire [3:0]instrret_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(301[16:30])
    wire [3:0]n5624;
    
    wire n31874, n32011, n29539, n29008, n40, n28508, n27180, 
        n8_adj_3110, n32014, n11559;
    wire [3:0]n658;
    
    wire n20, mstatus_mie, n29155, n31174, n31690;
    wire [3:0]n5671;
    
    wire n30666, n31689, instr_complete_N_1650, instr_complete_N_1649, 
        instr_complete_N_1648;
    wire [3:0]n234;
    
    wire n30669, n29351, n30696, n31171, n18076, n30699, n10513;
    wire [2:0]n5054;
    
    wire n31909, n31586, n31587, n31891, n33494;
    wire [3:0]mul_out_3__N_1510;
    
    wire n31843, n21568, n8_adj_3112, n29164, n29153, n29154, n29156, 
        n29157, n31352, n29010, n15837, n31873;
    wire [4:0]increment_result_3__N_1925;
    
    wire n27558, n31787, n28436;
    wire [3:0]csr_read_3__N_1439;
    
    wire n28664, n31688, n18009, n32330, n32328;
    wire [3:0]csr_read_3__N_1451;
    
    FD1P3IX mie__i0 (.D(n30581), .SP(clk_c_enable_274), .CD(n31841), .CK(clk_c), 
            .Q(mie[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i0.GSR = "DISABLED";
    FD1P3IX mcause__i0 (.D(n611[0]), .SP(clk_c_enable_251), .CD(n31980), 
            .CK(clk_c), .Q(mcause[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i0.GSR = "DISABLED";
    FD1P3IX mip_reg__i16 (.D(n979[0]), .SP(clk_c_enable_234), .CD(n31841), 
            .CK(clk_c), .Q(mip_reg[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mip_reg__i16.GSR = "DISABLED";
    FD1S3IX time_hi__i0 (.D(n1[0]), .CK(clk_c), .CD(n31980), .Q(time_hi[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i0.GSR = "DISABLED";
    LUT4 cy_I_0_3_lut_rep_685_3_lut_4_lut (.A(n31988), .B(counter_hi[2]), 
         .C(cy_c), .D(instr_retired), .Z(n31890)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam cy_I_0_3_lut_rep_685_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX shift_amt__i1 (.D(n92[0]), .SP(clk_c_enable_80), .CK(clk_c), 
            .Q(shift_amt[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i1.GSR = "DISABLED";
    FD1P3AX shift_amt__i5 (.D(n92[0]), .SP(clk_c_enable_77), .CK(clk_c), 
            .Q(shift_amt_adj_3116[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i5.GSR = "DISABLED";
    FD1P3AX shift_amt__i4 (.D(n92[3]), .SP(clk_c_enable_80), .CK(clk_c), 
            .Q(shift_amt_adj_3116[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i4.GSR = "DISABLED";
    FD1P3AX shift_amt__i3 (.D(n92[2]), .SP(clk_c_enable_80), .CK(clk_c), 
            .Q(shift_amt_adj_3116[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i3.GSR = "DISABLED";
    FD1P3AX shift_amt__i2 (.D(n92[1]), .SP(clk_c_enable_80), .CK(clk_c), 
            .Q(shift_amt[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(125[12] 130[8])
    defparam shift_amt__i2.GSR = "DISABLED";
    FD1S3IX instr_retired_518 (.D(instr_complete_N_1647), .CK(clk_c), .CD(n18324), 
            .Q(instr_retired)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(303[12] 305[8])
    defparam instr_retired_518.GSR = "DISABLED";
    FD1S3AX cmp_511 (.D(cmp_out), .CK(clk_c), .Q(cmp)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(117[12] 120[8])
    defparam cmp_511.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i0 (.D(tmp_data[4]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i0.GSR = "DISABLED";
    FD1P3AX mepc_i0_i0 (.D(mepc[4]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i0.GSR = "DISABLED";
    FD1P3AX last_interrupt_req_i0_i0 (.D(\ui_in_sync[0] ), .SP(clk_c_enable_449), 
            .CK(clk_c), .Q(last_interrupt_req[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam last_interrupt_req_i0_i0.GSR = "DISABLED";
    FD1S3AX cy_510 (.D(cy_out), .CK(clk_c), .Q(cy_adj_3108)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(117[12] 120[8])
    defparam cy_510.GSR = "DISABLED";
    FD1P3BX mstatus_mte_523 (.D(mstatus_mte_N_1703), .SP(clk_c_enable_137), 
            .CK(clk_c), .PD(n31980), .Q(mstatus_mte)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(384[18] 390[12])
    defparam mstatus_mte_523.GSR = "DISABLED";
    LUT4 n5655_bdd_3_lut (.A(n32095), .B(n31588), .C(\imm[10] ), .Z(n31589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n5655_bdd_3_lut.init = 16'hcaca;
    LUT4 i4755_2_lut_rep_707_3_lut_4_lut (.A(n31988), .B(counter_hi[2]), 
         .C(cycle_count_wide[0]), .D(cy_adj_3109), .Z(n31912)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i4755_2_lut_rep_707_3_lut_4_lut.init = 16'hf010;
    LUT4 cy_I_0_3_lut_rep_719_4_lut (.A(n31988), .B(counter_hi[2]), .C(n31959), 
         .D(cy_adj_3108), .Z(n31924)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam cy_I_0_3_lut_rep_719_4_lut.init = 16'hfe10;
    LUT4 i4753_2_lut_3_lut_4_lut (.A(n31988), .B(counter_hi[2]), .C(cycle_count_wide[0]), 
         .D(cy_adj_3109), .Z(increment_result_3__N_1911[0])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i4753_2_lut_3_lut_4_lut.init = 16'h0fe1;
    LUT4 i1_4_lut_4_lut_4_lut (.A(n31744), .B(n31738), .C(n27838), .D(n31742), 
         .Z(n26648)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i15539_4_lut_then_4_lut (.A(\imm[1] ), .B(mcause[4]), .C(counter_hi[4]), 
         .D(counter_hi[3]), .Z(n32094)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i15539_4_lut_then_4_lut.init = 16'h0008;
    LUT4 i15539_4_lut_else_4_lut (.A(mcause[0]), .B(\imm[1] ), .C(counter_hi[4]), 
         .D(counter_hi[3]), .Z(n32093)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i15539_4_lut_else_4_lut.init = 16'h0008;
    LUT4 i1_4_lut_4_lut_4_lut_adj_279 (.A(n31744), .B(n31738), .C(n27934), 
         .D(n31742), .Z(n26764)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_279.init = 16'h0040;
    LUT4 n30953_bdd_4_lut_then_4_lut (.A(mie[14]), .B(mie[6]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n32098)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !((C+!(D))+!B)) */ ;
    defparam n30953_bdd_4_lut_then_4_lut.init = 16'hac00;
    LUT4 n30953_bdd_4_lut_else_4_lut (.A(mie[10]), .B(mie[2]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n32097)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !((C+!(D))+!B)) */ ;
    defparam n30953_bdd_4_lut_else_4_lut.init = 16'hac00;
    LUT4 i1_4_lut_4_lut_4_lut_adj_280 (.A(n31744), .B(n31738), .C(n27874), 
         .D(n31742), .Z(n26794)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_280.init = 16'h0040;
    LUT4 tmp_data_in_3__I_124_i1_3_lut (.A(tmp_data_in_3__N_1582[0]), .B(data_rs1[0]), 
         .C(n5737), .Z(tmp_data_in_3__N_1514[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_124_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_4_lut_adj_281 (.A(n31744), .B(n31738), .C(n27810), 
         .D(n31742), .Z(n2804)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_281.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_282 (.A(n31744), .B(n31738), .C(n27886), 
         .D(n31742), .Z(n26788)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_282.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_283 (.A(n31744), .B(n31738), .C(n28020), 
         .D(n31742), .Z(n2498)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_283.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_284 (.A(n31744), .B(n31738), .C(n27960), 
         .D(n31742), .Z(n3402)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_284.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_285 (.A(n31744), .B(n31738), .C(n28068), 
         .D(n31742), .Z(n26807)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_285.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_286 (.A(n31744), .B(n31738), .C(n28080), 
         .D(n31742), .Z(n26889)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_286.init = 16'h0040;
    LUT4 i3_rep_528_4_lut (.A(n31744), .B(n27672), .C(n31738), .D(n31758), 
         .Z(n31733)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i3_rep_528_4_lut.init = 16'h4000;
    LUT4 i3129_4_lut_4_lut_4_lut (.A(n31744), .B(n31738), .C(n27862), 
         .D(n31742), .Z(n2592)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i3129_4_lut_4_lut_4_lut.init = 16'hffbf;
    LUT4 i1_4_lut_4_lut_4_lut_adj_287 (.A(n31744), .B(n9894), .C(n27728), 
         .D(n31742), .Z(n27734)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_287.init = 16'h0010;
    LUT4 debug_branch_N_446_31__bdd_3_lut (.A(\next_pc_for_core[7] ), .B(\next_pc_for_core[3] ), 
         .C(counter_hi[2]), .Z(n32329)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam debug_branch_N_446_31__bdd_3_lut.init = 16'hacac;
    LUT4 i1_4_lut_4_lut_4_lut_adj_288 (.A(n31744), .B(n31738), .C(n27910), 
         .D(n31742), .Z(n26776)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_288.init = 16'h0040;
    LUT4 next_pc_for_core_23__bdd_4_lut (.A(\next_pc_for_core[23] ), .B(\next_pc_for_core[19] ), 
         .C(counter_hi[3]), .D(counter_hi[2]), .Z(n32326)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam next_pc_for_core_23__bdd_4_lut.init = 16'h0a0c;
    LUT4 i1_4_lut_4_lut_4_lut_adj_289 (.A(n31744), .B(n31738), .C(n28116), 
         .D(n31742), .Z(n26871)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_289.init = 16'h0040;
    LUT4 i1_4_lut_rep_530_4_lut_4_lut (.A(n31744), .B(n31738), .C(n27946), 
         .D(n31742), .Z(n31735)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_rep_530_4_lut_4_lut.init = 16'h0040;
    LUT4 next_pc_for_core_23__bdd_3_lut (.A(\next_pc_for_core[15] ), .B(\next_pc_for_core[11] ), 
         .C(counter_hi[2]), .Z(n32327)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam next_pc_for_core_23__bdd_3_lut.init = 16'hacac;
    LUT4 n30969_bdd_4_lut (.A(n30969), .B(n30968), .C(counter_hi[2]), 
         .D(n4874), .Z(csr_read_3__N_1447[1])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n30969_bdd_4_lut.init = 16'hca00;
    LUT4 i1_4_lut_4_lut_4_lut_adj_290 (.A(n31744), .B(n31738), .C(n27922), 
         .D(n31742), .Z(n26770)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_290.init = 16'h0040;
    LUT4 i11_4_lut (.A(\alu_op[0] ), .B(\alu_op[3] ), .C(\alu_op[1] ), 
         .D(\alu_op_in[2] ), .Z(n5737)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i11_4_lut.init = 16'hca0a;
    LUT4 i26324_4_lut_4_lut_4_lut (.A(n31744), .B(n31738), .C(n29006), 
         .D(n31742), .Z(n28881)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i26324_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_291 (.A(n31744), .B(n9894), .C(n27738), 
         .D(n31742), .Z(n27744)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_291.init = 16'h0010;
    LUT4 i1_4_lut_4_lut_4_lut_adj_292 (.A(n31744), .B(n31738), .C(n27898), 
         .D(n31742), .Z(n26782)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_292.init = 16'h0040;
    LUT4 instr_12__bdd_3_lut_28472_4_lut_4_lut (.A(n31744), .B(n31738), 
         .C(n30947), .D(n31853), .Z(n30949)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam instr_12__bdd_3_lut_28472_4_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_4_lut (.A(n31744), .B(n27790), .C(n12), .D(n9894), 
         .Z(n27796)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_293 (.A(n31744), .B(n31738), .C(n28128), 
         .D(n31742), .Z(n26827)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_293.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_294 (.A(n31744), .B(n31738), .C(n28140), 
         .D(n31742), .Z(n26905)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_294.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_295 (.A(n31744), .B(n31738), .C(n28054), 
         .D(n31742), .Z(n26814)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_295.init = 16'h0040;
    LUT4 i27901_4_lut (.A(n26019), .B(n31894), .C(n28972), .D(n31875), 
         .Z(n1160)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;
    defparam i27901_4_lut.init = 16'h5040;
    FD1P3AX load_done_515 (.D(n8289), .SP(clk_c_enable_249), .CK(clk_c), 
            .Q(load_done)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(232[12] 235[8])
    defparam load_done_515.GSR = "DISABLED";
    LUT4 i26414_2_lut (.A(\imm[2] ), .B(\imm[6] ), .Z(n28972)) /* synthesis lut_function=(A (B)) */ ;
    defparam i26414_2_lut.init = 16'h8888;
    LUT4 i5218_2_lut (.A(time_hi[0]), .B(clk_c_enable_233), .Z(n1[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam i5218_2_lut.init = 16'h6666;
    LUT4 n30989_bdd_4_lut (.A(n30989), .B(n30988), .C(counter_hi[2]), 
         .D(n4874), .Z(csr_read_3__N_1447[3])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n30989_bdd_4_lut.init = 16'hca00;
    LUT4 i1_4_lut_4_lut_adj_296 (.A(n31744), .B(n27576), .C(n31738), .D(n31720), 
         .Z(n26800)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_296.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_adj_297 (.A(n31744), .B(n31838), .C(n9894), .D(is_jalr_N_1370), 
         .Z(n27724)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_adj_297.init = 16'h0100;
    LUT4 i1_4_lut_4_lut_4_lut_adj_298 (.A(n31744), .B(n31738), .C(n28040), 
         .D(n31742), .Z(n26821)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_298.init = 16'h0040;
    LUT4 i1_4_lut (.A(stall_core), .B(instr_complete_N_1647), .C(clk_c_enable_36), 
         .D(n28204), .Z(n26993)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut.init = 16'h8000;
    LUT4 i15342_2_lut_4_lut (.A(mstatus_mte), .B(is_double_fault_r), .C(n31893), 
         .D(n31878), .Z(mstatus_mte_N_1703)) /* synthesis lut_function=(A (B+!(D))+!A (B+(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(365[28:90])
    defparam i15342_2_lut_4_lut.init = 16'hdcff;
    LUT4 i1_4_lut_4_lut_4_lut_adj_299 (.A(n31744), .B(n31738), .C(n28092), 
         .D(n31742), .Z(n26883)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_299.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_300 (.A(n31744), .B(n31738), .C(n28104), 
         .D(n31742), .Z(n26877)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_300.init = 16'h0040;
    LUT4 i1_4_lut_4_lut_4_lut_adj_301 (.A(n31744), .B(n31738), .C(n27824), 
         .D(n31742), .Z(n26656)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_adj_301.init = 16'h0040;
    LUT4 i26554_3_lut (.A(cycle_count_wide[1]), .B(time_count[1]), .C(\imm[0] ), 
         .Z(n29171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26554_3_lut.init = 16'hcaca;
    LUT4 mux_3522_i2_4_lut (.A(n5633[1]), .B(mepc[1]), .C(\imm[0] ), .D(n26121), 
         .Z(n5665[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3522_i2_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_302 (.A(cycle[0]), .B(n10486), .C(n32004), .D(n31981), 
         .Z(instr_complete_N_1652)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;
    defparam i1_4_lut_adj_302.init = 16'h6aaa;
    LUT4 n30870_bdd_3_lut_4_lut (.A(\alu_op[0] ), .B(n32008), .C(n30868), 
         .D(n30870), .Z(cmp_out)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam n30870_bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_3036_i1_3_lut_4_lut (.A(\alu_op[0] ), .B(n32008), .C(alu_b_in[0]), 
         .D(alu_a_in[0]), .Z(n4913[0])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam mux_3036_i1_3_lut_4_lut.init = 16'hfdd0;
    LUT4 mux_3036_i4_3_lut_4_lut (.A(\alu_op[0] ), .B(n32008), .C(\alu_b_in[3] ), 
         .D(alu_a_in[3]), .Z(n4913[3])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam mux_3036_i4_3_lut_4_lut.init = 16'hfdd0;
    LUT4 mux_3036_i2_3_lut_4_lut (.A(\alu_op[0] ), .B(n32008), .C(alu_b_in[1]), 
         .D(alu_a_in[1]), .Z(n4913[1])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam mux_3036_i2_3_lut_4_lut.init = 16'hfdd0;
    LUT4 mux_3036_i3_3_lut_4_lut (.A(\alu_op[0] ), .B(n32008), .C(alu_b_in[2]), 
         .D(alu_a_in[2]), .Z(n4913[2])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (C+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(106[28:55])
    defparam mux_3036_i3_3_lut_4_lut.init = 16'hfdd0;
    LUT4 i1_4_lut_adj_303 (.A(n10727), .B(n26148), .C(n28518), .D(n7754), 
         .Z(n26149)) /* synthesis lut_function=(A (B)+!A !((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_303.init = 16'h888c;
    LUT4 i1_3_lut_4_lut (.A(instr_complete_N_1647), .B(clk_c_enable_36), 
         .C(cycle[1]), .D(cycle[0]), .Z(n24774)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_4_lut.init = 16'h0770;
    LUT4 csr_read_3__I_128_i4_4_lut (.A(mcause[3]), .B(n28520), .C(n31949), 
         .D(n31946), .Z(csr_read_3__N_1455[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(490[33] 493[57])
    defparam csr_read_3__I_128_i4_4_lut.init = 16'hca0a;
    PFUMX i28409 (.BLUT(n31353), .ALUT(n31351), .C0(n31956), .Z(debug_reg_wen));
    LUT4 i1_2_lut_4_lut (.A(stall_core), .B(instr_complete_N_1647), .C(n31917), 
         .D(n4325), .Z(\additional_mem_ops_2__N_749[0] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_4_lut.init = 16'h7f80;
    LUT4 interrupt_core_I_32_2_lut_rep_536_4_lut (.A(stall_core), .B(instr_complete_N_1647), 
         .C(n31943), .D(n27018), .Z(n31741)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam interrupt_core_I_32_2_lut_rep_536_4_lut.init = 16'h80ff;
    LUT4 i26546_4_lut (.A(n32040), .B(mepc[2]), .C(\imm[6] ), .D(clk_c_enable_543), 
         .Z(n29163)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i26546_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_4_lut_adj_304 (.A(stall_core), .B(instr_complete_N_1647), 
         .C(n31943), .D(is_load), .Z(n844)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_4_lut_adj_304.init = 16'h80ff;
    LUT4 i1_2_lut_4_lut_adj_305 (.A(stall_core), .B(instr_complete_N_1647), 
         .C(n31943), .D(n26290), .Z(clk_c_enable_527)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_2_lut_4_lut_adj_305.init = 16'hff80;
    FD1P3IX time_hi__i2 (.D(n498[2]), .SP(clk_c_enable_233), .CD(n31980), 
            .CK(clk_c), .Q(time_hi[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i2.GSR = "DISABLED";
    FD1P3IX time_hi__i1 (.D(n498[1]), .SP(clk_c_enable_233), .CD(n31980), 
            .CK(clk_c), .Q(time_hi[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(293[12] 296[8])
    defparam time_hi__i1.GSR = "DISABLED";
    LUT4 i2_rep_539 (.A(n32046), .B(interrupt_pending_N_1671), .C(instr_complete_N_1647), 
         .D(n27534), .Z(n31744)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i2_rep_539.init = 16'h4000;
    FD1P3IX mip_reg__i17 (.D(n25168), .SP(clk_c_enable_234), .CD(n31841), 
            .CK(clk_c), .Q(mip_reg[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mip_reg__i17.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_306 (.A(n32024), .B(n27089), .C(n32045), .D(n32023), 
         .Z(n27061)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(331[17] 350[24])
    defparam i1_4_lut_adj_306.init = 16'hfdfc;
    FD1P3IX mcause__i5 (.D(interrupt_core), .SP(clk_c_enable_251), .CD(n31980), 
            .CK(clk_c), .Q(mcause[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i5.GSR = "DISABLED";
    FD1P3IX mcause__i4 (.D(n611[4]), .SP(clk_c_enable_251), .CD(n31980), 
            .CK(clk_c), .Q(mcause[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i4.GSR = "DISABLED";
    FD1P3IX mcause__i3 (.D(n27308), .SP(clk_c_enable_251), .CD(n31980), 
            .CK(clk_c), .Q(mcause[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i3.GSR = "DISABLED";
    FD1P3IX mcause__i2 (.D(n611[2]), .SP(clk_c_enable_251), .CD(n31980), 
            .CK(clk_c), .Q(mcause[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i2.GSR = "DISABLED";
    FD1P3IX is_double_fault_r_520 (.D(n31938), .SP(clk_c_enable_249), .CD(n6096), 
            .CK(clk_c), .Q(is_double_fault_r)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(361[12] 364[8])
    defparam is_double_fault_r_520.GSR = "DISABLED";
    FD1P3AX mstatus_mpie_525 (.D(n6337), .SP(clk_c_enable_250), .CK(clk_c), 
            .Q(mstatus_mpie)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam mstatus_mpie_525.GSR = "DISABLED";
    FD1P3IX mcause__i1 (.D(n611[1]), .SP(clk_c_enable_251), .CD(n31980), 
            .CK(clk_c), .Q(mcause[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(326[12] 357[8])
    defparam mcause__i1.GSR = "DISABLED";
    FD1P3IX mie__i16 (.D(n25282), .SP(clk_c_enable_252), .CD(n31841), 
            .CK(clk_c), .Q(mie[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i16.GSR = "DISABLED";
    FD1P3IX mie__i15 (.D(n25292), .SP(clk_c_enable_258), .CD(n31841), 
            .CK(clk_c), .Q(mie[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i15.GSR = "DISABLED";
    FD1P3IX mie__i14 (.D(n926), .SP(clk_c_enable_258), .CD(n31841), .CK(clk_c), 
            .Q(mie[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i14.GSR = "DISABLED";
    FD1P3IX mie__i13 (.D(n927), .SP(clk_c_enable_258), .CD(n31841), .CK(clk_c), 
            .Q(mie[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i13.GSR = "DISABLED";
    FD1P3IX mie__i12 (.D(n928), .SP(clk_c_enable_258), .CD(n31841), .CK(clk_c), 
            .Q(mie[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i12.GSR = "DISABLED";
    FD1P3IX mie__i11 (.D(n25290), .SP(clk_c_enable_264), .CD(n31841), 
            .CK(clk_c), .Q(mie[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i11.GSR = "DISABLED";
    FD1P3IX mie__i10 (.D(n893), .SP(clk_c_enable_264), .CD(n31841), .CK(clk_c), 
            .Q(mie[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i10.GSR = "DISABLED";
    FD1P3IX mie__i9 (.D(n894), .SP(clk_c_enable_264), .CD(n31841), .CK(clk_c), 
            .Q(mie[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i9.GSR = "DISABLED";
    FD1P3IX mie__i8 (.D(n895), .SP(clk_c_enable_264), .CD(n31841), .CK(clk_c), 
            .Q(mie[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i8.GSR = "DISABLED";
    FD1P3IX mie__i7 (.D(n25288), .SP(clk_c_enable_269), .CD(n31841), .CK(clk_c), 
            .Q(mie[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i7.GSR = "DISABLED";
    FD1P3IX mie__i6 (.D(n860), .SP(clk_c_enable_269), .CD(n31841), .CK(clk_c), 
            .Q(mie[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i6.GSR = "DISABLED";
    FD1P3IX mie__i5 (.D(n861), .SP(clk_c_enable_269), .CD(n31841), .CK(clk_c), 
            .Q(mie[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i5.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n31949), .B(n31896), .C(n31876), .D(n31926), 
         .Z(clk_c_enable_137)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(398[22:52])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff4;
    FD1P3IX mie__i4 (.D(n862), .SP(clk_c_enable_269), .CD(n31841), .CK(clk_c), 
            .Q(mie[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i4.GSR = "DISABLED";
    FD1P3IX mie__i3 (.D(n25284), .SP(clk_c_enable_274), .CD(n31841), .CK(clk_c), 
            .Q(mie[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i3.GSR = "DISABLED";
    FD1P3IX mie__i2 (.D(n793), .SP(clk_c_enable_274), .CD(n31841), .CK(clk_c), 
            .Q(mie[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i2.GSR = "DISABLED";
    LUT4 mux_351_i2_3_lut_4_lut (.A(clk_c_enable_36), .B(n26597), .C(n5014[1]), 
         .D(n1766), .Z(\instr_write_offset_3__N_934[1] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_351_i2_3_lut_4_lut.init = 16'hf780;
    FD1P3IX mie__i1 (.D(n794), .SP(clk_c_enable_274), .CD(n31841), .CK(clk_c), 
            .Q(mie[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam mie__i1.GSR = "DISABLED";
    PFUMX i28384 (.BLUT(n31313), .ALUT(\debug_branch_N_450[1] ), .C0(n29329), 
          .Z(debug_rd_3__N_1571[1]));
    LUT4 mux_351_i1_3_lut_4_lut (.A(clk_c_enable_36), .B(n26597), .C(n5014[0]), 
         .D(n1767), .Z(\instr_write_offset_3__N_934[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_351_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_251_i1_3_lut (.A(mepc[0]), .B(data_rs1[0]), .C(n652), .Z(n653[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i1_3_lut.init = 16'hcaca;
    LUT4 i27493_3_lut_rep_541_4_lut (.A(n32005), .B(n31981), .C(n191[3]), 
         .D(shift_out[3]), .Z(n31746)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i27493_3_lut_rep_541_4_lut.init = 16'hf2d0;
    LUT4 i27777_3_lut_4_lut (.A(n32005), .B(n31981), .C(n15), .D(n32008), 
         .Z(n29550)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i27777_3_lut_4_lut.init = 16'hffdf;
    LUT4 i27454_4_lut_4_lut (.A(n32008), .B(n15), .C(n196[0]), .D(n191[0]), 
         .Z(debug_rd_3__N_1559[0])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;
    defparam i27454_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i27496_3_lut_4_lut_4_lut (.A(n32008), .B(debug_rd_3__N_1563[3]), 
         .C(n15), .D(n31746), .Z(debug_rd_3__N_1396[3])) /* synthesis lut_function=(A (B)+!A (C (D))) */ ;
    defparam i27496_3_lut_4_lut_4_lut.init = 16'hd888;
    LUT4 interrupt_core_I_31_2_lut_rep_533_3_lut_4_lut (.A(clk_c_enable_36), 
         .B(n26597), .C(n31743), .D(n27018), .Z(n31738)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (C+!(D))) */ ;
    defparam interrupt_core_I_31_2_lut_rep_533_3_lut_4_lut.init = 16'hf8ff;
    LUT4 mux_352_i1_3_lut_4_lut (.A(clk_c_enable_36), .B(n26597), .C(n5014[0]), 
         .D(n1768[0]), .Z(pc_2__N_932[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_352_i1_3_lut_4_lut.init = 16'hf780;
    PFUMX i28382 (.BLUT(n29665), .ALUT(n31311), .C0(counter_hi[4]), .Z(n31312));
    LUT4 debug_rd_3__I_0_i1_3_lut (.A(debug_rd_3__N_1392[0]), .B(debug_rd_3__N_1396[0]), 
         .C(n31956), .Z(debug_rd[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(176[18] 194[12])
    defparam debug_rd_3__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_540_3_lut_4_lut (.A(clk_c_enable_36), .B(n26597), 
         .C(instr_fetch_running), .D(was_early_branch), .Z(n31745)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (C))) */ ;
    defparam i1_2_lut_rep_540_3_lut_4_lut.init = 16'h0f07;
    LUT4 mux_352_i2_3_lut_4_lut (.A(clk_c_enable_36), .B(n26597), .C(n5014[1]), 
         .D(n1768[1]), .Z(pc_2__N_932[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam mux_352_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 i15627_2_lut_3_lut_4_lut_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .D(mip_reg[16]), .Z(csr_read_3__N_1459[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i15627_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0400;
    FD1P3IX cycle__i1 (.D(n24774), .SP(clk_c_enable_348), .CD(n31980), 
            .CK(clk_c), .Q(cycle[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam cycle__i1.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_307 (.A(n32024), .B(n32023), .C(n31), .D(n10548), 
         .Z(n27089)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[48:59])
    defparam i1_3_lut_4_lut_adj_307.init = 16'h0100;
    LUT4 i1_4_lut_adj_308 (.A(mip_reg[17]), .B(n31957), .C(\ui_in_sync[1] ), 
         .D(last_interrupt_req[1]), .Z(n17438)) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(321[17:24])
    defparam i1_4_lut_adj_308.init = 16'h88c8;
    LUT4 mux_251_i4_3_lut (.A(mepc[3]), .B(data_rs1_c[3]), .C(n652), .Z(n653[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i4_3_lut.init = 16'hcaca;
    LUT4 debug_rd_3__I_0_i4_4_lut (.A(debug_rd_3__N_1567[3]), .B(debug_rd_3__N_1392[3]), 
         .C(n31956), .D(debug_rd_3__N_1575), .Z(debug_rd[3])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(176[18] 194[12])
    defparam debug_rd_3__I_0_i4_4_lut.init = 16'hccca;
    LUT4 counter_hi_2__bdd_4_lut_28148 (.A(mie[4]), .B(mie[12]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n30944)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam counter_hi_2__bdd_4_lut_28148.init = 16'hcac0;
    LUT4 i1_4_lut_adj_309 (.A(n1160), .B(n28620), .C(n31842), .D(n14), 
         .Z(n21)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_4_lut_adj_309.init = 16'ha8a0;
    LUT4 i1_4_lut_adj_310 (.A(n28946), .B(n27176), .C(n18), .D(\imm[1] ), 
         .Z(n652)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_310.init = 16'h0004;
    LUT4 i1_4_lut_adj_311 (.A(\imm[2] ), .B(n31915), .C(\imm[0] ), .D(\imm[6] ), 
         .Z(n27176)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_311.init = 16'h4000;
    LUT4 mux_251_i3_3_lut (.A(mepc[2]), .B(data_rs1_c[2]), .C(n652), .Z(n653[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i3_3_lut.init = 16'hcaca;
    LUT4 mux_251_i2_3_lut (.A(mepc[1]), .B(data_rs1_c[1]), .C(n652), .Z(n653[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(371[28] 372[75])
    defparam mux_251_i2_3_lut.init = 16'hcaca;
    LUT4 counter_hi_2__bdd_4_lut_28154 (.A(mie[8]), .B(mie[0]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n30945)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam counter_hi_2__bdd_4_lut_28154.init = 16'hacaa;
    LUT4 i15349_4_lut (.A(mip_reg[16]), .B(n31957), .C(\ui_in_sync[0] ), 
         .D(last_interrupt_req[0]), .Z(n948[0])) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(447[18] 459[12])
    defparam i15349_4_lut.init = 16'h88c8;
    LUT4 i15346_4_lut (.A(n809[0]), .B(n1160), .C(data_rs1[0]), .D(n31915), 
         .Z(n822[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(434[22] 438[16])
    defparam i15346_4_lut.init = 16'hc088;
    LUT4 mie_0__bdd_4_lut (.A(mie[0]), .B(data_rs1[0]), .C(n31894), .D(n31892), 
         .Z(n30580)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A (B (D))) */ ;
    defparam mie_0__bdd_4_lut.init = 16'hee2a;
    FD1P3AX tmp_data_i0_i1 (.D(tmp_data[5]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i1.GSR = "DISABLED";
    LUT4 mux_149_i1_3_lut_4_lut (.A(load_done_N_1741), .B(n32004), .C(alu_out[0]), 
         .D(\data_rs2[0] ), .Z(tmp_data_in_3__N_1582[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 counter_hi_2__bdd_4_lut_29130 (.A(mie[9]), .B(mie[1]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n30969)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam counter_hi_2__bdd_4_lut_29130.init = 16'hacaa;
    LUT4 mux_149_i3_3_lut_4_lut (.A(load_done_N_1741), .B(n32004), .C(alu_out[2]), 
         .D(\data_rs2[2] ), .Z(tmp_data_in_3__N_1582[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 i64_3_lut_4_lut (.A(load_done_N_1741), .B(n32004), .C(alu_out[3]), 
         .D(n84), .Z(tmp_data_in_3__N_1582[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam i64_3_lut_4_lut.init = 16'hfb40;
    LUT4 counter_hi_2__bdd_4_lut_28169 (.A(mie[5]), .B(mie[13]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n30968)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam counter_hi_2__bdd_4_lut_28169.init = 16'hcac0;
    LUT4 mux_149_i2_3_lut_4_lut (.A(load_done_N_1741), .B(n32004), .C(alu_out[1]), 
         .D(\data_rs2[1] ), .Z(tmp_data_in_3__N_1582[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(253[14] 256[36])
    defparam mux_149_i2_3_lut_4_lut.init = 16'hfb40;
    PFUMX i28029 (.BLUT(n30704), .ALUT(n30701), .C0(n31956), .Z(debug_rd[2]));
    LUT4 i1_4_lut_adj_312 (.A(n31), .B(n10548), .C(n31973), .D(n32045), 
         .Z(interrupt_pending_N_1671)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[48:59])
    defparam i1_4_lut_adj_312.init = 16'hfffe;
    FD1P3AX tmp_data_i0_i2 (.D(tmp_data[6]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i2.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i3 (.D(tmp_data[7]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i3.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i4 (.D(tmp_data[8]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i4.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i5 (.D(tmp_data[9]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i5.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i6 (.D(tmp_data[10]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i6.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i7 (.D(tmp_data[11]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i7.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i8 (.D(tmp_data[12]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i8.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i9 (.D(tmp_data[13]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i9.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i10 (.D(tmp_data[14]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i10.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i11 (.D(tmp_data[15]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i11.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i12 (.D(tmp_data[16]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i12.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i13 (.D(tmp_data[17]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i13.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i14 (.D(tmp_data[18]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i14.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i15 (.D(tmp_data[19]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i15.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i16 (.D(tmp_data[20]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i16.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i17 (.D(tmp_data[21]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i17.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i18 (.D(tmp_data[22]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i18.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i19 (.D(tmp_data[23]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i19.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i20 (.D(tmp_data[24]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i20.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i21 (.D(tmp_data[25]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i21.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i22 (.D(tmp_data[26]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i22.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i23 (.D(tmp_data[27]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i23.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i24 (.D(tmp_data[28]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i24.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i25 (.D(tmp_data[29]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i25.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i26 (.D(tmp_data[30]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i26.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i27 (.D(tmp_data[31]), .SP(clk_c_enable_544), .CK(clk_c), 
            .Q(tmp_data[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i27.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i30 (.D(tmp_data_in[2]), .SP(clk_c_enable_544), 
            .CK(clk_c), .Q(tmp_data[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i30.GSR = "DISABLED";
    FD1P3AX tmp_data_i0_i31 (.D(tmp_data_in[3]), .SP(clk_c_enable_544), 
            .CK(clk_c), .Q(tmp_data[31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i31.GSR = "DISABLED";
    FD1P3AX mepc_i0_i1 (.D(mepc[5]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i1.GSR = "DISABLED";
    PFUMX i28026 (.BLUT(debug_branch_N_840[30]), .ALUT(n30702), .C0(n29329), 
          .Z(n30703));
    FD1P3AX mepc_i0_i2 (.D(mepc[6]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i2.GSR = "DISABLED";
    FD1P3AX mepc_i0_i3 (.D(mepc[7]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i3.GSR = "DISABLED";
    FD1P3AX mepc_i0_i4 (.D(mepc[8]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i4.GSR = "DISABLED";
    FD1P3AX mepc_i0_i5 (.D(mepc[9]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i5.GSR = "DISABLED";
    FD1P3AX mepc_i0_i6 (.D(mepc[10]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i6.GSR = "DISABLED";
    FD1P3AX mepc_i0_i7 (.D(mepc[11]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i7.GSR = "DISABLED";
    FD1P3AX mepc_i0_i8 (.D(mepc[12]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i8.GSR = "DISABLED";
    FD1P3AX mepc_i0_i9 (.D(mepc[13]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i9.GSR = "DISABLED";
    FD1P3AX mepc_i0_i10 (.D(mepc[14]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i10.GSR = "DISABLED";
    FD1P3AX mepc_i0_i11 (.D(mepc[15]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i11.GSR = "DISABLED";
    FD1P3AX mepc_i0_i12 (.D(mepc[16]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i12.GSR = "DISABLED";
    FD1P3AX mepc_i0_i13 (.D(mepc[17]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i13.GSR = "DISABLED";
    FD1P3AX mepc_i0_i14 (.D(mepc[18]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i14.GSR = "DISABLED";
    FD1P3AX mepc_i0_i15 (.D(mepc[19]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i15.GSR = "DISABLED";
    FD1P3AX mepc_i0_i16 (.D(mepc[20]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i16.GSR = "DISABLED";
    FD1P3AX mepc_i0_i17 (.D(mepc[21]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i17.GSR = "DISABLED";
    FD1P3AX mepc_i0_i18 (.D(mepc[22]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i18.GSR = "DISABLED";
    FD1P3AX mepc_i0_i19 (.D(mepc[23]), .SP(clk_c_enable_543), .CK(clk_c), 
            .Q(mepc[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i19.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(\next_fsm_state_3__N_3015[3] ), .B(mie[2]), .Z(n31)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    FD1P3AX last_interrupt_req_i0_i1 (.D(\ui_in_sync[1] ), .SP(clk_c_enable_449), 
            .CK(clk_c), .Q(last_interrupt_req[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(419[12] 460[8])
    defparam last_interrupt_req_i0_i1.GSR = "DISABLED";
    LUT4 i1_3_lut (.A(n32046), .B(rd[1]), .C(rd[0]), .Z(n28210)) /* synthesis lut_function=(!((B (C)+!B !(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut.init = 16'h2828;
    LUT4 equal_3547_i6_2_lut_rep_776 (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .Z(n31981)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam equal_3547_i6_2_lut_rep_776.init = 16'hdddd;
    LUT4 i1_4_lut_adj_313 (.A(fsm_state[2]), .B(n32025), .C(fsm_state[0]), 
         .D(mie[3]), .Z(n10548)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_313.init = 16'h0100;
    LUT4 i15334_3_lut_4_lut (.A(\alu_op[0] ), .B(\alu_op[1] ), .C(n32004), 
         .D(n32005), .Z(clk_c_enable_544)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i15334_3_lut_4_lut.init = 16'hd0ff;
    LUT4 i8256_4_lut (.A(debug_instr_valid), .B(n28318), .C(is_lui), .D(is_jal), 
         .Z(n10873)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(218[17:110])
    defparam i8256_4_lut.init = 16'haaa8;
    LUT4 i1_2_lut_3_lut_4_lut_adj_314 (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .C(mip_reg[17]), .D(n31948), .Z(n28620)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i1_2_lut_3_lut_4_lut_adj_314.init = 16'hd0f0;
    LUT4 i16135_3_lut_4_lut_4_lut_4_lut (.A(\alu_op[0] ), .B(\alu_op[1] ), 
         .C(data_rs1_c[3]), .D(n31948), .Z(n18719)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(60[21:41])
    defparam i16135_3_lut_4_lut_4_lut_4_lut.init = 16'he200;
    LUT4 mie_3__bdd_4_lut_28446 (.A(mie[3]), .B(mie[11]), .C(counter_hi[3]), 
         .D(counter_hi[4]), .Z(n30989)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;
    defparam mie_3__bdd_4_lut_28446.init = 16'hcacc;
    LUT4 n30987_bdd_3_lut (.A(n30987), .B(mie[15]), .C(counter_hi[3]), 
         .Z(n30988)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30987_bdd_3_lut.init = 16'hcaca;
    LUT4 mie_15__bdd_3_lut (.A(mie[7]), .B(mie[16]), .C(counter_hi[4]), 
         .Z(n30987)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam mie_15__bdd_3_lut.init = 16'hacac;
    LUT4 i27839_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n31966), .D(counter_hi[2]), .Z(clk_c_enable_169)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(482[33:47])
    defparam i27839_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_adj_315 (.A(is_branch), .B(is_jalr), .C(is_auipc), .D(is_system), 
         .Z(n28318)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(218[17:110])
    defparam i1_4_lut_adj_315.init = 16'hfffe;
    LUT4 equal_110_i5_2_lut_rep_742_3_lut (.A(n33486), .B(n33484), .C(counter_hi[2]), 
         .Z(n31947)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(482[33:47])
    defparam equal_110_i5_2_lut_rep_742_3_lut.init = 16'hfbfb;
    LUT4 i27686_4_lut (.A(n31841), .B(n28558), .C(n31854), .D(n18719), 
         .Z(clk_c_enable_536)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i27686_4_lut.init = 16'hfbfa;
    LUT4 i27844_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n31966), .D(counter_hi[2]), .Z(clk_c_enable_165)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(482[33:47])
    defparam i27844_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i27936_2_lut_rep_778 (.A(\imm[5] ), .B(\imm[3] ), .Z(n31983)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i27936_2_lut_rep_778.init = 16'h1111;
    LUT4 i1_3_lut_4_lut_adj_316 (.A(\imm[5] ), .B(\imm[3] ), .C(\imm[2] ), 
         .D(\imm[0] ), .Z(n28518)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_316.init = 16'hfffe;
    LUT4 i1_4_lut_adj_317 (.A(n27528), .B(cmp_out), .C(n32015), .D(mem_op[0]), 
         .Z(n26597)) /* synthesis lut_function=(A+!(B ((D)+!C)+!B !(C (D)))) */ ;
    defparam i1_4_lut_adj_317.init = 16'hbaea;
    LUT4 i1_4_lut_adj_318 (.A(\alu_op_in[2] ), .B(n31987), .C(\alu_op[1] ), 
         .D(\alu_op[0] ), .Z(n26175)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_318.init = 16'h0004;
    LUT4 i1_4_lut_adj_319 (.A(n31938), .B(n31926), .C(n31955), .D(interrupt_core), 
         .Z(n27528)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_319.init = 16'hfffe;
    LUT4 mux_73_i1_4_lut (.A(cmp), .B(tmp_data[0]), .C(n32008), .D(n32005), 
         .Z(n196[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(170[18] 174[35])
    defparam mux_73_i1_4_lut.init = 16'hca0a;
    LUT4 mux_72_i1_4_lut (.A(accum[0]), .B(alu_out[0]), .C(n32004), .D(d_3__N_1868[0]), 
         .Z(n191[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(174[17:35])
    defparam mux_72_i1_4_lut.init = 16'hc5ca;
    LUT4 tmp_data_in_3__I_124_i2_3_lut (.A(tmp_data_in_3__N_1582[1]), .B(data_rs1_c[1]), 
         .C(n5737), .Z(tmp_data_in_3__N_1514[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_124_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_783 (.A(n33486), .B(counter_hi[4]), .Z(n31988)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i1_2_lut_rep_783.init = 16'heeee;
    LUT4 equal_109_i5_2_lut_rep_741_3_lut (.A(n33486), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(n31946)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam equal_109_i5_2_lut_rep_741_3_lut.init = 16'hefef;
    LUT4 i27879_2_lut_rep_724_3_lut_3_lut_4_lut_3_lut (.A(counter_hi[3]), 
         .B(counter_hi[4]), .C(counter_hi[2]), .Z(n31929)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i27879_2_lut_rep_724_3_lut_3_lut_4_lut_3_lut.init = 16'h0404;
    LUT4 i27848_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_done_N_1741), .D(counter_hi[2]), .Z(clk_c_enable_77)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i27848_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_adj_320 (.A(n26486), .B(debug_rd_3__N_1575), .C(counter_hi[4]), 
         .D(n28374), .Z(load_top_bit_next_N_1731)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_320.init = 16'h0400;
    LUT4 i23998_2_lut (.A(n33486), .B(mem_op[0]), .Z(n26486)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i23998_2_lut.init = 16'h6666;
    LUT4 i1_3_lut_4_lut_adj_321 (.A(counter_hi[3]), .B(counter_hi[4]), .C(timer_interrupt), 
         .D(counter_hi[2]), .Z(n27288)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i1_3_lut_4_lut_adj_321.init = 16'h1000;
    LUT4 i1_3_lut_adj_322 (.A(mem_op[2]), .B(mem_op[1]), .C(counter_hi[2]), 
         .Z(n28374)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_adj_322.init = 16'h1010;
    LUT4 i27831_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n31966), .D(counter_hi[2]), .Z(clk_c_enable_181)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i27831_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_744_3_lut (.A(n33486), .B(n33484), .C(counter_hi[2]), 
         .Z(n31949)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i1_2_lut_rep_744_3_lut.init = 16'hfefe;
    LUT4 mux_72_i2_3_lut (.A(\mul_out[1] ), .B(alu_out[1]), .C(n32004), 
         .Z(n191[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(174[17:35])
    defparam mux_72_i2_3_lut.init = 16'hcaca;
    LUT4 i15512_2_lut_rep_740_3_lut_4_lut (.A(n33486), .B(n33484), .C(cy_adj_3109), 
         .D(counter_hi[2]), .Z(n31945)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i15512_2_lut_rep_740_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i27853_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_top_bit_next_N_1731), .D(counter_hi[2]), .Z(n18685)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i27853_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i27689_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_done_N_1741), .D(counter_hi[2]), .Z(clk_c_enable_80)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i27689_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(load_top_bit_next_N_1731), .D(counter_hi[2]), .Z(clk_c_enable_545)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i1_3_lut_adj_323 (.A(\alu_op_in[2] ), .B(\alu_op[1] ), .C(\alu_op[3] ), 
         .Z(n10486)) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam i1_3_lut_adj_323.init = 16'hfbfb;
    LUT4 equal_106_i6_1_lut_rep_715_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .Z(clk_c_enable_249)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam equal_106_i6_1_lut_rep_715_2_lut_3_lut.init = 16'h0101;
    LUT4 i27746_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n31966), .D(counter_hi[2]), .Z(clk_c_enable_184)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i27746_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i3941_2_lut_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(mstatus_mte), .D(counter_hi[2]), .Z(n6096)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i3941_2_lut_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 debug_rd_3__I_0_i2_3_lut_4_lut (.A(n31956), .B(debug_rd_3__N_1575), 
         .C(debug_rd_3__N_1392[1]), .D(debug_rd_3__N_1571[1]), .Z(debug_rd[1])) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(176[18] 194[12])
    defparam debug_rd_3__I_0_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_716_3_lut_3_lut_4_lut_3_lut (.A(n33486), .B(n33484), 
         .C(counter_hi[2]), .Z(n31957)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i1_2_lut_rep_716_3_lut_3_lut_4_lut_3_lut.init = 16'h4040;
    LUT4 i27470_3_lut (.A(n32185), .B(\timer_data[0] ), .C(is_timer_addr), 
         .Z(debug_branch_N_840[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam i27470_3_lut.init = 16'hcaca;
    LUT4 mux_72_i3_3_lut (.A(\mul_out[2] ), .B(alu_out[2]), .C(n32004), 
         .Z(n191[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(174[17:35])
    defparam mux_72_i3_3_lut.init = 16'hcaca;
    LUT4 i27921_3_lut (.A(data_out_3__N_1385), .B(is_timer_addr), .C(n29318), 
         .Z(n29329)) /* synthesis lut_function=(A+!(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam i27921_3_lut.init = 16'habab;
    LUT4 tmp_data_in_3__I_124_i3_4_lut (.A(data_rs1_c[2]), .B(mstatus_mte), 
         .C(n31896), .D(n31893), .Z(tmp_data_in_3__N_1514[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(251[14] 256[36])
    defparam tmp_data_in_3__I_124_i3_4_lut.init = 16'hca0a;
    LUT4 n30945_bdd_4_lut (.A(n30945), .B(n30944), .C(counter_hi[2]), 
         .D(n4874), .Z(csr_read_3__N_1447[0])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n30945_bdd_4_lut.init = 16'hca00;
    PFUMX i28306 (.BLUT(csr_read_3__N_1447[3]), .ALUT(n31172), .C0(\imm[6] ), 
          .Z(n31173));
    LUT4 i27484_3_lut (.A(n31319), .B(\timer_data[2] ), .C(is_timer_addr), 
         .Z(debug_branch_N_840[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam i27484_3_lut.init = 16'hcaca;
    LUT4 mux_72_i4_3_lut (.A(\mul_out[3] ), .B(alu_out[3]), .C(n32004), 
         .Z(n191[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(174[17:35])
    defparam mux_72_i4_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_324 (.A(tmp_data[30]), .B(tmp_data[31]), .C(cycle[0]), 
         .Z(instr_complete_N_1656)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_adj_324.init = 16'hf7f7;
    LUT4 cycle_0__I_0_548_3_lut (.A(cycle[0]), .B(cmp_out), .C(\alu_op[0] ), 
         .Z(instr_complete_N_1654)) /* synthesis lut_function=(A+!(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(224[34:67])
    defparam cycle_0__I_0_548_3_lut.init = 16'hbebe;
    LUT4 is_jal_I_0_2_lut_rep_794 (.A(is_jal), .B(is_jalr), .Z(n31999)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam is_jal_I_0_2_lut_rep_794.init = 16'heeee;
    LUT4 mux_87_i4_3_lut (.A(\debug_branch_N_450[3] ), .B(load_top_bit), 
         .C(data_out_3__N_1385), .Z(debug_rd_3__N_1571[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(182[17:35])
    defparam mux_87_i4_3_lut.init = 16'hcaca;
    LUT4 i5743_2_lut_rep_750_3_lut (.A(is_jal), .B(is_jalr), .C(debug_instr_valid), 
         .Z(n31955)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(201[37:54])
    defparam i5743_2_lut_rep_750_3_lut.init = 16'he0e0;
    LUT4 mux_3526_i1_3_lut (.A(n31589), .B(n29158), .C(n5670), .Z(n5677[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3526_i1_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_325 (.A(n31948), .B(n46), .C(\imm[7] ), .Z(n9033)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(190[18] 194[12])
    defparam i1_3_lut_adj_325.init = 16'h0808;
    LUT4 i1_4_lut_adj_326 (.A(n26148), .B(n10727), .C(\imm[7] ), .D(\imm[11] ), 
         .Z(n5670)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_326.init = 16'h0008;
    LUT4 i1_4_lut_adj_327 (.A(\imm[1] ), .B(n31983), .C(\imm[0] ), .D(\imm[2] ), 
         .Z(n10727)) /* synthesis lut_function=(!(A+((C (D)+!C !(D))+!B))) */ ;
    defparam i1_4_lut_adj_327.init = 16'h0440;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(counter_hi[2]), .D(mip_reg[17]), .Z(csr_read_3__N_1459[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i1_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0400;
    LUT4 i7103_3_lut_rep_751_4_lut (.A(is_alu_imm), .B(is_alu_reg), .C(is_auipc), 
         .D(debug_instr_valid), .Z(n31956)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(225[22:46])
    defparam i7103_3_lut_rep_751_4_lut.init = 16'hfe00;
    LUT4 i5748_2_lut_3_lut (.A(is_alu_imm), .B(is_alu_reg), .C(debug_instr_valid), 
         .Z(debug_rd_3__N_1401)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(225[22:46])
    defparam i5748_2_lut_3_lut.init = 16'he0e0;
    FD1P3IX tmp_data_i0_i28 (.D(tmp_data_in_3__N_1514[0]), .SP(clk_c_enable_544), 
            .CD(n11557), .CK(clk_c), .Q(tmp_data[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i28.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_799 (.A(\alu_op[3] ), .B(\alu_op[1] ), .C(\alu_op_in[2] ), 
         .Z(n32004)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_rep_799.init = 16'hf7f7;
    PFUMX i28009 (.BLUT(n30667), .ALUT(n30665), .C0(n32008), .Z(n30668));
    LUT4 i27732_2_lut_rep_800 (.A(cycle[0]), .B(cycle[1]), .Z(n32005)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam i27732_2_lut_rep_800.init = 16'h2222;
    LUT4 n194_bdd_2_lut_28186_3_lut (.A(cycle[0]), .B(cycle[1]), .C(tmp_data[1]), 
         .Z(n30665)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam n194_bdd_2_lut_28186_3_lut.init = 16'h2020;
    LUT4 i15642_2_lut_3_lut (.A(cycle[0]), .B(cycle[1]), .C(tmp_data[3]), 
         .Z(debug_rd_3__N_1563[3])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam i15642_2_lut_3_lut.init = 16'h2020;
    LUT4 n193_bdd_2_lut_3_lut (.A(cycle[0]), .B(cycle[1]), .C(tmp_data[2]), 
         .Z(n30695)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(168[34:44])
    defparam n193_bdd_2_lut_3_lut.init = 16'h2020;
    LUT4 i1_3_lut_rep_803 (.A(\alu_op[1] ), .B(\alu_op_in[2] ), .C(\alu_op[3] ), 
         .Z(n32008)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_803.init = 16'h8080;
    LUT4 i5235_2_lut_rep_621_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in[2]), .Z(n31826)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i5235_2_lut_rep_621_4_lut_4_lut.init = 16'h857a;
    LUT4 i5236_2_lut_rep_622_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(\alu_b_in[3] ), .Z(n31827)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i5236_2_lut_rep_622_4_lut_4_lut.init = 16'h857a;
    LUT4 i15760_3_lut_rep_754_3_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .Z(n31959)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;
    defparam i15760_3_lut_rep_754_3_lut.init = 16'h7a7a;
    LUT4 i5220_2_lut_rep_620_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in[0]), .Z(n31825)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i5220_2_lut_rep_620_4_lut_4_lut.init = 16'h857a;
    LUT4 i27948_2_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), .C(\alu_op[3] ), 
         .D(debug_rd_3__N_413), .Z(n29243)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i27948_2_lut_4_lut.init = 16'hff80;
    LUT4 i5234_2_lut_rep_651_4_lut_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(alu_b_in[1]), .Z(n31856)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A !(C (D)+!C !(D))) */ ;
    defparam i5234_2_lut_rep_651_4_lut_4_lut.init = 16'h857a;
    LUT4 i15311_2_lut_rep_755_4_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .D(\alu_op[0] ), .Z(n31960)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;
    defparam i15311_2_lut_rep_755_4_lut.init = 16'h7f00;
    LUT4 i15637_2_lut_rep_774_3_lut (.A(\alu_op[1] ), .B(\alu_op_in[2] ), 
         .C(\alu_op[3] ), .Z(n31979)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i15637_2_lut_rep_774_3_lut.init = 16'h2a2a;
    LUT4 mux_3501_i4_4_lut_4_lut (.A(\imm[0] ), .B(\imm[1] ), .C(instrret_count[3]), 
         .D(\cycle_count_wide[3] ), .Z(n5624[3])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam mux_3501_i4_4_lut_4_lut.init = 16'h7340;
    LUT4 mux_3501_i3_4_lut_4_lut (.A(\imm[0] ), .B(\imm[1] ), .C(instrret_count[2]), 
         .D(cycle_count_wide[2]), .Z(n5626)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam mux_3501_i3_4_lut_4_lut.init = 16'h7340;
    LUT4 i1_3_lut_4_lut_adj_328 (.A(n31946), .B(n31874), .C(counter_hi[4]), 
         .D(n32049), .Z(clk_c_enable_258)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(429[18] 459[12])
    defparam i1_3_lut_4_lut_adj_328.init = 16'h2000;
    LUT4 i27784_2_lut_rep_806 (.A(\imm[1] ), .B(\imm[0] ), .Z(n32011)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i27784_2_lut_rep_806.init = 16'hbbbb;
    LUT4 i27792_2_lut_3_lut (.A(\imm[1] ), .B(\imm[0] ), .C(\imm[10] ), 
         .Z(n29539)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i27792_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i1_3_lut_4_lut_adj_329 (.A(n31875), .B(data_rs1[0]), .C(n29008), 
         .D(mie[12]), .Z(n928)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_329.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_330 (.A(n31875), .B(data_rs1[0]), .C(n29008), 
         .D(mie[8]), .Z(n895)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_330.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_331 (.A(n31875), .B(data_rs1[0]), .C(n29008), 
         .D(mie[4]), .Z(n862)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_331.init = 16'h8f88;
    LUT4 i1_4_lut_4_lut_adj_332 (.A(\imm[2] ), .B(n31983), .C(n40), .D(n28508), 
         .Z(n27180)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_4_lut_4_lut_adj_332.init = 16'h4000;
    LUT4 i1_3_lut_4_lut_adj_333 (.A(data_rs1_c[1]), .B(n31875), .C(n8_adj_3110), 
         .D(mie[13]), .Z(n927)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_333.init = 16'h8f88;
    LUT4 i1_2_lut_rep_809 (.A(\imm[9] ), .B(\imm[8] ), .Z(n32014)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_809.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_334 (.A(data_rs1_c[1]), .B(n31875), .C(n8_adj_3110), 
         .D(mie[9]), .Z(n894)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_334.init = 16'h8f88;
    LUT4 i1_2_lut_rep_721_3_lut (.A(\imm[9] ), .B(\imm[8] ), .C(n26175), 
         .Z(n31926)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_721_3_lut.init = 16'h8080;
    LUT4 i1_3_lut_4_lut_adj_335 (.A(data_rs1_c[1]), .B(n31875), .C(n8_adj_3110), 
         .D(mie[5]), .Z(n861)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_335.init = 16'h8f88;
    LUT4 i15650_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[30]), 
         .D(n26175), .Z(\addr_out[26] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i15650_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i1_3_lut_4_lut_adj_336 (.A(\imm[9] ), .B(\imm[8] ), .C(\imm[4] ), 
         .D(\imm[10] ), .Z(n26148)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_336.init = 16'h0008;
    LUT4 i15649_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[29]), 
         .D(n26175), .Z(\addr_out[25] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i15649_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i1_3_lut_4_lut_adj_337 (.A(data_rs1_c[1]), .B(n31875), .C(n8_adj_3110), 
         .D(mie[1]), .Z(n794)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_4_lut_adj_337.init = 16'h8f88;
    LUT4 i15648_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[28]), 
         .D(n26175), .Z(\addr_out[24] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i15648_2_lut_3_lut_4_lut.init = 16'h70f0;
    FD1P3IX mepc_i0_i23 (.D(n658[3]), .SP(clk_c_enable_543), .CD(n11559), 
            .CK(clk_c), .Q(mepc[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i23.GSR = "DISABLED";
    FD1P3IX mepc_i0_i22 (.D(n658[2]), .SP(clk_c_enable_543), .CD(n11559), 
            .CK(clk_c), .Q(mepc[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i22.GSR = "DISABLED";
    FD1P3IX mepc_i0_i21 (.D(n658[1]), .SP(clk_c_enable_543), .CD(n11559), 
            .CK(clk_c), .Q(mepc[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i21.GSR = "DISABLED";
    LUT4 i15651_2_lut_3_lut_4_lut (.A(\imm[9] ), .B(\imm[8] ), .C(tmp_data[31]), 
         .D(n26175), .Z(\addr_out[27] )) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;
    defparam i15651_2_lut_3_lut_4_lut.init = 16'h70f0;
    LUT4 i1_3_lut_4_lut_adj_338 (.A(n31875), .B(data_rs1_c[3]), .C(n20), 
         .D(mie[16]), .Z(n25282)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_338.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_339 (.A(n31875), .B(data_rs1_c[3]), .C(n20), 
         .D(mie[15]), .Z(n25292)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_339.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_340 (.A(n31875), .B(data_rs1_c[3]), .C(n20), 
         .D(mie[11]), .Z(n25290)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_340.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_341 (.A(n31875), .B(data_rs1_c[3]), .C(n20), 
         .D(mie[7]), .Z(n25288)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_341.init = 16'h8f88;
    LUT4 i1_3_lut_4_lut_adj_342 (.A(n31875), .B(data_rs1_c[3]), .C(n20), 
         .D(mie[3]), .Z(n25284)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam i1_3_lut_4_lut_adj_342.init = 16'h8f88;
    LUT4 mstatus_mie_I_153_3_lut_4_lut (.A(n31875), .B(data_rs1_c[3]), .C(n31926), 
         .D(mstatus_mpie), .Z(mstatus_mie_N_1709)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(406[22] 407[72])
    defparam mstatus_mie_I_153_3_lut_4_lut.init = 16'hf808;
    FD1P3AX mstatus_mie_524 (.D(mstatus_mie_N_1707), .SP(clk_c_enable_536), 
            .CK(clk_c), .Q(mstatus_mie)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam mstatus_mie_524.GSR = "DISABLED";
    LUT4 mux_3526_i4_3_lut (.A(n29155), .B(n31174), .C(n5670), .Z(n5677[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam mux_3526_i4_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_343 (.A(stall_core), .B(instr_complete_N_1647), .C(clk_c_enable_36), 
         .D(n28210), .Z(n26997)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_343.init = 16'h8000;
    LUT4 i1_4_lut_adj_344 (.A(stall_core), .B(instr_complete_N_1647), .C(clk_c_enable_36), 
         .D(n28222), .Z(n26995)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_344.init = 16'h8000;
    LUT4 mux_327_i1_4_lut (.A(n31894), .B(data_rs1[0]), .C(n31892), .D(mip_reg[16]), 
         .Z(n809[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(437[22:76])
    defparam mux_327_i1_4_lut.init = 16'hf2c0;
    LUT4 i1_4_lut_adj_345 (.A(stall_core), .B(instr_complete_N_1647), .C(n31917), 
         .D(n109), .Z(n26996)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_345.init = 16'h8000;
    LUT4 i1_2_lut_rep_818 (.A(mip_reg[17]), .B(mie[1]), .Z(n32023)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(321[17:24])
    defparam i1_2_lut_rep_818.init = 16'h8888;
    LUT4 and_454_i1_2_lut_rep_819 (.A(mip_reg[16]), .B(mie[0]), .Z(n32024)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[48:59])
    defparam and_454_i1_2_lut_rep_819.init = 16'h8888;
    LUT4 i1_2_lut_rep_768_3_lut_4_lut (.A(mip_reg[16]), .B(mie[0]), .C(mie[1]), 
         .D(mip_reg[17]), .Z(n31973)) /* synthesis lut_function=(A (B+(C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[48:59])
    defparam i1_2_lut_rep_768_3_lut_4_lut.init = 16'hf888;
    LUT4 i26322_2_lut_rep_820 (.A(fsm_state[1]), .B(fsm_state[3]), .Z(n32025)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26322_2_lut_rep_820.init = 16'heeee;
    LUT4 i1_2_lut_rep_758_3_lut (.A(fsm_state[1]), .B(fsm_state[3]), .C(fsm_state[2]), 
         .Z(n31963)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_758_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_727_3_lut_4_lut (.A(fsm_state[1]), .B(fsm_state[3]), 
         .C(fsm_state[0]), .D(fsm_state[2]), .Z(n31932)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_727_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_346 (.A(fsm_state[1]), .B(fsm_state[3]), 
         .C(next_bit), .D(fsm_state[2]), .Z(n28800)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_346.init = 16'hf0e0;
    LUT4 i27373_3_lut_4_lut (.A(\imm[10] ), .B(\imm[1] ), .C(n31690), 
         .D(n29171), .Z(n5671[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(468[9] 512[16])
    defparam i27373_3_lut_4_lut.init = 16'hf2d0;
    FD1P3IX mepc_i0_i20 (.D(n658[0]), .SP(clk_c_enable_543), .CD(n11559), 
            .CK(clk_c), .Q(mepc[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(367[12] 375[8])
    defparam mepc_i0_i20.GSR = "DISABLED";
    FD1S3AX cycle__i0 (.D(n31389), .CK(clk_c), .Q(cycle[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(206[12] 212[8])
    defparam cycle__i0.GSR = "DISABLED";
    LUT4 i15336_2_lut (.A(\data_rs2[0] ), .B(data_out_3__N_1385), .Z(\data_out_slice[0] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i15336_2_lut.init = 16'h2222;
    LUT4 i8257_4_lut (.A(mem_op[1]), .B(mem_op[0]), .C(n33484), .D(n33486), 
         .Z(data_out_3__N_1385)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[13] 272[50])
    defparam i8257_4_lut.init = 16'h5150;
    LUT4 n194_bdd_4_lut_28187 (.A(n191[1]), .B(shift_out[1]), .C(n32005), 
         .D(n31981), .Z(n30666)) /* synthesis lut_function=(A (B+((D)+!C))+!A !(((D)+!C)+!B)) */ ;
    defparam n194_bdd_4_lut_28187.init = 16'haaca;
    FD1P3IX tmp_data_i0_i29 (.D(tmp_data_in_3__N_1514[1]), .SP(clk_c_enable_544), 
            .CD(n11557), .CK(clk_c), .Q(tmp_data[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(262[12] 265[8])
    defparam tmp_data_i0_i29.GSR = "DISABLED";
    LUT4 is_load_I_0_2_lut (.A(is_load), .B(is_store), .Z(n9710)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(237[58:79])
    defparam is_load_I_0_2_lut.init = 16'heeee;
    FD1P3IX load_top_bit_513 (.D(\debug_branch_N_450[3] ), .SP(clk_c_enable_545), 
            .CD(n18685), .CK(clk_c), .Q(load_top_bit)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(156[12] 157[43])
    defparam load_top_bit_513.GSR = "DISABLED";
    LUT4 equal_108_i3_2_lut (.A(cycle[0]), .B(cycle[1]), .Z(load_done_N_1741)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(237[42:54])
    defparam equal_108_i3_2_lut.init = 16'heeee;
    LUT4 imm_10__bdd_3_lut_3_lut_4_lut (.A(n31988), .B(counter_hi[2]), .C(\imm[1] ), 
         .D(mcause[1]), .Z(n31689)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam imm_10__bdd_3_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 gnd_bdd_2_lut_28015 (.A(n30666), .B(n15), .Z(n30667)) /* synthesis lut_function=(A (B)) */ ;
    defparam gnd_bdd_2_lut_28015.init = 16'h8888;
    LUT4 i26577_3_lut_3_lut (.A(counter_hi[4]), .B(n29739), .C(n13), .Z(n29194)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i26577_3_lut_3_lut.init = 16'he4e4;
    PFUMX debug_rd_3__I_122_i4 (.BLUT(debug_rd_3__N_1571[3]), .ALUT(debug_rd_3__N_1396[3]), 
          .C0(n31956), .Z(debug_rd_3__N_1392[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    L6MUX21 instr_complete_I_131 (.D0(instr_complete_N_1650), .D1(instr_complete_N_1649), 
            .SD(n29243), .Z(instr_complete_N_1648)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX instr_complete_I_132 (.BLUT(instr_complete_N_1654), .ALUT(instr_complete_N_1656), 
          .C0(debug_rd_3__N_413), .Z(instr_complete_N_1649)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 n29137_bdd_3_lut_28190 (.A(n29137), .B(n234[1]), .C(n29330), 
         .Z(n30669)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n29137_bdd_3_lut_28190.init = 16'hacac;
    PFUMX tmp_data_in_3__I_0_i4 (.BLUT(tmp_data_in_3__N_1582[3]), .ALUT(tmp_data_in_3__N_1514[3]), 
          .C0(n29351), .Z(tmp_data_in[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 n30669_bdd_3_lut_28013 (.A(n30669), .B(n30668), .C(n31956), .Z(debug_rd_3__N_1392[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30669_bdd_3_lut_28013.init = 16'hcaca;
    LUT4 debug_branch_N_840_30__bdd_4_lut (.A(n30696), .B(n30695), .C(n15), 
         .D(n32008), .Z(n30701)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (B (D))) */ ;
    defparam debug_branch_N_840_30__bdd_4_lut.init = 16'hcca0;
    L6MUX21 debug_rd_3__I_122_i1 (.D0(debug_rd_3__N_1567[0]), .D1(debug_rd_3__N_1571[0]), 
            .SD(debug_rd_3__N_1575), .Z(debug_rd_3__N_1392[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX tmp_data_in_3__I_0_i3 (.BLUT(tmp_data_in_3__N_1582[2]), .ALUT(tmp_data_in_3__N_1514[2]), 
          .C0(n29351), .Z(tmp_data_in[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 n31173_bdd_3_lut (.A(n31173), .B(n31171), .C(\imm[0] ), .Z(n31174)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31173_bdd_3_lut.init = 16'hcaca;
    LUT4 i5190_2_lut (.A(\imm[6] ), .B(\imm[1] ), .Z(n7754)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i5190_2_lut.init = 16'h6666;
    PFUMX mux_87_i1 (.BLUT(debug_branch_N_840[28]), .ALUT(\debug_branch_N_450[0] ), 
          .C0(n29329), .Z(debug_rd_3__N_1571[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_2_lut_adj_347 (.A(\imm[6] ), .B(\imm[10] ), .Z(n28508)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_347.init = 16'h4444;
    LUT4 i67_4_lut (.A(n18076), .B(n32014), .C(\imm[4] ), .D(n32044), 
         .Z(n40)) /* synthesis lut_function=(A (B (C))+!A !(C+(D))) */ ;
    defparam i67_4_lut.init = 16'h8085;
    LUT4 i15495_2_lut_rep_834 (.A(counter_hi[3]), .B(counter_hi[2]), .Z(n32039)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15495_2_lut_rep_834.init = 16'heeee;
    LUT4 debug_branch_N_840_30__bdd_3_lut (.A(n29190), .B(data_out_3__N_1385), 
         .C(load_top_bit), .Z(n30702)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam debug_branch_N_840_30__bdd_3_lut.init = 16'he2e2;
    LUT4 i15509_2_lut (.A(\imm[1] ), .B(\imm[0] ), .Z(n18076)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15509_2_lut.init = 16'h8888;
    LUT4 n29149_bdd_3_lut_28744 (.A(n29149), .B(n234[2]), .C(n29330), 
         .Z(n30699)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n29149_bdd_3_lut_28744.init = 16'hacac;
    PFUMX mux_93_i1 (.BLUT(\debug_branch_N_446[28] ), .ALUT(n238), .C0(n29240), 
          .Z(debug_rd_3__N_1567[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX debug_rd_3__I_121_i1 (.BLUT(shift_out[0]), .ALUT(debug_rd_3__N_1559[0]), 
          .C0(n29550), .Z(debug_rd_3__N_1396[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 csr_read_3__N_1447_3__bdd_4_lut (.A(n31932), .B(n31949), .C(n27288), 
         .D(n31947), .Z(n31172)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C+!(D)))) */ ;
    defparam csr_read_3__N_1447_3__bdd_4_lut.init = 16'hc044;
    LUT4 data_ready_sync_I_0_3_lut_4_lut (.A(n31988), .B(counter_hi[2]), 
         .C(n31768), .D(data_ready_sync), .Z(data_ready_core)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam data_ready_sync_I_0_3_lut_4_lut.init = 16'hfe10;
    LUT4 n193_bdd_4_lut_28741 (.A(n191[2]), .B(shift_out[2]), .C(n32005), 
         .D(n31981), .Z(n30696)) /* synthesis lut_function=(A (B+((D)+!C))+!A !(((D)+!C)+!B)) */ ;
    defparam n193_bdd_4_lut_28741.init = 16'haaca;
    LUT4 i15902_2_lut_rep_839 (.A(\imm[8] ), .B(\imm[9] ), .Z(n32044)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15902_2_lut_rep_839.init = 16'heeee;
    LUT4 i1_2_lut_rep_733_3_lut (.A(\imm[8] ), .B(\imm[9] ), .C(n26175), 
         .Z(n31938)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_733_3_lut.init = 16'h1010;
    LUT4 i15341_2_lut_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), .C(n10513), 
         .D(n26175), .Z(n5054[0])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i15341_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 is_trap_I_0_586_2_lut_rep_691_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), 
         .C(interrupt_core), .D(n26175), .Z(n31896)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam is_trap_I_0_586_2_lut_rep_691_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i1_2_lut_rep_704_3_lut_4_lut (.A(\imm[8] ), .B(\imm[9] ), .C(interrupt_core), 
         .D(n26175), .Z(n31909)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i1_2_lut_rep_704_3_lut_4_lut.init = 16'hf1f0;
    LUT4 and_454_i17_2_lut_rep_840 (.A(timer_interrupt), .B(mie[16]), .Z(n32045)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[48:59])
    defparam and_454_i17_2_lut_rep_840.init = 16'h8888;
    LUT4 i15655_2_lut_3_lut (.A(timer_interrupt), .B(mie[16]), .C(interrupt_core), 
         .Z(n611[2])) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[48:59])
    defparam i15655_2_lut_3_lut.init = 16'h8080;
    LUT4 i15656_2_lut_3_lut (.A(timer_interrupt), .B(mie[16]), .C(interrupt_core), 
         .Z(n611[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[48:59])
    defparam i15656_2_lut_3_lut.init = 16'h7070;
    LUT4 i15420_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[20] ), 
         .D(\next_pc_for_core[16] ), .Z(n225)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i15420_4_lut_4_lut.init = 16'h5140;
    LUT4 c_2__N_1861_1__bdd_4_lut_28049_4_lut (.A(n33486), .B(counter_hi[2]), 
         .C(\pc[23] ), .D(\pc[19] ), .Z(n30741)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam c_2__N_1861_1__bdd_4_lut_28049_4_lut.init = 16'h5140;
    LUT4 c_2__N_1861_1__bdd_4_lut_4_lut (.A(n33486), .B(counter_hi[2]), 
         .C(\pc[21] ), .D(\pc[17] ), .Z(n30802)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam c_2__N_1861_1__bdd_4_lut_4_lut.init = 16'h5140;
    LUT4 i1_3_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(n33484), 
         .Z(n4874)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i1_3_lut_3_lut.init = 16'hf4f4;
    LUT4 i15422_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[22] ), 
         .D(\next_pc_for_core[18] ), .Z(n227)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i15422_4_lut_4_lut.init = 16'h5140;
    LUT4 i15399_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\pc[20] ), 
         .D(\pc[16] ), .Z(n225_adj_1)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i15399_4_lut_4_lut.init = 16'h5140;
    LUT4 c_2__N_1861_1__bdd_4_lut_28083_4_lut (.A(n33486), .B(counter_hi[2]), 
         .C(\pc[22] ), .D(\pc[18] ), .Z(n30746)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam c_2__N_1861_1__bdd_4_lut_28083_4_lut.init = 16'h5140;
    LUT4 i15421_4_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[2]), .C(\next_pc_for_core[21] ), 
         .D(\next_pc_for_core[17] ), .Z(n226)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[44:52])
    defparam i15421_4_lut_4_lut.init = 16'h5140;
    LUT4 csr_read_3__N_1463_1__bdd_3_lut_28534_3_lut_4_lut (.A(n31988), .B(counter_hi[2]), 
         .C(\cycle_count_wide[3] ), .D(\imm[1] ), .Z(n31586)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam csr_read_3__N_1463_1__bdd_3_lut_28534_3_lut_4_lut.init = 16'h11f0;
    LUT4 i15663_4_lut (.A(data_rs1_c[3]), .B(n32008), .C(\debug_branch_N_442[31] ), 
         .D(alu_a_in_3__N_1552), .Z(alu_a_in[3])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i15663_4_lut.init = 16'h3022;
    LUT4 i15662_4_lut (.A(data_rs1_c[2]), .B(n32008), .C(\debug_branch_N_442[30] ), 
         .D(alu_a_in_3__N_1552), .Z(alu_a_in[2])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i15662_4_lut.init = 16'h3022;
    LUT4 imm_3__I_0_i3_3_lut (.A(\debug_rd_3__N_405[30] ), .B(\data_rs2[2] ), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 imm_3__I_0_i2_3_lut (.A(\debug_rd_3__N_405[29] ), .B(\data_rs2[1] ), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 i15358_4_lut (.A(n157), .B(n32008), .C(\debug_branch_N_442[28] ), 
         .D(n29220), .Z(alu_a_in[0])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i15358_4_lut.init = 16'h2230;
    LUT4 imm_3__I_0_i1_3_lut (.A(\debug_rd_3__N_405[28] ), .B(\data_rs2[0] ), 
         .C(alu_b_in_3__N_1504), .Z(alu_b_in[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:69])
    defparam imm_3__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 i5733_3_lut (.A(debug_instr_valid), .B(is_alu_reg), .C(is_branch), 
         .Z(alu_b_in_3__N_1504)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(109[27:52])
    defparam i5733_3_lut.init = 16'ha8a8;
    LUT4 i5732_3_lut (.A(debug_instr_valid), .B(is_auipc), .C(is_jal), 
         .Z(alu_a_in_3__N_1552)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(108[27:47])
    defparam i5732_3_lut.init = 16'ha8a8;
    LUT4 i15661_4_lut (.A(data_rs1_c[1]), .B(n32008), .C(\debug_branch_N_442[29] ), 
         .D(alu_a_in_3__N_1552), .Z(alu_a_in[1])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(107[27] 108[63])
    defparam i15661_4_lut.init = 16'h3022;
    LUT4 i1_2_lut_rep_688_3_lut_4_lut (.A(n31988), .B(counter_hi[2]), .C(n26175), 
         .D(n32044), .Z(n31893)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam i1_2_lut_rep_688_3_lut_4_lut.init = 16'h0010;
    LUT4 csr_read_3__N_1463_1__bdd_3_lut_28605 (.A(cycle_count_wide[0]), .B(instrret_count[0]), 
         .C(\imm[1] ), .Z(n31587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam csr_read_3__N_1463_1__bdd_3_lut_28605.init = 16'hcaca;
    PFUMX mux_91_i3 (.BLUT(n29147), .ALUT(\debug_branch_N_446[30] ), .C0(n29333), 
          .Z(n234[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    PFUMX mux_91_i2 (.BLUT(n29135), .ALUT(\debug_branch_N_446[29] ), .C0(n29333), 
          .Z(n234[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_adj_348 (.A(\imm[2] ), .B(n31891), .C(n31947), 
         .D(n31946), .Z(clk_c_enable_274)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_2_lut_3_lut_4_lut_adj_348.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_349 (.A(\imm[2] ), .B(n31891), .C(n15604), 
         .D(n31946), .Z(clk_c_enable_264)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_2_lut_3_lut_4_lut_adj_349.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_adj_350 (.A(\imm[2] ), .B(n31891), .C(n31947), 
         .D(n31957), .Z(clk_c_enable_269)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(480[13:20])
    defparam i1_3_lut_4_lut_adj_350.init = 16'h2000;
    LUT4 i15653_2_lut (.A(\data_rs2[2] ), .B(data_out_3__N_1385), .Z(\data_out_slice[2] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i15653_2_lut.init = 16'h2222;
    LUT4 i15652_2_lut (.A(\data_rs2[1] ), .B(data_out_3__N_1385), .Z(\data_out_slice[1] )) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(271[9] 273[26])
    defparam i15652_2_lut.init = 16'h2222;
    PFUMX i27966 (.BLUT(n30580), .ALUT(n33494), .C0(n31915), .Z(n30581));
    LUT4 n30699_bdd_3_lut (.A(n30699), .B(n30703), .C(debug_rd_3__N_1575), 
         .Z(n30704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30699_bdd_3_lut.init = 16'hcaca;
    PFUMX mux_443_i1 (.BLUT(n822[0]), .ALUT(n948[0]), .C0(n31947), .Z(n979[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 data_rs1_3__I_0_i1_2_lut (.A(data_rs1[0]), .B(cycle[0]), .Z(mul_out_3__N_1510[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i1_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i2_2_lut (.A(data_rs1_c[1]), .B(cycle[0]), .Z(mul_out_3__N_1510[1])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i2_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_351 (.A(n31909), .B(n31972), .C(n10873), .D(instr_complete_N_1648), 
         .Z(instr_complete_N_1647)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i1_3_lut_4_lut_adj_351.init = 16'hfffe;
    LUT4 data_rs1_3__I_0_i3_2_lut (.A(data_rs1_c[2]), .B(cycle[0]), .Z(mul_out_3__N_1510[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i3_2_lut.init = 16'h8888;
    LUT4 data_rs1_3__I_0_i4_2_lut (.A(data_rs1_c[3]), .B(cycle[0]), .Z(mul_out_3__N_1510[3])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[47:71])
    defparam data_rs1_3__I_0_i4_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_686 (.A(\imm[6] ), .B(n26019), .Z(n31891)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_686.init = 16'heeee;
    PFUMX i34 (.BLUT(n21), .ALUT(n17438), .C0(n31947), .Z(n25168));
    LUT4 i1_2_lut_rep_669_3_lut (.A(\imm[6] ), .B(n26019), .C(\imm[2] ), 
         .Z(n31874)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_669_3_lut.init = 16'hefef;
    LUT4 i1_3_lut_4_lut_adj_352 (.A(\imm[6] ), .B(n26019), .C(\imm[2] ), 
         .D(n31949), .Z(n28558)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_352.init = 16'hfffe;
    LUT4 i27837_2_lut_3_lut_4_lut (.A(\imm[6] ), .B(n26019), .C(n31946), 
         .D(\imm[2] ), .Z(clk_c_enable_252)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i27837_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_637_3_lut_4_lut (.A(\alu_op[0] ), .B(n31914), .C(data_rs1_c[1]), 
         .D(n31915), .Z(n31842)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_637_3_lut_4_lut.init = 16'hf040;
    LUT4 i8880_2_lut_rep_638_3_lut_4_lut (.A(\alu_op[0] ), .B(n31914), .C(data_rs1_c[3]), 
         .D(n31915), .Z(n31843)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i8880_2_lut_rep_638_3_lut_4_lut.init = 16'hf040;
    LUT4 i1_2_lut_3_lut_4_lut_adj_353 (.A(\alu_op[0] ), .B(n31914), .C(data_rs1_c[2]), 
         .D(n31915), .Z(n21568)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_353.init = 16'hf040;
    LUT4 n31312_bdd_3_lut (.A(n31312), .B(\timer_data[1] ), .C(is_timer_addr), 
         .Z(n31313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n31312_bdd_3_lut.init = 16'hcaca;
    LUT4 is_double_fault_I_0_3_lut_rep_671_4_lut (.A(n31949), .B(n31938), 
         .C(is_double_fault_r), .D(mstatus_mte), .Z(n31876)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(248[27:99])
    defparam is_double_fault_I_0_3_lut_rep_671_4_lut.init = 16'hf0f4;
    LUT4 i25_3_lut_4_lut (.A(\alu_op[0] ), .B(n31914), .C(data_rs1_c[3]), 
         .D(n31915), .Z(n20)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i25_3_lut_4_lut.init = 16'h8f80;
    LUT4 i13_3_lut_4_lut (.A(\alu_op[0] ), .B(n31914), .C(data_rs1_c[1]), 
         .D(n31915), .Z(n8_adj_3110)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i13_3_lut_4_lut.init = 16'h8f80;
    LUT4 i26448_3_lut_4_lut (.A(\alu_op[0] ), .B(n31914), .C(data_rs1[0]), 
         .D(n31915), .Z(n29008)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i26448_3_lut_4_lut.init = 16'hff80;
    LUT4 i13_3_lut_4_lut_adj_354 (.A(\alu_op[0] ), .B(n31914), .C(data_rs1_c[2]), 
         .D(n31915), .Z(n8_adj_3112)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i13_3_lut_4_lut_adj_354.init = 16'h8f80;
    LUT4 n13_bdd_3_lut_28386 (.A(\mem_data_from_read[17] ), .B(counter_hi[2]), 
         .C(\mem_data_from_read[21] ), .Z(n31310)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n13_bdd_3_lut_28386.init = 16'he2e2;
    LUT4 i26404_2_lut_rep_649_3_lut_4_lut (.A(n31938), .B(interrupt_core), 
         .C(n31926), .D(n31949), .Z(n31854)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i26404_2_lut_rep_649_3_lut_4_lut.init = 16'hf0fe;
    LUT4 mux_252_i2_3_lut_4_lut (.A(n31938), .B(interrupt_core), .C(\debug_branch_N_442[29] ), 
         .D(n653[1]), .Z(n658[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i3_3_lut_4_lut (.A(n31938), .B(interrupt_core), .C(\debug_branch_N_442[30] ), 
         .D(n653[2]), .Z(n658[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_252_i4_3_lut_4_lut (.A(n31938), .B(interrupt_core), .C(\debug_branch_N_442[31] ), 
         .D(n653[3]), .Z(n658[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam mux_252_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4546_3_lut (.A(time_hi[2]), .B(time_hi[1]), .C(time_hi[0]), 
         .Z(n498[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(295[55:71])
    defparam i4546_3_lut.init = 16'h6a6a;
    L6MUX21 mux_3526_i3 (.D0(n5671[2]), .D1(n29164), .SD(n5670), .Z(n5677[2]));
    PFUMX mux_3526_i2 (.BLUT(n5671[1]), .ALUT(n5665[1]), .C0(n5670), .Z(n5677[1]));
    LUT4 i4539_2_lut (.A(time_hi[1]), .B(time_hi[0]), .Z(n498[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(295[55:71])
    defparam i4539_2_lut.init = 16'h6666;
    LUT4 i4425_2_lut_4_lut (.A(tmp_data[6]), .B(mepc[2]), .C(n31926), 
         .D(\addr_offset[2] ), .Z(n701)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(267[23:65])
    defparam i4425_2_lut_4_lut.init = 16'h35ca;
    PFUMX mux_252_i1 (.BLUT(n653[0]), .ALUT(n29012), .C0(n31896), .Z(n658[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    L6MUX21 i26538 (.D0(n29153), .D1(n29154), .SD(\imm[10] ), .Z(n29155));
    L6MUX21 i26541 (.D0(n29156), .D1(n29157), .SD(\imm[0] ), .Z(n29158));
    PFUMX i26547 (.BLUT(n29162), .ALUT(n29163), .C0(\imm[0] ), .Z(n29164));
    LUT4 debug_rd_3__N_1575_bdd_4_lut_28707 (.A(n31948), .B(n31999), .C(debug_instr_valid), 
         .D(is_lui), .Z(n31352)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam debug_rd_3__N_1575_bdd_4_lut_28707.init = 16'hfaea;
    LUT4 n31352_bdd_2_lut (.A(n31352), .B(debug_rd_3__N_1575), .Z(n31353)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n31352_bdd_2_lut.init = 16'heeee;
    LUT4 debug_rd_3__N_1575_bdd_4_lut_28408 (.A(\alu_op[3] ), .B(\alu_op[1] ), 
         .C(\alu_op_in[2] ), .D(cycle[0]), .Z(n31351)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam debug_rd_3__N_1575_bdd_4_lut_28408.init = 16'hfff7;
    LUT4 i1_4_lut_adj_355 (.A(n10513), .B(n31938), .C(\debug_rd_3__N_405[28] ), 
         .D(interrupt_core), .Z(n27308)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_355.init = 16'h0004;
    LUT4 i1_3_lut_adj_356 (.A(\debug_rd_3__N_405[30] ), .B(\debug_rd_3__N_405[29] ), 
         .C(\debug_rd_3__N_405[31] ), .Z(n10513)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(353[26:40])
    defparam i1_3_lut_adj_356.init = 16'hfefe;
    LUT4 i1_4_lut_adj_357 (.A(n31841), .B(n29010), .C(n31878), .D(n18719), 
         .Z(clk_c_enable_250)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;
    defparam i1_4_lut_adj_357.init = 16'hfbfa;
    LUT4 i26450_4_lut (.A(n31926), .B(n31891), .C(n31946), .D(\imm[2] ), 
         .Z(n29010)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i26450_4_lut.init = 16'hfffe;
    LUT4 i15218_4_lut (.A(n31843), .B(n31841), .C(mstatus_mie), .D(n31878), 
         .Z(n6337)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(394[12] 414[8])
    defparam i15218_4_lut.init = 16'h3022;
    LUT4 i1_4_lut_adj_358 (.A(n32045), .B(n10548), .C(n31973), .D(n31), 
         .Z(n15837)) /* synthesis lut_function=(A+!(B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(331[17] 350[24])
    defparam i1_4_lut_adj_358.init = 16'hafae;
    LUT4 i1_3_lut_adj_359 (.A(mie[14]), .B(n21568), .C(n8_adj_3112), .Z(n926)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_359.init = 16'hcece;
    LUT4 i27684_3_lut_4_lut (.A(n31938), .B(interrupt_core), .C(n31949), 
         .D(rst_reg_n), .Z(clk_c_enable_251)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(66[25:48])
    defparam i27684_3_lut_4_lut.init = 16'h0eff;
    LUT4 i1_3_lut_adj_360 (.A(mie[10]), .B(n21568), .C(n8_adj_3112), .Z(n893)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_360.init = 16'hcece;
    LUT4 i1_3_lut_adj_361 (.A(mie[6]), .B(n21568), .C(n8_adj_3112), .Z(n860)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_361.init = 16'hcece;
    LUT4 i1_3_lut_adj_362 (.A(mie[2]), .B(n21568), .C(n8_adj_3112), .Z(n793)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(77[10:22])
    defparam i1_3_lut_adj_362.init = 16'hcece;
    PFUMX mux_233_i1 (.BLUT(n5054[0]), .ALUT(n27061), .C0(interrupt_core), 
          .Z(n611[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 i1_3_lut_rep_537_4_lut (.A(clk_c_enable_36), .B(n32046), .C(instr_complete_N_1647), 
         .D(stall_core), .Z(n31742)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_rep_537_4_lut.init = 16'h8000;
    PFUMX mux_3506_i2 (.BLUT(csr_read_3__N_1447[1]), .ALUT(csr_read_3__N_1459[1]), 
          .C0(\imm[6] ), .Z(n5633[1]));
    LUT4 tmp_data_in_3__I_124_i4_4_lut_4_lut_4_lut (.A(n31949), .B(data_rs1_c[3]), 
         .C(interrupt_core), .D(n31938), .Z(tmp_data_in_3__N_1514[3])) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam tmp_data_in_3__I_124_i4_4_lut_4_lut_4_lut.init = 16'h505c;
    LUT4 i4783_2_lut_rep_668_4_lut_4_lut (.A(n31949), .B(instrret_count[0]), 
         .C(instr_retired), .D(cy_c), .Z(n31873)) /* synthesis lut_function=(A (B (D))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i4783_2_lut_rep_668_4_lut_4_lut.init = 16'hc840;
    LUT4 cy_I_0_3_lut_rep_684_4_lut_4_lut (.A(n31949), .B(cy), .C(time_pulse_r), 
         .D(n10573), .Z(n31889)) /* synthesis lut_function=(A (B)+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam cy_I_0_3_lut_rep_684_4_lut_4_lut.init = 16'hd8dd;
    LUT4 i15915_4_lut_4_lut (.A(n31949), .B(\imm[1] ), .C(mcause[2]), 
         .D(mstatus_mte), .Z(n9538)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i15915_4_lut_4_lut.init = 16'h5140;
    LUT4 i4846_2_lut_rep_667_4_lut_4_lut (.A(n31949), .B(\mtime_out[0] ), 
         .C(n31913), .D(cy), .Z(n31872)) /* synthesis lut_function=(A (B (D))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i4846_2_lut_rep_667_4_lut_4_lut.init = 16'hc840;
    LUT4 i4781_2_lut_4_lut_4_lut (.A(n31949), .B(instrret_count[0]), .C(instr_retired), 
         .D(cy_c), .Z(increment_result_3__N_1925[0])) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i4781_2_lut_4_lut_4_lut.init = 16'h369c;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n31949), .B(cmp), .C(alu_b_in[1]), .D(alu_a_in[1]), 
         .Z(n27558)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(166[50:62])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd00d;
    LUT4 i4729_2_lut_rep_582_3_lut_4_lut (.A(cy_adj_3108), .B(n31959), .C(n31949), 
         .D(alu_b_in[0]), .Z(n31787)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A ((C+(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(111[18:70])
    defparam i4729_2_lut_rep_582_3_lut_4_lut.init = 16'h208c;
    LUT4 i1_2_lut_3_lut_4_lut_adj_363 (.A(cy_adj_3108), .B(n31959), .C(n31949), 
         .D(alu_b_in[0]), .Z(n28436)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(111[18:70])
    defparam i1_2_lut_3_lut_4_lut_adj_363.init = 16'h9f60;
    LUT4 tmp_data_31__I_0_542_i24_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[23]), 
         .D(tmp_data[27]), .Z(\addr_out[23] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i1_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[0]), 
         .D(tmp_data[4]), .Z(\addr_out[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i2_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[1]), 
         .D(tmp_data[5]), .Z(\addr_out[1] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i3_3_lut_rep_693_4_lut (.A(n32014), .B(n26175), 
         .C(mepc[2]), .D(tmp_data[6]), .Z(n31898)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i3_3_lut_rep_693_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i23_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[22]), 
         .D(tmp_data[26]), .Z(\addr_out[22] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i22_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[21]), 
         .D(tmp_data[25]), .Z(\addr_out[21] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i21_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[20]), 
         .D(tmp_data[24]), .Z(\addr_out[20] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i20_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[19]), 
         .D(tmp_data[23]), .Z(\addr_out[19] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i19_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[18]), 
         .D(tmp_data[22]), .Z(\addr_out[18] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i18_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[17]), 
         .D(tmp_data[21]), .Z(\addr_out[17] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i17_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[16]), 
         .D(tmp_data[20]), .Z(\addr_out[16] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i16_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[15]), 
         .D(tmp_data[19]), .Z(\addr_out[15] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i15_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[14]), 
         .D(tmp_data[18]), .Z(\addr_out[14] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i14_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[13]), 
         .D(tmp_data[17]), .Z(\addr_out[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i14_3_lut_4_lut.init = 16'hf780;
    PFUMX i26539 (.BLUT(csr_read_3__N_1447[0]), .ALUT(csr_read_3__N_1459[0]), 
          .C0(\imm[6] ), .Z(n29156));
    LUT4 tmp_data_31__I_0_542_i13_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[12]), 
         .D(tmp_data[16]), .Z(\addr_out[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i12_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[11]), 
         .D(tmp_data[15]), .Z(\addr_out[11] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i11_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[10]), 
         .D(tmp_data[14]), .Z(\addr_out[10] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i10_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[9]), 
         .D(tmp_data[13]), .Z(\addr_out[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i9_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[8]), 
         .D(tmp_data[12]), .Z(\addr_out[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i8_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[7]), 
         .D(tmp_data[11]), .Z(\addr_out[7] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i7_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[6]), 
         .D(tmp_data[10]), .Z(\addr_out[6] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i6_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[5]), 
         .D(tmp_data[9]), .Z(\addr_out[5] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 tmp_data_31__I_0_542_i5_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[4]), 
         .D(tmp_data[8]), .Z(\addr_out[4] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i5_3_lut_4_lut.init = 16'hf780;
    PFUMX i26536 (.BLUT(csr_read_3__N_1439[3]), .ALUT(csr_read_3__N_1455[3]), 
          .C0(\imm[1] ), .Z(n29153));
    LUT4 tmp_data_31__I_0_542_i4_3_lut_4_lut (.A(n32014), .B(n26175), .C(mepc[3]), 
         .D(tmp_data[7]), .Z(\addr_out[3] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam tmp_data_31__I_0_542_i4_3_lut_4_lut.init = 16'hf780;
    PFUMX i66 (.BLUT(n26149), .ALUT(n27180), .C0(\imm[11] ), .Z(n46));
    LUT4 mux_3121_i2_4_lut_4_lut (.A(n31946), .B(n31949), .C(mstatus_mpie), 
         .D(mstatus_mie), .Z(csr_read_3__N_1439[3])) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(471[33:47])
    defparam mux_3121_i2_4_lut_4_lut.init = 16'h7340;
    LUT4 i1_4_lut_adj_364 (.A(n28946), .B(n18), .C(\imm[0] ), .D(\imm[1] ), 
         .Z(n26019)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_364.init = 16'hfffe;
    LUT4 i26388_4_lut (.A(n28664), .B(\imm[4] ), .C(\imm[9] ), .D(n31983), 
         .Z(n28946)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i26388_4_lut.init = 16'hefff;
    LUT4 i1_2_lut_adj_365 (.A(\imm[10] ), .B(\imm[11] ), .Z(n28664)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(496[13:20])
    defparam i1_2_lut_adj_365.init = 16'heeee;
    LUT4 imm_lo_11__I_0_534_i18_2_lut (.A(\imm[7] ), .B(\imm[8] ), .Z(n18)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(487[13:20])
    defparam imm_lo_11__I_0_534_i18_2_lut.init = 16'hbbbb;
    LUT4 i13246_3_lut_4_lut (.A(n32044), .B(n26175), .C(n15837), .D(interrupt_core), 
         .Z(n611[1])) /* synthesis lut_function=(A (C (D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i13246_3_lut_4_lut.init = 16'hf044;
    LUT4 i1_4_lut_4_lut_4_lut_rep_864 (.A(n31744), .B(n31738), .C(n27960), 
         .D(n31742), .Z(n33493)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(462[32:59])
    defparam i1_4_lut_4_lut_4_lut_rep_864.init = 16'h0040;
    LUT4 i8931_2_lut_3_lut_4_lut (.A(n32044), .B(n26175), .C(clk_c_enable_544), 
         .D(interrupt_core), .Z(n11557)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i8931_2_lut_3_lut_4_lut.init = 16'hf040;
    PFUMX i28596 (.BLUT(n31689), .ALUT(n31688), .C0(\imm[10] ), .Z(n31690));
    LUT4 i27918_2_lut_3_lut_4_lut (.A(n32044), .B(n26175), .C(n5737), 
         .D(interrupt_core), .Z(n29351)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i27918_2_lut_3_lut_4_lut.init = 16'hfff4;
    PFUMX instr_complete_I_133 (.BLUT(instr_complete_N_1651), .ALUT(instr_complete_N_1652), 
          .C0(debug_rd_3__N_1401), .Z(instr_complete_N_1650)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=72, LSE_RCOL=6, LSE_LLINE=322, LSE_RLINE=368 */ ;
    LUT4 tmp_data_in_3__N_1581_I_0_588_2_lut_rep_673_3_lut_4_lut (.A(n32044), 
         .B(n26175), .C(n31949), .D(interrupt_core), .Z(n31878)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C)+!B (C+!(D))))) */ ;
    defparam tmp_data_in_3__N_1581_I_0_588_2_lut_rep_673_3_lut_4_lut.init = 16'h0f04;
    PFUMX mux_3524_i3 (.BLUT(time_count[2]), .ALUT(n5661), .C0(n29539), 
          .Z(n5671[2]));
    LUT4 i1_4_lut_adj_366 (.A(stall_core), .B(clk_c_enable_36), .C(n32046), 
         .D(\addr_offset[2] ), .Z(n28282)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_4_lut_adj_366.init = 16'h8000;
    LUT4 i1_3_lut_rep_538_4_lut (.A(clk_c_enable_36), .B(n32046), .C(instr_complete_N_1647), 
         .D(stall_core), .Z(n31743)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_rep_538_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_adj_367 (.A(clk_c_enable_36), .B(n32046), .C(stall_core), 
         .D(\next_pc_offset[3] ), .Z(n27604)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(217[9] 229[12])
    defparam i1_3_lut_4_lut_adj_367.init = 16'h2000;
    LUT4 i1_4_lut_adj_368 (.A(n31888), .B(instr_complete_N_1648), .C(n18009), 
         .D(n10873), .Z(n18086)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(220[18] 228[36])
    defparam i1_4_lut_adj_368.init = 16'hffef;
    LUT4 i15442_2_lut (.A(cycle[0]), .B(cycle[1]), .Z(n18009)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15442_2_lut.init = 16'h8888;
    PFUMX i26537 (.BLUT(time_count[3]), .ALUT(n5624[3]), .C0(n32011), 
          .Z(n29154));
    L6MUX21 i28739 (.D0(n32330), .D1(n32328), .SD(n29330), .Z(debug_rd_3__N_1567[3]));
    PFUMX i28737 (.BLUT(n32329), .ALUT(\debug_branch_N_446[31] ), .C0(n29333), 
          .Z(n32330));
    LUT4 i1_3_lut_4_lut_3_lut_4_lut_4_lut (.A(n31987), .B(\alu_op[0] ), 
         .C(\alu_op[1] ), .D(data_rs1_c[1]), .Z(n14)) /* synthesis lut_function=(!((B ((D)+!C)+!B !(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(75[19:52])
    defparam i1_3_lut_4_lut_3_lut_4_lut_4_lut.init = 16'h20a0;
    PFUMX i28735 (.BLUT(n32327), .ALUT(n32326), .C0(counter_hi[4]), .Z(n32328));
    PFUMX i26540 (.BLUT(\csr_read_3__N_1443[0] ), .ALUT(csr_read_3__N_1451[0]), 
          .C0(\imm[6] ), .Z(n29157));
    PFUMX i28634 (.BLUT(n32097), .ALUT(n32098), .C0(counter_hi[2]), .Z(\csr_read_3__N_1447[2] ));
    PFUMX i28632 (.BLUT(n32093), .ALUT(n32094), .C0(counter_hi[2]), .Z(n32095));
    LUT4 imm_10__bdd_3_lut_28595_3_lut_4_lut (.A(n31988), .B(counter_hi[2]), 
         .C(instrret_count[1]), .D(\imm[0] ), .Z(n31688)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(150[15:31])
    defparam imm_10__bdd_3_lut_28595_3_lut_4_lut.init = 16'h11f0;
    PFUMX i28535 (.BLUT(n31587), .ALUT(n31586), .C0(\imm[0] ), .Z(n31588));
    tinyqv_mul multiplier (.accum({accum}), .clk_c(clk_c), .mul_out_3__N_1510({mul_out_3__N_1510}), 
            .\tmp_data[0] (tmp_data[0]), .\tmp_data[1] (tmp_data[1]), .\tmp_data[2] (tmp_data[2]), 
            .\tmp_data[3] (tmp_data[3]), .\tmp_data[4] (tmp_data[4]), .\tmp_data[5] (tmp_data[5]), 
            .\tmp_data[6] (tmp_data[6]), .\tmp_data[7] (tmp_data[7]), .\tmp_data[8] (tmp_data[8]), 
            .\tmp_data[9] (tmp_data[9]), .\tmp_data[10] (tmp_data[10]), 
            .\tmp_data[11] (tmp_data[11]), .\tmp_data[12] (tmp_data[12]), 
            .\tmp_data[13] (tmp_data[13]), .\tmp_data[14] (tmp_data[14]), 
            .\tmp_data[15] (tmp_data[15]), .d_3__N_1868({d_3__N_1868}), 
            .GND_net(GND_net), .VCC_net(VCC_net), .\next_accum[5] (\next_accum[5] ), 
            .\next_accum[6] (\next_accum[6] ), .\next_accum[7] (\next_accum[7] ), 
            .\next_accum[8] (\next_accum[8] ), .\next_accum[9] (\next_accum[9] ), 
            .\next_accum[10] (\next_accum[10] ), .\next_accum[11] (\next_accum[11] ), 
            .\next_accum[12] (\next_accum[12] ), .\next_accum[13] (\next_accum[13] ), 
            .\next_accum[14] (\next_accum[14] ), .\next_accum[15] (\next_accum[15] ), 
            .\next_accum[16] (\next_accum[16] ), .\next_accum[17] (\next_accum[17] ), 
            .\next_accum[18] (\next_accum[18] ), .\next_accum[19] (\next_accum[19] ), 
            .\next_accum[4] (\next_accum[4] ), .\cycle[0] (cycle[0]), .data_rs1({data_rs1_c[3:1], 
            data_rs1[0]})) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(139[31:97])
    tinyqv_shifter i_shift (.\shift_amt[1] (shift_amt[1]), .\shift_amt[0] (shift_amt[0]), 
            .\shift_amt[2] (shift_amt_adj_3116[2]), .\shift_amt[3] (shift_amt_adj_3116[3]), 
            .tmp_data({tmp_data}), .\alu_op_in[2] (\alu_op_in[2] ), .n33486(n33486), 
            .\alu_op[3] (\alu_op[3] ), .shift_out({shift_out}), .\counter_hi[2] (counter_hi[2]), 
            .n33484(n33484), .\shift_amt[4] (shift_amt_adj_3116[4]), .\counter_hi[4] (counter_hi[4])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(133[20:81])
    tinyqv_registers i_registers (.rd({rd}), .debug_reg_wen(debug_reg_wen), 
            .rs2({rs2}), .n12(n12_adj_2), .n11(n11), .n9(n9), .n8(n8), 
            .rs1({rs1}), .clk_c(clk_c), .return_addr({return_addr}), .\registers[5][7] (\registers[5][7] ), 
            .\registers[6][7] (\registers[6][7] ), .\registers[7][7] (\registers[7][7] ), 
            .debug_rd({debug_rd}), .counter_hi({counter_hi}), .clk_c_enable_543(clk_c_enable_543), 
            .mstatus_mie(mstatus_mie), .interrupt_pending_N_1671(interrupt_pending_N_1671), 
            .n27480(n27480), .was_early_branch(was_early_branch), .n26597(n26597), 
            .n31747(n31747), .rst_reg_n(rst_reg_n), .n18086(n18086), .clk_c_enable_348(clk_c_enable_348), 
            .no_write_in_progress(no_write_in_progress), .n27534(n27534), 
            .time_hi({time_hi}), .\cycle_count_wide[6] (cycle_count_wide[6]), 
            .\time_count[3] (time_count[3]), .\cycle_count_wide[4] (cycle_count_wide[4]), 
            .\time_count[1] (time_count[1]), .n28150(n28150), .n27762(n27762), 
            .\cycle_count_wide[5] (cycle_count_wide[5]), .\time_count[2] (time_count[2]), 
            .n27018(n27018), .n28182(n28182), .n15604(n15604), .n29747(n29747), 
            .\data_rs2[1] (\data_rs2[1] ), .n4(n4), .\reg_access[3][2] (\reg_access[3][2] ), 
            .n33484(n33484), .\mcause[5] (mcause[5]), .n28520(n28520), 
            .n30165(n30165), .n30166(n30166), .n30169(n30169), .n33486(n33486), 
            .n31748(n31748), .n32046(n32046), .n31917(n31917), .n30167(n30167), 
            .n31943(n31943), .clk_c_enable_36(clk_c_enable_36), .\mepc[0] (mepc[0]), 
            .\csr_read_3__N_1451[0] (csr_read_3__N_1451[0]), .n30168(n30168), 
            .n11559(n11559), .\imm[6] (\imm[6] ), .n26121(n26121), .\mepc[3] (mepc[3]), 
            .n31171(n31171), .data_rs1({data_rs1_c[3:1], data_rs1[0]}), 
            .\data_rs2[0] (\data_rs2[0] ), .\data_rs2[2] (\data_rs2[2] ), 
            .n33494(n33494)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(91[9:103])
    tinyqv_counter_U0 i_instrret (.cy(cy_c), .clk_c(clk_c), .n31980(n31980), 
            .\increment_result_3__N_1925[0] (increment_result_3__N_1925[0]), 
            .instrret_count({instrret_count}), .n31873(n31873), .n31890(n31890)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(307[20] 315[6])
    \tinyqv_counter(OUTPUT_WIDTH=7)  i_cycles (.cy(cy_adj_3109), .clk_c(clk_c), 
            .n31980(n31980), .\increment_result_3__N_1911[0] (increment_result_3__N_1911[0]), 
            .cycle_count_wide({cycle_count_wide[6:4], \cycle_count_wide[3] , 
            cycle_count_wide[2:0]}), .n31912(n31912), .n31945(n31945), 
            .n31870(n31870), .n31949(n31949)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(281[40] 290[6])
    tinyqv_alu i_alu (.alu_a_in({alu_a_in}), .n31826(n31826), .n31827(n31827), 
            .n30868(n30868), .n28436(n28436), .alu_b_in({\alu_b_in[3] , 
            alu_b_in[2:0]}), .\alu_op_in[2] (\alu_op_in[2] ), .n31959(n31959), 
            .n31924(n31924), .n31787(n31787), .n31856(n31856), .cy_out(cy_out), 
            .n27558(n27558), .n4913({n4913}), .n31979(n31979), .n30870(n30870), 
            .n31825(n31825), .n31960(n31960), .alu_out({alu_out})) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/core.v(115[16:93])
    
endmodule
//
// Verilog Description of module tinyqv_mul
//

module tinyqv_mul (accum, clk_c, mul_out_3__N_1510, \tmp_data[0] , \tmp_data[1] , 
            \tmp_data[2] , \tmp_data[3] , \tmp_data[4] , \tmp_data[5] , 
            \tmp_data[6] , \tmp_data[7] , \tmp_data[8] , \tmp_data[9] , 
            \tmp_data[10] , \tmp_data[11] , \tmp_data[12] , \tmp_data[13] , 
            \tmp_data[14] , \tmp_data[15] , d_3__N_1868, GND_net, VCC_net, 
            \next_accum[5] , \next_accum[6] , \next_accum[7] , \next_accum[8] , 
            \next_accum[9] , \next_accum[10] , \next_accum[11] , \next_accum[12] , 
            \next_accum[13] , \next_accum[14] , \next_accum[15] , \next_accum[16] , 
            \next_accum[17] , \next_accum[18] , \next_accum[19] , \next_accum[4] , 
            \cycle[0] , data_rs1) /* synthesis syn_module_defined=1 */ ;
    output [15:0]accum;
    input clk_c;
    input [3:0]mul_out_3__N_1510;
    input \tmp_data[0] ;
    input \tmp_data[1] ;
    input \tmp_data[2] ;
    input \tmp_data[3] ;
    input \tmp_data[4] ;
    input \tmp_data[5] ;
    input \tmp_data[6] ;
    input \tmp_data[7] ;
    input \tmp_data[8] ;
    input \tmp_data[9] ;
    input \tmp_data[10] ;
    input \tmp_data[11] ;
    input \tmp_data[12] ;
    input \tmp_data[13] ;
    input \tmp_data[14] ;
    input \tmp_data[15] ;
    output [19:0]d_3__N_1868;
    input GND_net;
    input VCC_net;
    input \next_accum[5] ;
    input \next_accum[6] ;
    input \next_accum[7] ;
    input \next_accum[8] ;
    input \next_accum[9] ;
    input \next_accum[10] ;
    input \next_accum[11] ;
    input \next_accum[12] ;
    input \next_accum[13] ;
    input \next_accum[14] ;
    input \next_accum[15] ;
    input \next_accum[16] ;
    input \next_accum[17] ;
    input \next_accum[18] ;
    input \next_accum[19] ;
    input \next_accum[4] ;
    input \cycle[0] ;
    input [3:0]data_rs1;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [15:0]accum_15__N_1888;
    
    wire n7, n28638;
    
    FD1S3AX accum_i0 (.D(accum_15__N_1888[0]), .CK(clk_c), .Q(accum[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i0.GSR = "DISABLED";
    MULT18X18D a_3__I_0_11_mult_2 (.A17(GND_net), .A16(GND_net), .A15(GND_net), 
            .A14(GND_net), .A13(GND_net), .A12(GND_net), .A11(GND_net), 
            .A10(GND_net), .A9(GND_net), .A8(GND_net), .A7(GND_net), 
            .A6(GND_net), .A5(GND_net), .A4(GND_net), .A3(mul_out_3__N_1510[3]), 
            .A2(mul_out_3__N_1510[2]), .A1(mul_out_3__N_1510[1]), .A0(mul_out_3__N_1510[0]), 
            .B17(GND_net), .B16(GND_net), .B15(\tmp_data[15] ), .B14(\tmp_data[14] ), 
            .B13(\tmp_data[13] ), .B12(\tmp_data[12] ), .B11(\tmp_data[11] ), 
            .B10(\tmp_data[10] ), .B9(\tmp_data[9] ), .B8(\tmp_data[8] ), 
            .B7(\tmp_data[7] ), .B6(\tmp_data[6] ), .B5(\tmp_data[5] ), 
            .B4(\tmp_data[4] ), .B3(\tmp_data[3] ), .B2(\tmp_data[2] ), 
            .B1(\tmp_data[1] ), .B0(\tmp_data[0] ), .C17(GND_net), .C16(GND_net), 
            .C15(GND_net), .C14(GND_net), .C13(GND_net), .C12(GND_net), 
            .C11(GND_net), .C10(GND_net), .C9(GND_net), .C8(GND_net), 
            .C7(GND_net), .C6(GND_net), .C5(GND_net), .C4(GND_net), 
            .C3(GND_net), .C2(GND_net), .C1(GND_net), .C0(GND_net), 
            .SIGNEDA(GND_net), .SIGNEDB(GND_net), .SOURCEA(GND_net), .SOURCEB(GND_net), 
            .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), .CLK0(GND_net), 
            .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), .CE0(VCC_net), 
            .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), .RST0(GND_net), 
            .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), .SRIA14(GND_net), 
            .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), .SRIA10(GND_net), 
            .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), .SRIA6(GND_net), 
            .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), .SRIA2(GND_net), 
            .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), .SRIB16(GND_net), 
            .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), .SRIB12(GND_net), 
            .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), .SRIB8(GND_net), 
            .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), .SRIB4(GND_net), 
            .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), .SRIB0(GND_net), 
            .P19(d_3__N_1868[19]), .P18(d_3__N_1868[18]), .P17(d_3__N_1868[17]), 
            .P16(d_3__N_1868[16]), .P15(d_3__N_1868[15]), .P14(d_3__N_1868[14]), 
            .P13(d_3__N_1868[13]), .P12(d_3__N_1868[12]), .P11(d_3__N_1868[11]), 
            .P10(d_3__N_1868[10]), .P9(d_3__N_1868[9]), .P8(d_3__N_1868[8]), 
            .P7(d_3__N_1868[7]), .P6(d_3__N_1868[6]), .P5(d_3__N_1868[5]), 
            .P4(d_3__N_1868[4]), .P3(d_3__N_1868[3]), .P2(d_3__N_1868[2]), 
            .P1(d_3__N_1868[1]), .P0(d_3__N_1868[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(105[52:83])
    defparam a_3__I_0_11_mult_2.REG_INPUTA_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTA_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTA_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTB_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_INPUTC_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_PIPELINE_RST = "RST0";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_CE = "CE0";
    defparam a_3__I_0_11_mult_2.REG_OUTPUT_RST = "RST0";
    defparam a_3__I_0_11_mult_2.CLK0_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK1_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK2_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.CLK3_DIV = "ENABLED";
    defparam a_3__I_0_11_mult_2.HIGHSPEED_CLK = "NONE";
    defparam a_3__I_0_11_mult_2.GSR = "DISABLED";
    defparam a_3__I_0_11_mult_2.CAS_MATCH_REG = "FALSE";
    defparam a_3__I_0_11_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam a_3__I_0_11_mult_2.MULT_BYPASS = "DISABLED";
    defparam a_3__I_0_11_mult_2.RESETMODE = "SYNC";
    LUT4 accum_15__I_0_i2_3_lut (.A(accum[5]), .B(\next_accum[5] ), .C(n7), 
         .Z(accum_15__N_1888[1])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i2_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i3_3_lut (.A(accum[6]), .B(\next_accum[6] ), .C(n7), 
         .Z(accum_15__N_1888[2])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i3_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i4_3_lut (.A(accum[7]), .B(\next_accum[7] ), .C(n7), 
         .Z(accum_15__N_1888[3])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i4_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i5_3_lut (.A(accum[8]), .B(\next_accum[8] ), .C(n7), 
         .Z(accum_15__N_1888[4])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i5_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i6_3_lut (.A(accum[9]), .B(\next_accum[9] ), .C(n7), 
         .Z(accum_15__N_1888[5])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i6_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i7_3_lut (.A(accum[10]), .B(\next_accum[10] ), .C(n7), 
         .Z(accum_15__N_1888[6])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i7_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i8_3_lut (.A(accum[11]), .B(\next_accum[11] ), .C(n7), 
         .Z(accum_15__N_1888[7])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i8_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i9_3_lut (.A(accum[12]), .B(\next_accum[12] ), .C(n7), 
         .Z(accum_15__N_1888[8])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i9_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i10_3_lut (.A(accum[13]), .B(\next_accum[13] ), .C(n7), 
         .Z(accum_15__N_1888[9])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i10_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i11_3_lut (.A(accum[14]), .B(\next_accum[14] ), .C(n7), 
         .Z(accum_15__N_1888[10])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i11_3_lut.init = 16'hacac;
    LUT4 accum_15__I_0_i12_3_lut (.A(accum[15]), .B(\next_accum[15] ), .C(n7), 
         .Z(accum_15__N_1888[11])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i12_3_lut.init = 16'hacac;
    FD1S3IX accum_i12 (.D(\next_accum[16] ), .CK(clk_c), .CD(n7), .Q(accum[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i12.GSR = "DISABLED";
    FD1S3AX accum_i1 (.D(accum_15__N_1888[1]), .CK(clk_c), .Q(accum[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i1.GSR = "DISABLED";
    FD1S3AX accum_i2 (.D(accum_15__N_1888[2]), .CK(clk_c), .Q(accum[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i2.GSR = "DISABLED";
    FD1S3AX accum_i3 (.D(accum_15__N_1888[3]), .CK(clk_c), .Q(accum[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i3.GSR = "DISABLED";
    FD1S3AX accum_i4 (.D(accum_15__N_1888[4]), .CK(clk_c), .Q(accum[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i4.GSR = "DISABLED";
    FD1S3AX accum_i5 (.D(accum_15__N_1888[5]), .CK(clk_c), .Q(accum[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i5.GSR = "DISABLED";
    FD1S3AX accum_i6 (.D(accum_15__N_1888[6]), .CK(clk_c), .Q(accum[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i6.GSR = "DISABLED";
    FD1S3AX accum_i7 (.D(accum_15__N_1888[7]), .CK(clk_c), .Q(accum[7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i7.GSR = "DISABLED";
    FD1S3AX accum_i8 (.D(accum_15__N_1888[8]), .CK(clk_c), .Q(accum[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i8.GSR = "DISABLED";
    FD1S3AX accum_i9 (.D(accum_15__N_1888[9]), .CK(clk_c), .Q(accum[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i9.GSR = "DISABLED";
    FD1S3AX accum_i10 (.D(accum_15__N_1888[10]), .CK(clk_c), .Q(accum[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i10.GSR = "DISABLED";
    FD1S3AX accum_i11 (.D(accum_15__N_1888[11]), .CK(clk_c), .Q(accum[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i11.GSR = "DISABLED";
    FD1S3IX accum_i13 (.D(\next_accum[17] ), .CK(clk_c), .CD(n7), .Q(accum[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i13.GSR = "DISABLED";
    FD1S3IX accum_i14 (.D(\next_accum[18] ), .CK(clk_c), .CD(n7), .Q(accum[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i14.GSR = "DISABLED";
    FD1S3IX accum_i15 (.D(\next_accum[19] ), .CK(clk_c), .CD(n7), .Q(accum[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=31, LSE_RCOL=97, LSE_LLINE=139, LSE_RLINE=139 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(107[12] 109[8])
    defparam accum_i15.GSR = "DISABLED";
    LUT4 accum_15__I_0_i1_3_lut (.A(accum[4]), .B(\next_accum[4] ), .C(n7), 
         .Z(accum_15__N_1888[0])) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:88])
    defparam accum_15__I_0_i1_3_lut.init = 16'hacac;
    LUT4 i27829_4_lut (.A(\cycle[0] ), .B(n28638), .C(data_rs1[3]), .D(data_rs1[0]), 
         .Z(n7)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:32])
    defparam i27829_4_lut.init = 16'h5557;
    LUT4 i1_2_lut (.A(data_rs1[2]), .B(data_rs1[1]), .Z(n28638)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(108[18:32])
    defparam i1_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module tinyqv_shifter
//

module tinyqv_shifter (\shift_amt[1] , \shift_amt[0] , \shift_amt[2] , 
            \shift_amt[3] , tmp_data, \alu_op_in[2] , n33486, \alu_op[3] , 
            shift_out, \counter_hi[2] , n33484, \shift_amt[4] , \counter_hi[4] ) /* synthesis syn_module_defined=1 */ ;
    input \shift_amt[1] ;
    input \shift_amt[0] ;
    input \shift_amt[2] ;
    input \shift_amt[3] ;
    input [31:0]tmp_data;
    input \alu_op_in[2] ;
    input n33486;
    input \alu_op[3] ;
    output [3:0]shift_out;
    input \counter_hi[2] ;
    input n33484;
    input \shift_amt[4] ;
    input \counter_hi[4] ;
    
    
    wire n117, n121, n30162, n29698, n29583, n29584;
    wire [5:0]shift_amt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[16:25])
    
    wire n29589, n47, n49, n113, n43, n45, n109, n36, n38, 
        n29580, n32, n34, n29579;
    wire [31:0]a_for_shift_right;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[17:34])
    
    wire n31998, n129, n46, n29585, n29586, n29590, n58, n60, 
        n29687, n32032, n29844, n4, n54, n56, n29686, n50, n52, 
        n29685, n48, n29684, n42, n44, n29683, n29601, n29602, 
        n30164, n29609, n40, n29682, n29603, n29604, n29610, n125, 
        n29699, n29681;
    wire [65:0]dr_3__N_1864;
    
    wire n9417, n29605, n29606, n30163, n29611, n9415, n9413, 
        n8720, n63, n62, n29688, n51, n53, n55, n57, n59, 
        n61, n29607, n29608, n29612, n39, n41, n105, n35, n37, 
        n101, n29696, n29689, n33, n29690, n29691, n29591, n29592, 
        n29613, n29614, n29693, n29694, n29700, n29701, n29692, 
        n29697, n29587, n29588, n29582, n29581;
    
    PFUMX i27081 (.BLUT(n117), .ALUT(n121), .C0(n30162), .Z(n29698));
    PFUMX i26972 (.BLUT(n29583), .ALUT(n29584), .C0(shift_amt[2]), .Z(n29589));
    LUT4 top_bit_I_0_i113_3_lut (.A(n47), .B(n49), .C(\shift_amt[1] ), 
         .Z(n113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i113_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i109_3_lut (.A(n43), .B(n45), .C(\shift_amt[1] ), 
         .Z(n109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i109_3_lut.init = 16'hcaca;
    LUT4 i26963_3_lut (.A(n36), .B(n38), .C(\shift_amt[1] ), .Z(n29580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26963_3_lut.init = 16'hcaca;
    LUT4 i26962_3_lut (.A(n32), .B(n34), .C(\shift_amt[1] ), .Z(n29579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26962_3_lut.init = 16'hcaca;
    LUT4 i6222_4_lut (.A(a_for_shift_right[31]), .B(n31998), .C(\shift_amt[0] ), 
         .D(\shift_amt[1] ), .Z(n129)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam i6222_4_lut.init = 16'hccca;
    LUT4 top_bit_I_0_i46_3_lut (.A(a_for_shift_right[14]), .B(a_for_shift_right[15]), 
         .C(\shift_amt[0] ), .Z(n46)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i46_3_lut.init = 16'hcaca;
    PFUMX i26973 (.BLUT(n29585), .ALUT(n29586), .C0(shift_amt[2]), .Z(n29590));
    LUT4 i27070_3_lut (.A(n58), .B(n60), .C(\shift_amt[1] ), .Z(n29687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27070_3_lut.init = 16'hcaca;
    LUT4 i4717_3_lut_4_lut (.A(\shift_amt[2] ), .B(n32032), .C(n29844), 
         .D(\shift_amt[3] ), .Z(n4)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[28:55])
    defparam i4717_3_lut_4_lut.init = 16'h2f02;
    LUT4 i2_3_lut_4_lut (.A(\shift_amt[2] ), .B(n32032), .C(n29844), .D(\shift_amt[3] ), 
         .Z(shift_amt[3])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(80[28:55])
    defparam i2_3_lut_4_lut.init = 16'hd22d;
    LUT4 i27069_3_lut (.A(n54), .B(n56), .C(\shift_amt[1] ), .Z(n29686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27069_3_lut.init = 16'hcaca;
    LUT4 i27068_3_lut (.A(n50), .B(n52), .C(\shift_amt[1] ), .Z(n29685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27068_3_lut.init = 16'hcaca;
    LUT4 i27067_3_lut (.A(n46), .B(n48), .C(\shift_amt[1] ), .Z(n29684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27067_3_lut.init = 16'hcaca;
    LUT4 i27066_3_lut (.A(n42), .B(n44), .C(\shift_amt[1] ), .Z(n29683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27066_3_lut.init = 16'hcaca;
    PFUMX i26992 (.BLUT(n29601), .ALUT(n29602), .C0(n30164), .Z(n29609));
    LUT4 i27065_3_lut (.A(n38), .B(n40), .C(\shift_amt[1] ), .Z(n29682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27065_3_lut.init = 16'hcaca;
    PFUMX i26993 (.BLUT(n29603), .ALUT(n29604), .C0(n30164), .Z(n29610));
    PFUMX i27082 (.BLUT(n125), .ALUT(n129), .C0(n30162), .Z(n29699));
    LUT4 i27064_3_lut (.A(n34), .B(n36), .C(\shift_amt[1] ), .Z(n29681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27064_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i45_3_lut (.A(a_for_shift_right[13]), .B(a_for_shift_right[14]), 
         .C(\shift_amt[0] ), .Z(n45)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i45_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i47_4_lut (.A(tmp_data[16]), .B(tmp_data[15]), .C(\alu_op_in[2] ), 
         .D(\shift_amt[0] ), .Z(n47)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A !((C (D)+!C !(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i47_4_lut.init = 16'hacca;
    LUT4 i6817_3_lut (.A(dr_3__N_1864[31]), .B(dr_3__N_1864[34]), .C(\alu_op_in[2] ), 
         .Z(n9417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i6817_3_lut.init = 16'hcaca;
    LUT4 i27632_2_lut (.A(n33486), .B(\alu_op_in[2] ), .Z(n29844)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i27632_2_lut.init = 16'h6666;
    PFUMX i26994 (.BLUT(n29605), .ALUT(n29606), .C0(n30163), .Z(n29611));
    LUT4 i6815_3_lut (.A(dr_3__N_1864[32]), .B(dr_3__N_1864[33]), .C(\alu_op_in[2] ), 
         .Z(n9415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i6815_3_lut.init = 16'hcaca;
    LUT4 i6813_3_lut (.A(dr_3__N_1864[33]), .B(dr_3__N_1864[32]), .C(\alu_op_in[2] ), 
         .Z(n9413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i6813_3_lut.init = 16'hcaca;
    LUT4 i15511_2_lut_rep_793 (.A(tmp_data[31]), .B(\alu_op[3] ), .Z(n31998)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i15511_2_lut_rep_793.init = 16'h8888;
    LUT4 i6818_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n9417), .Z(shift_out[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i6818_3_lut_4_lut.init = 16'h8f80;
    LUT4 i6129_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n8720), .Z(shift_out[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i6129_3_lut_4_lut.init = 16'h8f80;
    LUT4 i6814_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n9413), .Z(shift_out[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i6814_3_lut_4_lut.init = 16'h8f80;
    LUT4 top_bit_I_0_i63_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), 
         .C(\shift_amt[0] ), .D(a_for_shift_right[31]), .Z(n63)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam top_bit_I_0_i63_3_lut_4_lut.init = 16'h8f80;
    LUT4 i27071_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(\shift_amt[1] ), 
         .D(n62), .Z(n29688)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i27071_3_lut_4_lut.init = 16'h8f80;
    LUT4 i6816_3_lut_4_lut (.A(tmp_data[31]), .B(\alu_op[3] ), .C(shift_amt[5]), 
         .D(n9415), .Z(shift_out[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(69[20:40])
    defparam i6816_3_lut_4_lut.init = 16'h8f80;
    LUT4 top_bit_I_0_i51_3_lut (.A(a_for_shift_right[19]), .B(a_for_shift_right[20]), 
         .C(\shift_amt[0] ), .Z(n51)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i51_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i53_3_lut (.A(a_for_shift_right[21]), .B(a_for_shift_right[22]), 
         .C(\shift_amt[0] ), .Z(n53)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i53_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i22_3_lut (.A(tmp_data[10]), .B(tmp_data[21]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i23_3_lut (.A(tmp_data[9]), .B(tmp_data[22]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i20_3_lut (.A(tmp_data[12]), .B(tmp_data[19]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i21_3_lut (.A(tmp_data[11]), .B(tmp_data[20]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i55_3_lut (.A(a_for_shift_right[23]), .B(a_for_shift_right[24]), 
         .C(\shift_amt[0] ), .Z(n55)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i55_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i57_3_lut (.A(a_for_shift_right[25]), .B(a_for_shift_right[26]), 
         .C(\shift_amt[0] ), .Z(n57)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i57_3_lut.init = 16'hcaca;
    LUT4 i6128_3_lut (.A(dr_3__N_1864[34]), .B(dr_3__N_1864[31]), .C(\alu_op_in[2] ), 
         .Z(n8720)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(91[16:68])
    defparam i6128_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i26_3_lut (.A(tmp_data[6]), .B(tmp_data[25]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i27_3_lut (.A(tmp_data[5]), .B(tmp_data[26]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i24_3_lut (.A(tmp_data[8]), .B(tmp_data[23]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i24_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i59_3_lut (.A(a_for_shift_right[27]), .B(a_for_shift_right[28]), 
         .C(\shift_amt[0] ), .Z(n59)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i59_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i61_3_lut (.A(a_for_shift_right[29]), .B(a_for_shift_right[30]), 
         .C(\shift_amt[0] ), .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i61_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i25_3_lut (.A(tmp_data[7]), .B(tmp_data[24]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i7_3_lut (.A(tmp_data[25]), .B(tmp_data[6]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i7_3_lut.init = 16'hcaca;
    PFUMX i26995 (.BLUT(n29607), .ALUT(n29608), .C0(n30163), .Z(n29612));
    LUT4 top_bit_I_0_i105_3_lut (.A(n39), .B(n41), .C(\shift_amt[1] ), 
         .Z(n105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i105_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i101_3_lut (.A(n35), .B(n37), .C(\shift_amt[1] ), 
         .Z(n101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i101_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i34_3_lut (.A(a_for_shift_right[2]), .B(a_for_shift_right[3]), 
         .C(\shift_amt[0] ), .Z(n34)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i34_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i36_3_lut (.A(a_for_shift_right[4]), .B(a_for_shift_right[5]), 
         .C(\shift_amt[0] ), .Z(n36)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i36_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i38_3_lut (.A(a_for_shift_right[6]), .B(a_for_shift_right[7]), 
         .C(\shift_amt[0] ), .Z(n38)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i38_3_lut.init = 16'hcaca;
    PFUMX i27079 (.BLUT(n101), .ALUT(n105), .C0(n30164), .Z(n29696));
    LUT4 i27630_2_lut_rep_827 (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .Z(n32032)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i27630_2_lut_rep_827.init = 16'h6666;
    LUT4 i4704_rep_123_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .C(\shift_amt[2] ), .Z(n30162)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4704_rep_123_2_lut_3_lut.init = 16'h6969;
    LUT4 i4704_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), .C(\shift_amt[2] ), 
         .Z(shift_amt[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4704_2_lut_3_lut.init = 16'h6969;
    LUT4 i4704_rep_125_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .C(\shift_amt[2] ), .Z(n30164)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4704_rep_125_2_lut_3_lut.init = 16'h6969;
    LUT4 i4704_rep_124_2_lut_3_lut (.A(\counter_hi[2] ), .B(\alu_op_in[2] ), 
         .C(\shift_amt[2] ), .Z(n30163)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4704_rep_124_2_lut_3_lut.init = 16'h6969;
    LUT4 i26991_3_lut (.A(n61), .B(n63), .C(\shift_amt[1] ), .Z(n29608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26991_3_lut.init = 16'hcaca;
    LUT4 i26990_3_lut (.A(n57), .B(n59), .C(\shift_amt[1] ), .Z(n29607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26990_3_lut.init = 16'hcaca;
    LUT4 i26989_3_lut (.A(n53), .B(n55), .C(\shift_amt[1] ), .Z(n29606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26989_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i16_3_lut (.A(tmp_data[16]), .B(tmp_data[15]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i16_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i125_3_lut (.A(n59), .B(n61), .C(\shift_amt[1] ), 
         .Z(n125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i125_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i15_3_lut (.A(tmp_data[17]), .B(tmp_data[14]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 i26988_3_lut (.A(n49), .B(n51), .C(\shift_amt[1] ), .Z(n29605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26988_3_lut.init = 16'hcaca;
    LUT4 i4724_3_lut_4_lut (.A(n33484), .B(\alu_op_in[2] ), .C(n4), .D(\shift_amt[4] ), 
         .Z(shift_amt[5])) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A (B (C (D))+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i4724_3_lut_4_lut.init = 16'hf990;
    LUT4 i2_3_lut_4_lut_adj_278 (.A(\counter_hi[4] ), .B(\alu_op_in[2] ), 
         .C(n4), .D(\shift_amt[4] ), .Z(shift_amt[4])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(79[20:52])
    defparam i2_3_lut_4_lut_adj_278.init = 16'h9669;
    LUT4 i26987_3_lut (.A(n45), .B(n47), .C(\shift_amt[1] ), .Z(n29604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26987_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i32_3_lut (.A(a_for_shift_right[0]), .B(a_for_shift_right[1]), 
         .C(\shift_amt[0] ), .Z(n32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i32_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i1_3_lut (.A(tmp_data[31]), .B(tmp_data[0]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 i26986_3_lut (.A(n41), .B(n43), .C(\shift_amt[1] ), .Z(n29603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26986_3_lut.init = 16'hcaca;
    PFUMX i27072 (.BLUT(n29681), .ALUT(n29682), .C0(n30164), .Z(n29689));
    LUT4 top_bit_I_0_i48_3_lut (.A(a_for_shift_right[16]), .B(a_for_shift_right[17]), 
         .C(\shift_amt[0] ), .Z(n48)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i48_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i17_3_lut (.A(tmp_data[15]), .B(tmp_data[16]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i17_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i50_3_lut (.A(a_for_shift_right[18]), .B(a_for_shift_right[19]), 
         .C(\shift_amt[0] ), .Z(n50)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i50_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i18_3_lut (.A(tmp_data[14]), .B(tmp_data[17]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i19_3_lut (.A(tmp_data[13]), .B(tmp_data[18]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i52_3_lut (.A(a_for_shift_right[20]), .B(a_for_shift_right[21]), 
         .C(\shift_amt[0] ), .Z(n52)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i52_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i54_3_lut (.A(a_for_shift_right[22]), .B(a_for_shift_right[23]), 
         .C(\shift_amt[0] ), .Z(n54)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i54_3_lut.init = 16'hcaca;
    LUT4 i26985_3_lut (.A(n37), .B(n39), .C(\shift_amt[1] ), .Z(n29602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26985_3_lut.init = 16'hcaca;
    LUT4 i26984_3_lut (.A(n33), .B(n35), .C(\shift_amt[1] ), .Z(n29601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26984_3_lut.init = 16'hcaca;
    LUT4 i26969_3_lut (.A(n60), .B(n62), .C(\shift_amt[1] ), .Z(n29586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26969_3_lut.init = 16'hcaca;
    LUT4 i26968_3_lut (.A(n56), .B(n58), .C(\shift_amt[1] ), .Z(n29585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26968_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i56_3_lut (.A(a_for_shift_right[24]), .B(a_for_shift_right[25]), 
         .C(\shift_amt[0] ), .Z(n56)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i56_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i58_3_lut (.A(a_for_shift_right[26]), .B(a_for_shift_right[27]), 
         .C(\shift_amt[0] ), .Z(n58)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i58_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i28_3_lut (.A(tmp_data[4]), .B(tmp_data[27]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i60_3_lut (.A(a_for_shift_right[28]), .B(a_for_shift_right[29]), 
         .C(\shift_amt[0] ), .Z(n60)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i60_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i62_3_lut (.A(a_for_shift_right[30]), .B(a_for_shift_right[31]), 
         .C(\shift_amt[0] ), .Z(n62)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i62_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i31_3_lut (.A(tmp_data[1]), .B(tmp_data[30]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i32_3_lut (.A(tmp_data[0]), .B(tmp_data[31]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i29_3_lut (.A(tmp_data[3]), .B(tmp_data[28]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i30_3_lut (.A(tmp_data[2]), .B(tmp_data[29]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i30_3_lut.init = 16'hcaca;
    PFUMX i27073 (.BLUT(n29683), .ALUT(n29684), .C0(n30163), .Z(n29690));
    LUT4 top_bit_I_0_i41_3_lut (.A(a_for_shift_right[9]), .B(a_for_shift_right[10]), 
         .C(\shift_amt[0] ), .Z(n41)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i41_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i12_3_lut (.A(tmp_data[20]), .B(tmp_data[11]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i12_3_lut.init = 16'hcaca;
    PFUMX i27074 (.BLUT(n29685), .ALUT(n29686), .C0(n30163), .Z(n29691));
    L6MUX21 i26976 (.D0(n29591), .D1(n29592), .SD(shift_amt[4]), .Z(dr_3__N_1864[31]));
    L6MUX21 i26998 (.D0(n29613), .D1(n29614), .SD(shift_amt[4]), .Z(dr_3__N_1864[32]));
    L6MUX21 i27078 (.D0(n29693), .D1(n29694), .SD(shift_amt[4]), .Z(dr_3__N_1864[33]));
    L6MUX21 i27085 (.D0(n29700), .D1(n29701), .SD(shift_amt[4]), .Z(dr_3__N_1864[34]));
    LUT4 a_0__I_0_i13_3_lut (.A(tmp_data[19]), .B(tmp_data[12]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i13_3_lut.init = 16'hcaca;
    PFUMX i27075 (.BLUT(n29687), .ALUT(n29688), .C0(n30162), .Z(n29692));
    LUT4 top_bit_I_0_i43_3_lut (.A(a_for_shift_right[11]), .B(a_for_shift_right[12]), 
         .C(\shift_amt[0] ), .Z(n43)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i43_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i44_3_lut (.A(a_for_shift_right[12]), .B(a_for_shift_right[13]), 
         .C(\shift_amt[0] ), .Z(n44)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i44_3_lut.init = 16'hcaca;
    LUT4 i26967_3_lut (.A(n52), .B(n54), .C(\shift_amt[1] ), .Z(n29584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26967_3_lut.init = 16'hcaca;
    LUT4 i26966_3_lut (.A(n48), .B(n50), .C(\shift_amt[1] ), .Z(n29583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26966_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i121_3_lut (.A(n55), .B(n57), .C(\shift_amt[1] ), 
         .Z(n121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i121_3_lut.init = 16'hcaca;
    PFUMX i27080 (.BLUT(n109), .ALUT(n113), .C0(n30162), .Z(n29697));
    L6MUX21 i26974 (.D0(n29587), .D1(n29588), .SD(shift_amt[3]), .Z(n29591));
    L6MUX21 i26975 (.D0(n29589), .D1(n29590), .SD(shift_amt[3]), .Z(n29592));
    L6MUX21 i26996 (.D0(n29609), .D1(n29610), .SD(shift_amt[3]), .Z(n29613));
    L6MUX21 i26997 (.D0(n29611), .D1(n29612), .SD(shift_amt[3]), .Z(n29614));
    LUT4 top_bit_I_0_i117_3_lut (.A(n51), .B(n53), .C(\shift_amt[1] ), 
         .Z(n117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i117_3_lut.init = 16'hcaca;
    L6MUX21 i27076 (.D0(n29689), .D1(n29690), .SD(shift_amt[3]), .Z(n29693));
    L6MUX21 i27077 (.D0(n29691), .D1(n29692), .SD(shift_amt[3]), .Z(n29694));
    L6MUX21 i27083 (.D0(n29696), .D1(n29697), .SD(shift_amt[3]), .Z(n29700));
    L6MUX21 i27084 (.D0(n29698), .D1(n29699), .SD(shift_amt[3]), .Z(n29701));
    LUT4 top_bit_I_0_i40_3_lut (.A(a_for_shift_right[8]), .B(a_for_shift_right[9]), 
         .C(\shift_amt[0] ), .Z(n40)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i40_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i42_3_lut (.A(a_for_shift_right[10]), .B(a_for_shift_right[11]), 
         .C(\shift_amt[0] ), .Z(n42)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i42_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i9_3_lut (.A(tmp_data[23]), .B(tmp_data[8]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i33_3_lut (.A(a_for_shift_right[1]), .B(a_for_shift_right[2]), 
         .C(\shift_amt[0] ), .Z(n33)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i33_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i35_3_lut (.A(a_for_shift_right[3]), .B(a_for_shift_right[4]), 
         .C(\shift_amt[0] ), .Z(n35)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i35_3_lut.init = 16'hcaca;
    LUT4 i26965_3_lut (.A(n44), .B(n46), .C(\shift_amt[1] ), .Z(n29582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26965_3_lut.init = 16'hcaca;
    LUT4 i26964_3_lut (.A(n40), .B(n42), .C(\shift_amt[1] ), .Z(n29581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26964_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i2_3_lut (.A(tmp_data[30]), .B(tmp_data[1]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i49_3_lut (.A(a_for_shift_right[17]), .B(a_for_shift_right[18]), 
         .C(\shift_amt[0] ), .Z(n49)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i49_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i3_3_lut (.A(tmp_data[29]), .B(tmp_data[2]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i10_3_lut (.A(tmp_data[22]), .B(tmp_data[9]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i4_3_lut (.A(tmp_data[28]), .B(tmp_data[3]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i4_3_lut.init = 16'hcaca;
    PFUMX i26970 (.BLUT(n29579), .ALUT(n29580), .C0(shift_amt[2]), .Z(n29587));
    PFUMX i26971 (.BLUT(n29581), .ALUT(n29582), .C0(shift_amt[2]), .Z(n29588));
    LUT4 a_0__I_0_i5_3_lut (.A(tmp_data[27]), .B(tmp_data[4]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i37_3_lut (.A(a_for_shift_right[5]), .B(a_for_shift_right[6]), 
         .C(\shift_amt[0] ), .Z(n37)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i37_3_lut.init = 16'hcaca;
    LUT4 top_bit_I_0_i39_3_lut (.A(a_for_shift_right[7]), .B(a_for_shift_right[8]), 
         .C(\shift_amt[0] ), .Z(n39)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(88[30:53])
    defparam top_bit_I_0_i39_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i11_3_lut (.A(tmp_data[21]), .B(tmp_data[10]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i14_3_lut (.A(tmp_data[18]), .B(tmp_data[13]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i8_3_lut (.A(tmp_data[24]), .B(tmp_data[7]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 a_0__I_0_i6_3_lut (.A(tmp_data[26]), .B(tmp_data[5]), .C(\alu_op_in[2] ), 
         .Z(a_for_shift_right[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(72[37] 77[8])
    defparam a_0__I_0_i6_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module tinyqv_registers
//

module tinyqv_registers (rd, debug_reg_wen, rs2, n12, n11, n9, n8, 
            rs1, clk_c, return_addr, \registers[5][7] , \registers[6][7] , 
            \registers[7][7] , debug_rd, counter_hi, clk_c_enable_543, 
            mstatus_mie, interrupt_pending_N_1671, n27480, was_early_branch, 
            n26597, n31747, rst_reg_n, n18086, clk_c_enable_348, no_write_in_progress, 
            n27534, time_hi, \cycle_count_wide[6] , \time_count[3] , 
            \cycle_count_wide[4] , \time_count[1] , n28150, n27762, 
            \cycle_count_wide[5] , \time_count[2] , n27018, n28182, 
            n15604, n29747, \data_rs2[1] , n4, \reg_access[3][2] , 
            n33484, \mcause[5] , n28520, n30165, n30166, n30169, 
            n33486, n31748, n32046, n31917, n30167, n31943, clk_c_enable_36, 
            \mepc[0] , \csr_read_3__N_1451[0] , n30168, n11559, \imm[6] , 
            n26121, \mepc[3] , n31171, data_rs1, \data_rs2[0] , \data_rs2[2] , 
            n33494) /* synthesis syn_module_defined=1 */ ;
    input [3:0]rd;
    input debug_reg_wen;
    input [3:0]rs2;
    output n12;
    output n11;
    output n9;
    output n8;
    input [3:0]rs1;
    input clk_c;
    output [23:1]return_addr;
    output \registers[5][7] ;
    output \registers[6][7] ;
    output \registers[7][7] ;
    input [3:0]debug_rd;
    input [4:2]counter_hi;
    output clk_c_enable_543;
    input mstatus_mie;
    input interrupt_pending_N_1671;
    output n27480;
    input was_early_branch;
    input n26597;
    output n31747;
    input rst_reg_n;
    input n18086;
    output clk_c_enable_348;
    input no_write_in_progress;
    output n27534;
    input [2:0]time_hi;
    input \cycle_count_wide[6] ;
    output \time_count[3] ;
    input \cycle_count_wide[4] ;
    output \time_count[1] ;
    input n28150;
    output n27762;
    input \cycle_count_wide[5] ;
    output \time_count[2] ;
    input n27018;
    output n28182;
    output n15604;
    output n29747;
    output \data_rs2[1] ;
    input n4;
    output \reg_access[3][2] ;
    input n33484;
    input \mcause[5] ;
    output n28520;
    output n30165;
    output n30166;
    output n30169;
    input n33486;
    output n31748;
    input n32046;
    output n31917;
    output n30167;
    output n31943;
    output clk_c_enable_36;
    input \mepc[0] ;
    output \csr_read_3__N_1451[0] ;
    output n30168;
    output n11559;
    input \imm[6] ;
    output n26121;
    input \mepc[3] ;
    output n31171;
    output [3:0]data_rs1;
    output \data_rs2[0] ;
    output \data_rs2[2] ;
    output n33494;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire n31752, n31751, n31750, n31749;
    wire [31:0]\registers[14] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[15] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[12] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[13] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[10] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[11] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[8] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[9] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n12_adj_3091, n11_adj_3092, n9_adj_3093, n8_adj_3094, n29725, 
        n29724, n29723, n29722;
    wire [31:0]\registers[6] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    wire [31:0]\registers[7] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n29721;
    wire [31:0]\registers[5] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire n29720, n29710, n29709, n29708, n29707, n29706, n29705, 
        n29673, n29672, n29671, n29670, n29669, n29668, n29644, 
        n29643, n29642, n29641, n29640, n29639;
    wire [31:0]\registers[1] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_1__2__N_1756, registers_1__1__N_1757, registers_1__0__N_1758;
    wire [31:0]\registers[2] ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(29[16:25])
    
    wire registers_2__3__N_1759, registers_2__2__N_1762, registers_2__1__N_1763, 
        registers_2__0__N_1764, registers_5__3__N_1765, registers_5__2__N_1768, 
        registers_5__1__N_1769, registers_5__0__N_1770, registers_6__3__N_1771, 
        registers_6__2__N_1774, registers_6__1__N_1775, registers_6__0__N_1776, 
        registers_7__3__N_1777, registers_7__2__N_1780, registers_7__1__N_1781, 
        registers_7__0__N_1782, registers_8__3__N_1783, registers_8__2__N_1786, 
        registers_8__1__N_1787, registers_8__0__N_1788, registers_9__3__N_1789, 
        registers_9__2__N_1792, registers_9__1__N_1793, registers_9__0__N_1794, 
        registers_10__3__N_1795, registers_10__2__N_1798, registers_10__1__N_1799, 
        registers_10__0__N_1800, registers_11__3__N_1801, registers_11__2__N_1804, 
        registers_11__1__N_1805, registers_11__0__N_1806, registers_12__3__N_1807, 
        registers_12__2__N_1810, registers_12__1__N_1811, registers_12__0__N_1812, 
        registers_13__3__N_1813, registers_13__2__N_1816, registers_13__1__N_1817, 
        registers_13__0__N_1818, registers_14__3__N_1819, registers_14__2__N_1822, 
        registers_14__1__N_1823, registers_14__0__N_1824, registers_15__3__N_1825, 
        registers_15__2__N_1828, registers_15__1__N_1829, registers_15__0__N_1830, 
        registers_1__3__N_1753, n31984, n31985, n29761, n31986, n29667, 
        n29666, n31989, n29703, n29704, n29711, n29718, n29719, 
        n29726, n29762, n29765, n29763, n29764, n29766, n29768, 
        n29769, n29772, n29770, n29771, n29773, n12_adj_3095, n11_adj_3096, 
        n9_adj_3097, n29740, n8_adj_3098, n5, n12_adj_3099, n11_adj_3100, 
        n9_adj_3101, n8_adj_3102, n29637, n29638, n29645, n5_adj_3103, 
        n29647, n29648, n29650, n29676, n29677, n29679, n29713, 
        n29714, n29716, n29728, n29729, n29731, n29742, n29743, 
        n29745, n5_adj_3104, n29741, n29674, n29744, n29646, n29675, 
        n29678, n29712, n29649, n29727, n29715, n29730;
    
    LUT4 i1_2_lut_rep_547_3_lut (.A(rd[1]), .B(rd[0]), .C(debug_reg_wen), 
         .Z(n31752)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_rep_547_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_546_3_lut (.A(rd[1]), .B(debug_reg_wen), .C(rd[0]), 
         .Z(n31751)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_546_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_545_3_lut (.A(rd[1]), .B(rd[0]), .C(debug_reg_wen), 
         .Z(n31750)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_545_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_544_3_lut (.A(rd[1]), .B(debug_reg_wen), .C(rd[0]), 
         .Z(n31749)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_rep_544_3_lut.init = 16'h0404;
    LUT4 rs2_3__I_0_Mux_3_i12_3_lut (.A(\registers[14] [7]), .B(\registers[15] [7]), 
         .C(rs2[0]), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i12_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i11_3_lut (.A(\registers[12] [7]), .B(\registers[13] [7]), 
         .C(rs2[0]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i9_3_lut (.A(\registers[10] [7]), .B(\registers[11] [7]), 
         .C(rs2[0]), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_3_i8_3_lut (.A(\registers[8] [7]), .B(\registers[9] [7]), 
         .C(rs2[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i12_3_lut (.A(\registers[14] [7]), .B(\registers[15] [7]), 
         .C(rs1[0]), .Z(n12_adj_3091)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i12_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i11_3_lut (.A(\registers[12] [7]), .B(\registers[13] [7]), 
         .C(rs1[0]), .Z(n11_adj_3092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i11_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i9_3_lut (.A(\registers[10] [7]), .B(\registers[11] [7]), 
         .C(rs1[0]), .Z(n9_adj_3093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_3_i8_3_lut (.A(\registers[8] [7]), .B(\registers[9] [7]), 
         .C(rs1[0]), .Z(n8_adj_3094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 i27108_3_lut (.A(\registers[14] [6]), .B(\registers[15] [6]), .C(rs2[0]), 
         .Z(n29725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27108_3_lut.init = 16'hcaca;
    LUT4 i27107_3_lut (.A(\registers[12] [6]), .B(\registers[13] [6]), .C(rs2[0]), 
         .Z(n29724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27107_3_lut.init = 16'hcaca;
    LUT4 i27106_3_lut (.A(\registers[10] [6]), .B(\registers[11] [6]), .C(rs2[0]), 
         .Z(n29723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27106_3_lut.init = 16'hcaca;
    LUT4 i27105_3_lut (.A(\registers[8] [6]), .B(\registers[9] [6]), .C(rs2[0]), 
         .Z(n29722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27105_3_lut.init = 16'hcaca;
    LUT4 i27104_3_lut (.A(\registers[6] [6]), .B(\registers[7] [6]), .C(rs2[0]), 
         .Z(n29721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27104_3_lut.init = 16'hcaca;
    LUT4 i27103_3_lut (.A(\registers[5] [6]), .B(rs2[0]), .Z(n29720)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27103_3_lut.init = 16'h8888;
    LUT4 i27093_3_lut (.A(\registers[14] [6]), .B(\registers[15] [6]), .C(rs1[0]), 
         .Z(n29710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27093_3_lut.init = 16'hcaca;
    LUT4 i27092_3_lut (.A(\registers[12] [6]), .B(\registers[13] [6]), .C(rs1[0]), 
         .Z(n29709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27092_3_lut.init = 16'hcaca;
    LUT4 i27091_3_lut (.A(\registers[10] [6]), .B(\registers[11] [6]), .C(rs1[0]), 
         .Z(n29708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27091_3_lut.init = 16'hcaca;
    LUT4 i27090_3_lut (.A(\registers[8] [6]), .B(\registers[9] [6]), .C(rs1[0]), 
         .Z(n29707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27090_3_lut.init = 16'hcaca;
    LUT4 i27089_3_lut (.A(\registers[6] [6]), .B(\registers[7] [6]), .C(rs1[0]), 
         .Z(n29706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27089_3_lut.init = 16'hcaca;
    LUT4 i27088_3_lut (.A(\registers[5] [6]), .B(rs1[0]), .Z(n29705)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27088_3_lut.init = 16'h8888;
    LUT4 i27056_3_lut (.A(\registers[14] [4]), .B(\registers[15] [4]), .C(rs1[0]), 
         .Z(n29673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27056_3_lut.init = 16'hcaca;
    LUT4 i27055_3_lut (.A(\registers[12] [4]), .B(\registers[13] [4]), .C(rs1[0]), 
         .Z(n29672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27055_3_lut.init = 16'hcaca;
    LUT4 i27054_3_lut (.A(\registers[10] [4]), .B(\registers[11] [4]), .C(rs1[0]), 
         .Z(n29671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27054_3_lut.init = 16'hcaca;
    LUT4 i27053_3_lut (.A(\registers[8] [4]), .B(\registers[9] [4]), .C(rs1[0]), 
         .Z(n29670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27053_3_lut.init = 16'hcaca;
    LUT4 i27052_3_lut (.A(\registers[6] [4]), .B(\registers[7] [4]), .C(rs1[0]), 
         .Z(n29669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27052_3_lut.init = 16'hcaca;
    LUT4 i27051_3_lut (.A(\registers[5] [4]), .B(rs1[0]), .Z(n29668)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27051_3_lut.init = 16'h8888;
    LUT4 i27027_3_lut (.A(\registers[14] [4]), .B(\registers[15] [4]), .C(rs2[0]), 
         .Z(n29644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27027_3_lut.init = 16'hcaca;
    LUT4 i27026_3_lut (.A(\registers[12] [4]), .B(\registers[13] [4]), .C(rs2[0]), 
         .Z(n29643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27026_3_lut.init = 16'hcaca;
    LUT4 i27025_3_lut (.A(\registers[10] [4]), .B(\registers[11] [4]), .C(rs2[0]), 
         .Z(n29642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27025_3_lut.init = 16'hcaca;
    LUT4 i27024_3_lut (.A(\registers[8] [4]), .B(\registers[9] [4]), .C(rs2[0]), 
         .Z(n29641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27024_3_lut.init = 16'hcaca;
    LUT4 i27023_3_lut (.A(\registers[6] [4]), .B(\registers[7] [4]), .C(rs2[0]), 
         .Z(n29640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27023_3_lut.init = 16'hcaca;
    LUT4 i27022_3_lut (.A(\registers[5] [4]), .B(rs2[0]), .Z(n29639)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27022_3_lut.init = 16'h8888;
    FD1S3AX \registers_1[[2__504  (.D(registers_1__2__N_1756), .CK(clk_c), 
            .Q(\registers[1] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[2__504 .GSR = "DISABLED";
    FD1S3AX \registers_1[[1__505  (.D(registers_1__1__N_1757), .CK(clk_c), 
            .Q(\registers[1] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[1__505 .GSR = "DISABLED";
    FD1S3AX \registers_1[[0__506  (.D(registers_1__0__N_1758), .CK(clk_c), 
            .Q(\registers[1] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[0__506 .GSR = "DISABLED";
    FD1S3AX \registers_1[[31__507  (.D(\registers[1] [3]), .CK(clk_c), .Q(return_addr[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[31__507 .GSR = "DISABLED";
    FD1S3AX \registers_1[[30__508  (.D(\registers[1] [2]), .CK(clk_c), .Q(return_addr[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[30__508 .GSR = "DISABLED";
    FD1S3AX \registers_1[[29__509  (.D(\registers[1] [1]), .CK(clk_c), .Q(return_addr[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[29__509 .GSR = "DISABLED";
    FD1S3AX \registers_1[[28__510  (.D(\registers[1] [0]), .CK(clk_c), .Q(return_addr[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[28__510 .GSR = "DISABLED";
    FD1S3AX \registers_1[[27__511  (.D(return_addr[23]), .CK(clk_c), .Q(return_addr[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[27__511 .GSR = "DISABLED";
    FD1S3AX \registers_1[[26__512  (.D(return_addr[22]), .CK(clk_c), .Q(return_addr[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[26__512 .GSR = "DISABLED";
    FD1S3AX \registers_1[[25__513  (.D(return_addr[21]), .CK(clk_c), .Q(return_addr[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[25__513 .GSR = "DISABLED";
    FD1S3AX \registers_1[[24__514  (.D(return_addr[20]), .CK(clk_c), .Q(return_addr[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[24__514 .GSR = "DISABLED";
    FD1S3AX \registers_1[[23__515  (.D(return_addr[19]), .CK(clk_c), .Q(return_addr[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[23__515 .GSR = "DISABLED";
    FD1S3AX \registers_1[[22__516  (.D(return_addr[18]), .CK(clk_c), .Q(return_addr[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[22__516 .GSR = "DISABLED";
    FD1S3AX \registers_1[[21__517  (.D(return_addr[17]), .CK(clk_c), .Q(return_addr[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[21__517 .GSR = "DISABLED";
    FD1S3AX \registers_1[[20__518  (.D(return_addr[16]), .CK(clk_c), .Q(return_addr[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[20__518 .GSR = "DISABLED";
    FD1S3AX \registers_1[[19__519  (.D(return_addr[15]), .CK(clk_c), .Q(return_addr[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[19__519 .GSR = "DISABLED";
    FD1S3AX \registers_1[[18__520  (.D(return_addr[14]), .CK(clk_c), .Q(return_addr[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[18__520 .GSR = "DISABLED";
    FD1S3AX \registers_1[[17__521  (.D(return_addr[13]), .CK(clk_c), .Q(return_addr[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[17__521 .GSR = "DISABLED";
    FD1S3AX \registers_1[[16__522  (.D(return_addr[12]), .CK(clk_c), .Q(return_addr[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[16__522 .GSR = "DISABLED";
    FD1S3AX \registers_1[[15__523  (.D(return_addr[11]), .CK(clk_c), .Q(return_addr[7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[15__523 .GSR = "DISABLED";
    FD1S3AX \registers_1[[14__524  (.D(return_addr[10]), .CK(clk_c), .Q(return_addr[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[14__524 .GSR = "DISABLED";
    FD1S3AX \registers_1[[13__525  (.D(return_addr[9]), .CK(clk_c), .Q(return_addr[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[13__525 .GSR = "DISABLED";
    FD1S3AX \registers_1[[12__526  (.D(return_addr[8]), .CK(clk_c), .Q(return_addr[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[12__526 .GSR = "DISABLED";
    FD1S3AX \registers_1[[11__527  (.D(return_addr[7]), .CK(clk_c), .Q(return_addr[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[11__527 .GSR = "DISABLED";
    FD1S3AX \registers_1[[10__528  (.D(return_addr[6]), .CK(clk_c), .Q(return_addr[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[10__528 .GSR = "DISABLED";
    FD1S3AX \registers_1[[9__529  (.D(return_addr[5]), .CK(clk_c), .Q(return_addr[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[9__529 .GSR = "DISABLED";
    FD1S3AX \registers_1[[8__530  (.D(return_addr[4]), .CK(clk_c), .Q(\registers[1] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[8__530 .GSR = "DISABLED";
    FD1S3AX \registers_1[[7__531  (.D(return_addr[3]), .CK(clk_c), .Q(\registers[1] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[7__531 .GSR = "DISABLED";
    FD1S3AX \registers_1[[6__532  (.D(return_addr[2]), .CK(clk_c), .Q(\registers[1] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[6__532 .GSR = "DISABLED";
    FD1S3AX \registers_1[[5__533  (.D(return_addr[1]), .CK(clk_c), .Q(\registers[1] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[5__533 .GSR = "DISABLED";
    FD1S3AX \registers_1[[4__534  (.D(\registers[1] [8]), .CK(clk_c), .Q(\registers[1] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_1[[4__534 .GSR = "DISABLED";
    FD1S3AX \registers_2[[3__535  (.D(registers_2__3__N_1759), .CK(clk_c), 
            .Q(\registers[2] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[3__535 .GSR = "DISABLED";
    FD1S3AX \registers_2[[2__536  (.D(registers_2__2__N_1762), .CK(clk_c), 
            .Q(\registers[2] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[2__536 .GSR = "DISABLED";
    FD1S3AX \registers_2[[1__537  (.D(registers_2__1__N_1763), .CK(clk_c), 
            .Q(\registers[2] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[1__537 .GSR = "DISABLED";
    FD1S3AX \registers_2[[0__538  (.D(registers_2__0__N_1764), .CK(clk_c), 
            .Q(\registers[2] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_2[[0__538 .GSR = "DISABLED";
    FD1S3AX \registers_2[[31__539  (.D(\registers[2] [3]), .CK(clk_c), .Q(\registers[2] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[31__539 .GSR = "DISABLED";
    FD1S3AX \registers_2[[30__540  (.D(\registers[2] [2]), .CK(clk_c), .Q(\registers[2] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[30__540 .GSR = "DISABLED";
    FD1S3AX \registers_2[[29__541  (.D(\registers[2] [1]), .CK(clk_c), .Q(\registers[2] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[29__541 .GSR = "DISABLED";
    FD1S3AX \registers_2[[28__542  (.D(\registers[2] [0]), .CK(clk_c), .Q(\registers[2] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[28__542 .GSR = "DISABLED";
    FD1S3AX \registers_2[[27__543  (.D(\registers[2] [31]), .CK(clk_c), 
            .Q(\registers[2] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[27__543 .GSR = "DISABLED";
    FD1S3AX \registers_2[[26__544  (.D(\registers[2] [30]), .CK(clk_c), 
            .Q(\registers[2] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[26__544 .GSR = "DISABLED";
    FD1S3AX \registers_2[[25__545  (.D(\registers[2] [29]), .CK(clk_c), 
            .Q(\registers[2] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[25__545 .GSR = "DISABLED";
    FD1S3AX \registers_2[[24__546  (.D(\registers[2] [28]), .CK(clk_c), 
            .Q(\registers[2] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[24__546 .GSR = "DISABLED";
    FD1S3AX \registers_2[[23__547  (.D(\registers[2] [27]), .CK(clk_c), 
            .Q(\registers[2] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[23__547 .GSR = "DISABLED";
    FD1S3AX \registers_2[[22__548  (.D(\registers[2] [26]), .CK(clk_c), 
            .Q(\registers[2] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[22__548 .GSR = "DISABLED";
    FD1S3AX \registers_2[[21__549  (.D(\registers[2] [25]), .CK(clk_c), 
            .Q(\registers[2] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[21__549 .GSR = "DISABLED";
    FD1S3AX \registers_2[[20__550  (.D(\registers[2] [24]), .CK(clk_c), 
            .Q(\registers[2] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[20__550 .GSR = "DISABLED";
    FD1S3AX \registers_2[[19__551  (.D(\registers[2] [23]), .CK(clk_c), 
            .Q(\registers[2] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[19__551 .GSR = "DISABLED";
    FD1S3AX \registers_2[[18__552  (.D(\registers[2] [22]), .CK(clk_c), 
            .Q(\registers[2] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[18__552 .GSR = "DISABLED";
    FD1S3AX \registers_2[[17__553  (.D(\registers[2] [21]), .CK(clk_c), 
            .Q(\registers[2] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[17__553 .GSR = "DISABLED";
    FD1S3AX \registers_2[[16__554  (.D(\registers[2] [20]), .CK(clk_c), 
            .Q(\registers[2] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[16__554 .GSR = "DISABLED";
    FD1S3AX \registers_2[[15__555  (.D(\registers[2] [19]), .CK(clk_c), 
            .Q(\registers[2] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[15__555 .GSR = "DISABLED";
    FD1S3AX \registers_2[[14__556  (.D(\registers[2] [18]), .CK(clk_c), 
            .Q(\registers[2] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[14__556 .GSR = "DISABLED";
    FD1S3AX \registers_2[[13__557  (.D(\registers[2] [17]), .CK(clk_c), 
            .Q(\registers[2] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[13__557 .GSR = "DISABLED";
    FD1S3AX \registers_2[[12__558  (.D(\registers[2] [16]), .CK(clk_c), 
            .Q(\registers[2] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[12__558 .GSR = "DISABLED";
    FD1S3AX \registers_2[[11__559  (.D(\registers[2] [15]), .CK(clk_c), 
            .Q(\registers[2] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[11__559 .GSR = "DISABLED";
    FD1S3AX \registers_2[[10__560  (.D(\registers[2] [14]), .CK(clk_c), 
            .Q(\registers[2] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[10__560 .GSR = "DISABLED";
    FD1S3AX \registers_2[[9__561  (.D(\registers[2] [13]), .CK(clk_c), .Q(\registers[2] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[9__561 .GSR = "DISABLED";
    FD1S3AX \registers_2[[8__562  (.D(\registers[2] [12]), .CK(clk_c), .Q(\registers[2] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[8__562 .GSR = "DISABLED";
    FD1S3AX \registers_2[[7__563  (.D(\registers[2] [11]), .CK(clk_c), .Q(\registers[2] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[7__563 .GSR = "DISABLED";
    FD1S3AX \registers_2[[6__564  (.D(\registers[2] [10]), .CK(clk_c), .Q(\registers[2] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[6__564 .GSR = "DISABLED";
    FD1S3AX \registers_2[[5__565  (.D(\registers[2] [9]), .CK(clk_c), .Q(\registers[2] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[5__565 .GSR = "DISABLED";
    FD1S3AX \registers_2[[4__566  (.D(\registers[2] [8]), .CK(clk_c), .Q(\registers[2] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_2[[4__566 .GSR = "DISABLED";
    FD1S3AX \registers_5[[3__567  (.D(registers_5__3__N_1765), .CK(clk_c), 
            .Q(\registers[5] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[3__567 .GSR = "DISABLED";
    FD1S3AX \registers_5[[2__568  (.D(registers_5__2__N_1768), .CK(clk_c), 
            .Q(\registers[5] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[2__568 .GSR = "DISABLED";
    FD1S3AX \registers_5[[1__569  (.D(registers_5__1__N_1769), .CK(clk_c), 
            .Q(\registers[5] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[1__569 .GSR = "DISABLED";
    FD1S3AX \registers_5[[0__570  (.D(registers_5__0__N_1770), .CK(clk_c), 
            .Q(\registers[5] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_5[[0__570 .GSR = "DISABLED";
    FD1S3AX \registers_5[[31__571  (.D(\registers[5] [3]), .CK(clk_c), .Q(\registers[5] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[31__571 .GSR = "DISABLED";
    FD1S3AX \registers_5[[30__572  (.D(\registers[5] [2]), .CK(clk_c), .Q(\registers[5] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[30__572 .GSR = "DISABLED";
    FD1S3AX \registers_5[[29__573  (.D(\registers[5] [1]), .CK(clk_c), .Q(\registers[5] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[29__573 .GSR = "DISABLED";
    FD1S3AX \registers_5[[28__574  (.D(\registers[5] [0]), .CK(clk_c), .Q(\registers[5] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[28__574 .GSR = "DISABLED";
    FD1S3AX \registers_5[[27__575  (.D(\registers[5] [31]), .CK(clk_c), 
            .Q(\registers[5] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[27__575 .GSR = "DISABLED";
    FD1S3AX \registers_5[[26__576  (.D(\registers[5] [30]), .CK(clk_c), 
            .Q(\registers[5] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[26__576 .GSR = "DISABLED";
    FD1S3AX \registers_5[[25__577  (.D(\registers[5] [29]), .CK(clk_c), 
            .Q(\registers[5] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[25__577 .GSR = "DISABLED";
    FD1S3AX \registers_5[[24__578  (.D(\registers[5] [28]), .CK(clk_c), 
            .Q(\registers[5] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[24__578 .GSR = "DISABLED";
    FD1S3AX \registers_5[[23__579  (.D(\registers[5] [27]), .CK(clk_c), 
            .Q(\registers[5] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[23__579 .GSR = "DISABLED";
    FD1S3AX \registers_5[[22__580  (.D(\registers[5] [26]), .CK(clk_c), 
            .Q(\registers[5] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[22__580 .GSR = "DISABLED";
    FD1S3AX \registers_5[[21__581  (.D(\registers[5] [25]), .CK(clk_c), 
            .Q(\registers[5] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[21__581 .GSR = "DISABLED";
    FD1S3AX \registers_5[[20__582  (.D(\registers[5] [24]), .CK(clk_c), 
            .Q(\registers[5] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[20__582 .GSR = "DISABLED";
    FD1S3AX \registers_5[[19__583  (.D(\registers[5] [23]), .CK(clk_c), 
            .Q(\registers[5] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[19__583 .GSR = "DISABLED";
    FD1S3AX \registers_5[[18__584  (.D(\registers[5] [22]), .CK(clk_c), 
            .Q(\registers[5] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[18__584 .GSR = "DISABLED";
    FD1S3AX \registers_5[[17__585  (.D(\registers[5] [21]), .CK(clk_c), 
            .Q(\registers[5] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[17__585 .GSR = "DISABLED";
    FD1S3AX \registers_5[[16__586  (.D(\registers[5] [20]), .CK(clk_c), 
            .Q(\registers[5] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[16__586 .GSR = "DISABLED";
    FD1S3AX \registers_5[[15__587  (.D(\registers[5] [19]), .CK(clk_c), 
            .Q(\registers[5] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[15__587 .GSR = "DISABLED";
    FD1S3AX \registers_5[[14__588  (.D(\registers[5] [18]), .CK(clk_c), 
            .Q(\registers[5] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[14__588 .GSR = "DISABLED";
    FD1S3AX \registers_5[[13__589  (.D(\registers[5] [17]), .CK(clk_c), 
            .Q(\registers[5] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[13__589 .GSR = "DISABLED";
    FD1S3AX \registers_5[[12__590  (.D(\registers[5] [16]), .CK(clk_c), 
            .Q(\registers[5] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[12__590 .GSR = "DISABLED";
    FD1S3AX \registers_5[[11__591  (.D(\registers[5] [15]), .CK(clk_c), 
            .Q(\registers[5] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[11__591 .GSR = "DISABLED";
    FD1S3AX \registers_5[[10__592  (.D(\registers[5] [14]), .CK(clk_c), 
            .Q(\registers[5] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[10__592 .GSR = "DISABLED";
    FD1S3AX \registers_5[[9__593  (.D(\registers[5] [13]), .CK(clk_c), .Q(\registers[5] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[9__593 .GSR = "DISABLED";
    FD1S3AX \registers_5[[8__594  (.D(\registers[5] [12]), .CK(clk_c), .Q(\registers[5] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[8__594 .GSR = "DISABLED";
    FD1S3AX \registers_5[[7__595  (.D(\registers[5] [11]), .CK(clk_c), .Q(\registers[5][7] )) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[7__595 .GSR = "DISABLED";
    FD1S3AX \registers_5[[6__596  (.D(\registers[5] [10]), .CK(clk_c), .Q(\registers[5] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[6__596 .GSR = "DISABLED";
    FD1S3AX \registers_5[[5__597  (.D(\registers[5] [9]), .CK(clk_c), .Q(\registers[5] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[5__597 .GSR = "DISABLED";
    FD1S3AX \registers_5[[4__598  (.D(\registers[5] [8]), .CK(clk_c), .Q(\registers[5] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_5[[4__598 .GSR = "DISABLED";
    FD1S3AX \registers_6[[3__599  (.D(registers_6__3__N_1771), .CK(clk_c), 
            .Q(\registers[6] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[3__599 .GSR = "DISABLED";
    FD1S3AX \registers_6[[2__600  (.D(registers_6__2__N_1774), .CK(clk_c), 
            .Q(\registers[6] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[2__600 .GSR = "DISABLED";
    FD1S3AX \registers_6[[1__601  (.D(registers_6__1__N_1775), .CK(clk_c), 
            .Q(\registers[6] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[1__601 .GSR = "DISABLED";
    FD1S3AX \registers_6[[0__602  (.D(registers_6__0__N_1776), .CK(clk_c), 
            .Q(\registers[6] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_6[[0__602 .GSR = "DISABLED";
    FD1S3AX \registers_6[[31__603  (.D(\registers[6] [3]), .CK(clk_c), .Q(\registers[6] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[31__603 .GSR = "DISABLED";
    FD1S3AX \registers_6[[30__604  (.D(\registers[6] [2]), .CK(clk_c), .Q(\registers[6] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[30__604 .GSR = "DISABLED";
    FD1S3AX \registers_6[[29__605  (.D(\registers[6] [1]), .CK(clk_c), .Q(\registers[6] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[29__605 .GSR = "DISABLED";
    FD1S3AX \registers_6[[28__606  (.D(\registers[6] [0]), .CK(clk_c), .Q(\registers[6] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[28__606 .GSR = "DISABLED";
    FD1S3AX \registers_6[[27__607  (.D(\registers[6] [31]), .CK(clk_c), 
            .Q(\registers[6] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[27__607 .GSR = "DISABLED";
    FD1S3AX \registers_6[[26__608  (.D(\registers[6] [30]), .CK(clk_c), 
            .Q(\registers[6] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[26__608 .GSR = "DISABLED";
    FD1S3AX \registers_6[[25__609  (.D(\registers[6] [29]), .CK(clk_c), 
            .Q(\registers[6] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[25__609 .GSR = "DISABLED";
    FD1S3AX \registers_6[[24__610  (.D(\registers[6] [28]), .CK(clk_c), 
            .Q(\registers[6] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[24__610 .GSR = "DISABLED";
    FD1S3AX \registers_6[[23__611  (.D(\registers[6] [27]), .CK(clk_c), 
            .Q(\registers[6] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[23__611 .GSR = "DISABLED";
    FD1S3AX \registers_6[[22__612  (.D(\registers[6] [26]), .CK(clk_c), 
            .Q(\registers[6] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[22__612 .GSR = "DISABLED";
    FD1S3AX \registers_6[[21__613  (.D(\registers[6] [25]), .CK(clk_c), 
            .Q(\registers[6] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[21__613 .GSR = "DISABLED";
    FD1S3AX \registers_6[[20__614  (.D(\registers[6] [24]), .CK(clk_c), 
            .Q(\registers[6] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[20__614 .GSR = "DISABLED";
    FD1S3AX \registers_6[[19__615  (.D(\registers[6] [23]), .CK(clk_c), 
            .Q(\registers[6] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[19__615 .GSR = "DISABLED";
    FD1S3AX \registers_6[[18__616  (.D(\registers[6] [22]), .CK(clk_c), 
            .Q(\registers[6] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[18__616 .GSR = "DISABLED";
    FD1S3AX \registers_6[[17__617  (.D(\registers[6] [21]), .CK(clk_c), 
            .Q(\registers[6] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[17__617 .GSR = "DISABLED";
    FD1S3AX \registers_6[[16__618  (.D(\registers[6] [20]), .CK(clk_c), 
            .Q(\registers[6] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[16__618 .GSR = "DISABLED";
    FD1S3AX \registers_6[[15__619  (.D(\registers[6] [19]), .CK(clk_c), 
            .Q(\registers[6] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[15__619 .GSR = "DISABLED";
    FD1S3AX \registers_6[[14__620  (.D(\registers[6] [18]), .CK(clk_c), 
            .Q(\registers[6] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[14__620 .GSR = "DISABLED";
    FD1S3AX \registers_6[[13__621  (.D(\registers[6] [17]), .CK(clk_c), 
            .Q(\registers[6] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[13__621 .GSR = "DISABLED";
    FD1S3AX \registers_6[[12__622  (.D(\registers[6] [16]), .CK(clk_c), 
            .Q(\registers[6] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[12__622 .GSR = "DISABLED";
    FD1S3AX \registers_6[[11__623  (.D(\registers[6] [15]), .CK(clk_c), 
            .Q(\registers[6] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[11__623 .GSR = "DISABLED";
    FD1S3AX \registers_6[[10__624  (.D(\registers[6] [14]), .CK(clk_c), 
            .Q(\registers[6] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[10__624 .GSR = "DISABLED";
    FD1S3AX \registers_6[[9__625  (.D(\registers[6] [13]), .CK(clk_c), .Q(\registers[6] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[9__625 .GSR = "DISABLED";
    FD1S3AX \registers_6[[8__626  (.D(\registers[6] [12]), .CK(clk_c), .Q(\registers[6] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[8__626 .GSR = "DISABLED";
    FD1S3AX \registers_6[[7__627  (.D(\registers[6] [11]), .CK(clk_c), .Q(\registers[6][7] )) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[7__627 .GSR = "DISABLED";
    FD1S3AX \registers_6[[6__628  (.D(\registers[6] [10]), .CK(clk_c), .Q(\registers[6] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[6__628 .GSR = "DISABLED";
    FD1S3AX \registers_6[[5__629  (.D(\registers[6] [9]), .CK(clk_c), .Q(\registers[6] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[5__629 .GSR = "DISABLED";
    FD1S3AX \registers_6[[4__630  (.D(\registers[6] [8]), .CK(clk_c), .Q(\registers[6] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_6[[4__630 .GSR = "DISABLED";
    FD1S3AX \registers_7[[3__631  (.D(registers_7__3__N_1777), .CK(clk_c), 
            .Q(\registers[7] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[3__631 .GSR = "DISABLED";
    FD1S3AX \registers_7[[2__632  (.D(registers_7__2__N_1780), .CK(clk_c), 
            .Q(\registers[7] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[2__632 .GSR = "DISABLED";
    FD1S3AX \registers_7[[1__633  (.D(registers_7__1__N_1781), .CK(clk_c), 
            .Q(\registers[7] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[1__633 .GSR = "DISABLED";
    FD1S3AX \registers_7[[0__634  (.D(registers_7__0__N_1782), .CK(clk_c), 
            .Q(\registers[7] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_7[[0__634 .GSR = "DISABLED";
    FD1S3AX \registers_7[[31__635  (.D(\registers[7] [3]), .CK(clk_c), .Q(\registers[7] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[31__635 .GSR = "DISABLED";
    FD1S3AX \registers_7[[30__636  (.D(\registers[7] [2]), .CK(clk_c), .Q(\registers[7] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[30__636 .GSR = "DISABLED";
    FD1S3AX \registers_7[[29__637  (.D(\registers[7] [1]), .CK(clk_c), .Q(\registers[7] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[29__637 .GSR = "DISABLED";
    FD1S3AX \registers_7[[28__638  (.D(\registers[7] [0]), .CK(clk_c), .Q(\registers[7] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[28__638 .GSR = "DISABLED";
    FD1S3AX \registers_7[[27__639  (.D(\registers[7] [31]), .CK(clk_c), 
            .Q(\registers[7] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[27__639 .GSR = "DISABLED";
    FD1S3AX \registers_7[[26__640  (.D(\registers[7] [30]), .CK(clk_c), 
            .Q(\registers[7] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[26__640 .GSR = "DISABLED";
    FD1S3AX \registers_7[[25__641  (.D(\registers[7] [29]), .CK(clk_c), 
            .Q(\registers[7] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[25__641 .GSR = "DISABLED";
    FD1S3AX \registers_7[[24__642  (.D(\registers[7] [28]), .CK(clk_c), 
            .Q(\registers[7] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[24__642 .GSR = "DISABLED";
    FD1S3AX \registers_7[[23__643  (.D(\registers[7] [27]), .CK(clk_c), 
            .Q(\registers[7] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[23__643 .GSR = "DISABLED";
    FD1S3AX \registers_7[[22__644  (.D(\registers[7] [26]), .CK(clk_c), 
            .Q(\registers[7] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[22__644 .GSR = "DISABLED";
    FD1S3AX \registers_7[[21__645  (.D(\registers[7] [25]), .CK(clk_c), 
            .Q(\registers[7] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[21__645 .GSR = "DISABLED";
    FD1S3AX \registers_7[[20__646  (.D(\registers[7] [24]), .CK(clk_c), 
            .Q(\registers[7] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[20__646 .GSR = "DISABLED";
    FD1S3AX \registers_7[[19__647  (.D(\registers[7] [23]), .CK(clk_c), 
            .Q(\registers[7] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[19__647 .GSR = "DISABLED";
    FD1S3AX \registers_7[[18__648  (.D(\registers[7] [22]), .CK(clk_c), 
            .Q(\registers[7] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[18__648 .GSR = "DISABLED";
    FD1S3AX \registers_7[[17__649  (.D(\registers[7] [21]), .CK(clk_c), 
            .Q(\registers[7] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[17__649 .GSR = "DISABLED";
    FD1S3AX \registers_7[[16__650  (.D(\registers[7] [20]), .CK(clk_c), 
            .Q(\registers[7] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[16__650 .GSR = "DISABLED";
    FD1S3AX \registers_7[[15__651  (.D(\registers[7] [19]), .CK(clk_c), 
            .Q(\registers[7] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[15__651 .GSR = "DISABLED";
    FD1S3AX \registers_7[[14__652  (.D(\registers[7] [18]), .CK(clk_c), 
            .Q(\registers[7] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[14__652 .GSR = "DISABLED";
    FD1S3AX \registers_7[[13__653  (.D(\registers[7] [17]), .CK(clk_c), 
            .Q(\registers[7] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[13__653 .GSR = "DISABLED";
    FD1S3AX \registers_7[[12__654  (.D(\registers[7] [16]), .CK(clk_c), 
            .Q(\registers[7] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[12__654 .GSR = "DISABLED";
    FD1S3AX \registers_7[[11__655  (.D(\registers[7] [15]), .CK(clk_c), 
            .Q(\registers[7] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[11__655 .GSR = "DISABLED";
    FD1S3AX \registers_7[[10__656  (.D(\registers[7] [14]), .CK(clk_c), 
            .Q(\registers[7] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[10__656 .GSR = "DISABLED";
    FD1S3AX \registers_7[[9__657  (.D(\registers[7] [13]), .CK(clk_c), .Q(\registers[7] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[9__657 .GSR = "DISABLED";
    FD1S3AX \registers_7[[8__658  (.D(\registers[7] [12]), .CK(clk_c), .Q(\registers[7] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[8__658 .GSR = "DISABLED";
    FD1S3AX \registers_7[[7__659  (.D(\registers[7] [11]), .CK(clk_c), .Q(\registers[7][7] )) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[7__659 .GSR = "DISABLED";
    FD1S3AX \registers_7[[6__660  (.D(\registers[7] [10]), .CK(clk_c), .Q(\registers[7] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[6__660 .GSR = "DISABLED";
    FD1S3AX \registers_7[[5__661  (.D(\registers[7] [9]), .CK(clk_c), .Q(\registers[7] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[5__661 .GSR = "DISABLED";
    FD1S3AX \registers_7[[4__662  (.D(\registers[7] [8]), .CK(clk_c), .Q(\registers[7] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_7[[4__662 .GSR = "DISABLED";
    FD1S3AX \registers_8[[3__663  (.D(registers_8__3__N_1783), .CK(clk_c), 
            .Q(\registers[8] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[3__663 .GSR = "DISABLED";
    FD1S3AX \registers_8[[2__664  (.D(registers_8__2__N_1786), .CK(clk_c), 
            .Q(\registers[8] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[2__664 .GSR = "DISABLED";
    FD1S3AX \registers_8[[1__665  (.D(registers_8__1__N_1787), .CK(clk_c), 
            .Q(\registers[8] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[1__665 .GSR = "DISABLED";
    FD1S3AX \registers_8[[0__666  (.D(registers_8__0__N_1788), .CK(clk_c), 
            .Q(\registers[8] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_8[[0__666 .GSR = "DISABLED";
    FD1S3AX \registers_8[[31__667  (.D(\registers[8] [3]), .CK(clk_c), .Q(\registers[8] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[31__667 .GSR = "DISABLED";
    FD1S3AX \registers_8[[30__668  (.D(\registers[8] [2]), .CK(clk_c), .Q(\registers[8] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[30__668 .GSR = "DISABLED";
    FD1S3AX \registers_8[[29__669  (.D(\registers[8] [1]), .CK(clk_c), .Q(\registers[8] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[29__669 .GSR = "DISABLED";
    FD1S3AX \registers_8[[28__670  (.D(\registers[8] [0]), .CK(clk_c), .Q(\registers[8] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[28__670 .GSR = "DISABLED";
    FD1S3AX \registers_8[[27__671  (.D(\registers[8] [31]), .CK(clk_c), 
            .Q(\registers[8] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[27__671 .GSR = "DISABLED";
    FD1S3AX \registers_8[[26__672  (.D(\registers[8] [30]), .CK(clk_c), 
            .Q(\registers[8] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[26__672 .GSR = "DISABLED";
    FD1S3AX \registers_8[[25__673  (.D(\registers[8] [29]), .CK(clk_c), 
            .Q(\registers[8] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[25__673 .GSR = "DISABLED";
    FD1S3AX \registers_8[[24__674  (.D(\registers[8] [28]), .CK(clk_c), 
            .Q(\registers[8] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[24__674 .GSR = "DISABLED";
    FD1S3AX \registers_8[[23__675  (.D(\registers[8] [27]), .CK(clk_c), 
            .Q(\registers[8] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[23__675 .GSR = "DISABLED";
    FD1S3AX \registers_8[[22__676  (.D(\registers[8] [26]), .CK(clk_c), 
            .Q(\registers[8] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[22__676 .GSR = "DISABLED";
    FD1S3AX \registers_8[[21__677  (.D(\registers[8] [25]), .CK(clk_c), 
            .Q(\registers[8] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[21__677 .GSR = "DISABLED";
    FD1S3AX \registers_8[[20__678  (.D(\registers[8] [24]), .CK(clk_c), 
            .Q(\registers[8] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[20__678 .GSR = "DISABLED";
    FD1S3AX \registers_8[[19__679  (.D(\registers[8] [23]), .CK(clk_c), 
            .Q(\registers[8] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[19__679 .GSR = "DISABLED";
    FD1S3AX \registers_8[[18__680  (.D(\registers[8] [22]), .CK(clk_c), 
            .Q(\registers[8] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[18__680 .GSR = "DISABLED";
    FD1S3AX \registers_8[[17__681  (.D(\registers[8] [21]), .CK(clk_c), 
            .Q(\registers[8] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[17__681 .GSR = "DISABLED";
    FD1S3AX \registers_8[[16__682  (.D(\registers[8] [20]), .CK(clk_c), 
            .Q(\registers[8] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[16__682 .GSR = "DISABLED";
    FD1S3AX \registers_8[[15__683  (.D(\registers[8] [19]), .CK(clk_c), 
            .Q(\registers[8] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[15__683 .GSR = "DISABLED";
    FD1S3AX \registers_8[[14__684  (.D(\registers[8] [18]), .CK(clk_c), 
            .Q(\registers[8] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[14__684 .GSR = "DISABLED";
    FD1S3AX \registers_8[[13__685  (.D(\registers[8] [17]), .CK(clk_c), 
            .Q(\registers[8] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[13__685 .GSR = "DISABLED";
    FD1S3AX \registers_8[[12__686  (.D(\registers[8] [16]), .CK(clk_c), 
            .Q(\registers[8] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[12__686 .GSR = "DISABLED";
    FD1S3AX \registers_8[[11__687  (.D(\registers[8] [15]), .CK(clk_c), 
            .Q(\registers[8] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[11__687 .GSR = "DISABLED";
    FD1S3AX \registers_8[[10__688  (.D(\registers[8] [14]), .CK(clk_c), 
            .Q(\registers[8] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[10__688 .GSR = "DISABLED";
    FD1S3AX \registers_8[[9__689  (.D(\registers[8] [13]), .CK(clk_c), .Q(\registers[8] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[9__689 .GSR = "DISABLED";
    FD1S3AX \registers_8[[8__690  (.D(\registers[8] [12]), .CK(clk_c), .Q(\registers[8] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[8__690 .GSR = "DISABLED";
    FD1S3AX \registers_8[[7__691  (.D(\registers[8] [11]), .CK(clk_c), .Q(\registers[8] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[7__691 .GSR = "DISABLED";
    FD1S3AX \registers_8[[6__692  (.D(\registers[8] [10]), .CK(clk_c), .Q(\registers[8] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[6__692 .GSR = "DISABLED";
    FD1S3AX \registers_8[[5__693  (.D(\registers[8] [9]), .CK(clk_c), .Q(\registers[8] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[5__693 .GSR = "DISABLED";
    FD1S3AX \registers_8[[4__694  (.D(\registers[8] [8]), .CK(clk_c), .Q(\registers[8] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_8[[4__694 .GSR = "DISABLED";
    FD1S3AX \registers_9[[3__695  (.D(registers_9__3__N_1789), .CK(clk_c), 
            .Q(\registers[9] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[3__695 .GSR = "DISABLED";
    FD1S3AX \registers_9[[2__696  (.D(registers_9__2__N_1792), .CK(clk_c), 
            .Q(\registers[9] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[2__696 .GSR = "DISABLED";
    FD1S3AX \registers_9[[1__697  (.D(registers_9__1__N_1793), .CK(clk_c), 
            .Q(\registers[9] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[1__697 .GSR = "DISABLED";
    FD1S3AX \registers_9[[0__698  (.D(registers_9__0__N_1794), .CK(clk_c), 
            .Q(\registers[9] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_9[[0__698 .GSR = "DISABLED";
    FD1S3AX \registers_9[[31__699  (.D(\registers[9] [3]), .CK(clk_c), .Q(\registers[9] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[31__699 .GSR = "DISABLED";
    FD1S3AX \registers_9[[30__700  (.D(\registers[9] [2]), .CK(clk_c), .Q(\registers[9] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[30__700 .GSR = "DISABLED";
    FD1S3AX \registers_9[[29__701  (.D(\registers[9] [1]), .CK(clk_c), .Q(\registers[9] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[29__701 .GSR = "DISABLED";
    FD1S3AX \registers_9[[28__702  (.D(\registers[9] [0]), .CK(clk_c), .Q(\registers[9] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[28__702 .GSR = "DISABLED";
    FD1S3AX \registers_9[[27__703  (.D(\registers[9] [31]), .CK(clk_c), 
            .Q(\registers[9] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[27__703 .GSR = "DISABLED";
    FD1S3AX \registers_9[[26__704  (.D(\registers[9] [30]), .CK(clk_c), 
            .Q(\registers[9] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[26__704 .GSR = "DISABLED";
    FD1S3AX \registers_9[[25__705  (.D(\registers[9] [29]), .CK(clk_c), 
            .Q(\registers[9] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[25__705 .GSR = "DISABLED";
    FD1S3AX \registers_9[[24__706  (.D(\registers[9] [28]), .CK(clk_c), 
            .Q(\registers[9] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[24__706 .GSR = "DISABLED";
    FD1S3AX \registers_9[[23__707  (.D(\registers[9] [27]), .CK(clk_c), 
            .Q(\registers[9] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[23__707 .GSR = "DISABLED";
    FD1S3AX \registers_9[[22__708  (.D(\registers[9] [26]), .CK(clk_c), 
            .Q(\registers[9] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[22__708 .GSR = "DISABLED";
    FD1S3AX \registers_9[[21__709  (.D(\registers[9] [25]), .CK(clk_c), 
            .Q(\registers[9] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[21__709 .GSR = "DISABLED";
    FD1S3AX \registers_9[[20__710  (.D(\registers[9] [24]), .CK(clk_c), 
            .Q(\registers[9] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[20__710 .GSR = "DISABLED";
    FD1S3AX \registers_9[[19__711  (.D(\registers[9] [23]), .CK(clk_c), 
            .Q(\registers[9] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[19__711 .GSR = "DISABLED";
    FD1S3AX \registers_9[[18__712  (.D(\registers[9] [22]), .CK(clk_c), 
            .Q(\registers[9] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[18__712 .GSR = "DISABLED";
    FD1S3AX \registers_9[[17__713  (.D(\registers[9] [21]), .CK(clk_c), 
            .Q(\registers[9] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[17__713 .GSR = "DISABLED";
    FD1S3AX \registers_9[[16__714  (.D(\registers[9] [20]), .CK(clk_c), 
            .Q(\registers[9] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[16__714 .GSR = "DISABLED";
    FD1S3AX \registers_9[[15__715  (.D(\registers[9] [19]), .CK(clk_c), 
            .Q(\registers[9] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[15__715 .GSR = "DISABLED";
    FD1S3AX \registers_9[[14__716  (.D(\registers[9] [18]), .CK(clk_c), 
            .Q(\registers[9] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[14__716 .GSR = "DISABLED";
    FD1S3AX \registers_9[[13__717  (.D(\registers[9] [17]), .CK(clk_c), 
            .Q(\registers[9] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[13__717 .GSR = "DISABLED";
    FD1S3AX \registers_9[[12__718  (.D(\registers[9] [16]), .CK(clk_c), 
            .Q(\registers[9] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[12__718 .GSR = "DISABLED";
    FD1S3AX \registers_9[[11__719  (.D(\registers[9] [15]), .CK(clk_c), 
            .Q(\registers[9] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[11__719 .GSR = "DISABLED";
    FD1S3AX \registers_9[[10__720  (.D(\registers[9] [14]), .CK(clk_c), 
            .Q(\registers[9] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[10__720 .GSR = "DISABLED";
    FD1S3AX \registers_9[[9__721  (.D(\registers[9] [13]), .CK(clk_c), .Q(\registers[9] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[9__721 .GSR = "DISABLED";
    FD1S3AX \registers_9[[8__722  (.D(\registers[9] [12]), .CK(clk_c), .Q(\registers[9] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[8__722 .GSR = "DISABLED";
    FD1S3AX \registers_9[[7__723  (.D(\registers[9] [11]), .CK(clk_c), .Q(\registers[9] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[7__723 .GSR = "DISABLED";
    FD1S3AX \registers_9[[6__724  (.D(\registers[9] [10]), .CK(clk_c), .Q(\registers[9] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[6__724 .GSR = "DISABLED";
    FD1S3AX \registers_9[[5__725  (.D(\registers[9] [9]), .CK(clk_c), .Q(\registers[9] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[5__725 .GSR = "DISABLED";
    FD1S3AX \registers_9[[4__726  (.D(\registers[9] [8]), .CK(clk_c), .Q(\registers[9] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_9[[4__726 .GSR = "DISABLED";
    FD1S3AX \registers_10[[3__727  (.D(registers_10__3__N_1795), .CK(clk_c), 
            .Q(\registers[10] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[3__727 .GSR = "DISABLED";
    FD1S3AX \registers_10[[2__728  (.D(registers_10__2__N_1798), .CK(clk_c), 
            .Q(\registers[10] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[2__728 .GSR = "DISABLED";
    FD1S3AX \registers_10[[1__729  (.D(registers_10__1__N_1799), .CK(clk_c), 
            .Q(\registers[10] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[1__729 .GSR = "DISABLED";
    FD1S3AX \registers_10[[0__730  (.D(registers_10__0__N_1800), .CK(clk_c), 
            .Q(\registers[10] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_10[[0__730 .GSR = "DISABLED";
    FD1S3AX \registers_10[[31__731  (.D(\registers[10] [3]), .CK(clk_c), 
            .Q(\registers[10] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[31__731 .GSR = "DISABLED";
    FD1S3AX \registers_10[[30__732  (.D(\registers[10] [2]), .CK(clk_c), 
            .Q(\registers[10] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[30__732 .GSR = "DISABLED";
    FD1S3AX \registers_10[[29__733  (.D(\registers[10] [1]), .CK(clk_c), 
            .Q(\registers[10] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[29__733 .GSR = "DISABLED";
    FD1S3AX \registers_10[[28__734  (.D(\registers[10] [0]), .CK(clk_c), 
            .Q(\registers[10] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[28__734 .GSR = "DISABLED";
    FD1S3AX \registers_10[[27__735  (.D(\registers[10] [31]), .CK(clk_c), 
            .Q(\registers[10] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[27__735 .GSR = "DISABLED";
    FD1S3AX \registers_10[[26__736  (.D(\registers[10] [30]), .CK(clk_c), 
            .Q(\registers[10] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[26__736 .GSR = "DISABLED";
    FD1S3AX \registers_10[[25__737  (.D(\registers[10] [29]), .CK(clk_c), 
            .Q(\registers[10] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[25__737 .GSR = "DISABLED";
    FD1S3AX \registers_10[[24__738  (.D(\registers[10] [28]), .CK(clk_c), 
            .Q(\registers[10] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[24__738 .GSR = "DISABLED";
    FD1S3AX \registers_10[[23__739  (.D(\registers[10] [27]), .CK(clk_c), 
            .Q(\registers[10] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[23__739 .GSR = "DISABLED";
    FD1S3AX \registers_10[[22__740  (.D(\registers[10] [26]), .CK(clk_c), 
            .Q(\registers[10] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[22__740 .GSR = "DISABLED";
    FD1S3AX \registers_10[[21__741  (.D(\registers[10] [25]), .CK(clk_c), 
            .Q(\registers[10] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[21__741 .GSR = "DISABLED";
    FD1S3AX \registers_10[[20__742  (.D(\registers[10] [24]), .CK(clk_c), 
            .Q(\registers[10] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[20__742 .GSR = "DISABLED";
    FD1S3AX \registers_10[[19__743  (.D(\registers[10] [23]), .CK(clk_c), 
            .Q(\registers[10] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[19__743 .GSR = "DISABLED";
    FD1S3AX \registers_10[[18__744  (.D(\registers[10] [22]), .CK(clk_c), 
            .Q(\registers[10] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[18__744 .GSR = "DISABLED";
    FD1S3AX \registers_10[[17__745  (.D(\registers[10] [21]), .CK(clk_c), 
            .Q(\registers[10] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[17__745 .GSR = "DISABLED";
    FD1S3AX \registers_10[[16__746  (.D(\registers[10] [20]), .CK(clk_c), 
            .Q(\registers[10] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[16__746 .GSR = "DISABLED";
    FD1S3AX \registers_10[[15__747  (.D(\registers[10] [19]), .CK(clk_c), 
            .Q(\registers[10] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[15__747 .GSR = "DISABLED";
    FD1S3AX \registers_10[[14__748  (.D(\registers[10] [18]), .CK(clk_c), 
            .Q(\registers[10] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[14__748 .GSR = "DISABLED";
    FD1S3AX \registers_10[[13__749  (.D(\registers[10] [17]), .CK(clk_c), 
            .Q(\registers[10] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[13__749 .GSR = "DISABLED";
    FD1S3AX \registers_10[[12__750  (.D(\registers[10] [16]), .CK(clk_c), 
            .Q(\registers[10] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[12__750 .GSR = "DISABLED";
    FD1S3AX \registers_10[[11__751  (.D(\registers[10] [15]), .CK(clk_c), 
            .Q(\registers[10] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[11__751 .GSR = "DISABLED";
    FD1S3AX \registers_10[[10__752  (.D(\registers[10] [14]), .CK(clk_c), 
            .Q(\registers[10] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[10__752 .GSR = "DISABLED";
    FD1S3AX \registers_10[[9__753  (.D(\registers[10] [13]), .CK(clk_c), 
            .Q(\registers[10] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[9__753 .GSR = "DISABLED";
    FD1S3AX \registers_10[[8__754  (.D(\registers[10] [12]), .CK(clk_c), 
            .Q(\registers[10] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[8__754 .GSR = "DISABLED";
    FD1S3AX \registers_10[[7__755  (.D(\registers[10] [11]), .CK(clk_c), 
            .Q(\registers[10] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[7__755 .GSR = "DISABLED";
    FD1S3AX \registers_10[[6__756  (.D(\registers[10] [10]), .CK(clk_c), 
            .Q(\registers[10] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[6__756 .GSR = "DISABLED";
    FD1S3AX \registers_10[[5__757  (.D(\registers[10] [9]), .CK(clk_c), 
            .Q(\registers[10] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[5__757 .GSR = "DISABLED";
    FD1S3AX \registers_10[[4__758  (.D(\registers[10] [8]), .CK(clk_c), 
            .Q(\registers[10] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_10[[4__758 .GSR = "DISABLED";
    FD1S3AX \registers_11[[3__759  (.D(registers_11__3__N_1801), .CK(clk_c), 
            .Q(\registers[11] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[3__759 .GSR = "DISABLED";
    FD1S3AX \registers_11[[2__760  (.D(registers_11__2__N_1804), .CK(clk_c), 
            .Q(\registers[11] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[2__760 .GSR = "DISABLED";
    FD1S3AX \registers_11[[1__761  (.D(registers_11__1__N_1805), .CK(clk_c), 
            .Q(\registers[11] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[1__761 .GSR = "DISABLED";
    FD1S3AX \registers_11[[0__762  (.D(registers_11__0__N_1806), .CK(clk_c), 
            .Q(\registers[11] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_11[[0__762 .GSR = "DISABLED";
    FD1S3AX \registers_11[[31__763  (.D(\registers[11] [3]), .CK(clk_c), 
            .Q(\registers[11] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[31__763 .GSR = "DISABLED";
    FD1S3AX \registers_11[[30__764  (.D(\registers[11] [2]), .CK(clk_c), 
            .Q(\registers[11] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[30__764 .GSR = "DISABLED";
    FD1S3AX \registers_11[[29__765  (.D(\registers[11] [1]), .CK(clk_c), 
            .Q(\registers[11] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[29__765 .GSR = "DISABLED";
    FD1S3AX \registers_11[[28__766  (.D(\registers[11] [0]), .CK(clk_c), 
            .Q(\registers[11] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[28__766 .GSR = "DISABLED";
    FD1S3AX \registers_11[[27__767  (.D(\registers[11] [31]), .CK(clk_c), 
            .Q(\registers[11] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[27__767 .GSR = "DISABLED";
    FD1S3AX \registers_11[[26__768  (.D(\registers[11] [30]), .CK(clk_c), 
            .Q(\registers[11] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[26__768 .GSR = "DISABLED";
    FD1S3AX \registers_11[[25__769  (.D(\registers[11] [29]), .CK(clk_c), 
            .Q(\registers[11] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[25__769 .GSR = "DISABLED";
    FD1S3AX \registers_11[[24__770  (.D(\registers[11] [28]), .CK(clk_c), 
            .Q(\registers[11] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[24__770 .GSR = "DISABLED";
    FD1S3AX \registers_11[[23__771  (.D(\registers[11] [27]), .CK(clk_c), 
            .Q(\registers[11] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[23__771 .GSR = "DISABLED";
    FD1S3AX \registers_11[[22__772  (.D(\registers[11] [26]), .CK(clk_c), 
            .Q(\registers[11] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[22__772 .GSR = "DISABLED";
    FD1S3AX \registers_11[[21__773  (.D(\registers[11] [25]), .CK(clk_c), 
            .Q(\registers[11] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[21__773 .GSR = "DISABLED";
    FD1S3AX \registers_11[[20__774  (.D(\registers[11] [24]), .CK(clk_c), 
            .Q(\registers[11] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[20__774 .GSR = "DISABLED";
    FD1S3AX \registers_11[[19__775  (.D(\registers[11] [23]), .CK(clk_c), 
            .Q(\registers[11] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[19__775 .GSR = "DISABLED";
    FD1S3AX \registers_11[[18__776  (.D(\registers[11] [22]), .CK(clk_c), 
            .Q(\registers[11] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[18__776 .GSR = "DISABLED";
    FD1S3AX \registers_11[[17__777  (.D(\registers[11] [21]), .CK(clk_c), 
            .Q(\registers[11] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[17__777 .GSR = "DISABLED";
    FD1S3AX \registers_11[[16__778  (.D(\registers[11] [20]), .CK(clk_c), 
            .Q(\registers[11] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[16__778 .GSR = "DISABLED";
    FD1S3AX \registers_11[[15__779  (.D(\registers[11] [19]), .CK(clk_c), 
            .Q(\registers[11] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[15__779 .GSR = "DISABLED";
    FD1S3AX \registers_11[[14__780  (.D(\registers[11] [18]), .CK(clk_c), 
            .Q(\registers[11] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[14__780 .GSR = "DISABLED";
    FD1S3AX \registers_11[[13__781  (.D(\registers[11] [17]), .CK(clk_c), 
            .Q(\registers[11] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[13__781 .GSR = "DISABLED";
    FD1S3AX \registers_11[[12__782  (.D(\registers[11] [16]), .CK(clk_c), 
            .Q(\registers[11] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[12__782 .GSR = "DISABLED";
    FD1S3AX \registers_11[[11__783  (.D(\registers[11] [15]), .CK(clk_c), 
            .Q(\registers[11] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[11__783 .GSR = "DISABLED";
    FD1S3AX \registers_11[[10__784  (.D(\registers[11] [14]), .CK(clk_c), 
            .Q(\registers[11] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[10__784 .GSR = "DISABLED";
    FD1S3AX \registers_11[[9__785  (.D(\registers[11] [13]), .CK(clk_c), 
            .Q(\registers[11] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[9__785 .GSR = "DISABLED";
    FD1S3AX \registers_11[[8__786  (.D(\registers[11] [12]), .CK(clk_c), 
            .Q(\registers[11] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[8__786 .GSR = "DISABLED";
    FD1S3AX \registers_11[[7__787  (.D(\registers[11] [11]), .CK(clk_c), 
            .Q(\registers[11] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[7__787 .GSR = "DISABLED";
    FD1S3AX \registers_11[[6__788  (.D(\registers[11] [10]), .CK(clk_c), 
            .Q(\registers[11] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[6__788 .GSR = "DISABLED";
    FD1S3AX \registers_11[[5__789  (.D(\registers[11] [9]), .CK(clk_c), 
            .Q(\registers[11] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[5__789 .GSR = "DISABLED";
    FD1S3AX \registers_11[[4__790  (.D(\registers[11] [8]), .CK(clk_c), 
            .Q(\registers[11] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_11[[4__790 .GSR = "DISABLED";
    FD1S3AX \registers_12[[3__791  (.D(registers_12__3__N_1807), .CK(clk_c), 
            .Q(\registers[12] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[3__791 .GSR = "DISABLED";
    FD1S3AX \registers_12[[2__792  (.D(registers_12__2__N_1810), .CK(clk_c), 
            .Q(\registers[12] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[2__792 .GSR = "DISABLED";
    FD1S3AX \registers_12[[1__793  (.D(registers_12__1__N_1811), .CK(clk_c), 
            .Q(\registers[12] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[1__793 .GSR = "DISABLED";
    FD1S3AX \registers_12[[0__794  (.D(registers_12__0__N_1812), .CK(clk_c), 
            .Q(\registers[12] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_12[[0__794 .GSR = "DISABLED";
    FD1S3AX \registers_12[[31__795  (.D(\registers[12] [3]), .CK(clk_c), 
            .Q(\registers[12] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[31__795 .GSR = "DISABLED";
    FD1S3AX \registers_12[[30__796  (.D(\registers[12] [2]), .CK(clk_c), 
            .Q(\registers[12] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[30__796 .GSR = "DISABLED";
    FD1S3AX \registers_12[[29__797  (.D(\registers[12] [1]), .CK(clk_c), 
            .Q(\registers[12] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[29__797 .GSR = "DISABLED";
    FD1S3AX \registers_12[[28__798  (.D(\registers[12] [0]), .CK(clk_c), 
            .Q(\registers[12] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[28__798 .GSR = "DISABLED";
    FD1S3AX \registers_12[[27__799  (.D(\registers[12] [31]), .CK(clk_c), 
            .Q(\registers[12] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[27__799 .GSR = "DISABLED";
    FD1S3AX \registers_12[[26__800  (.D(\registers[12] [30]), .CK(clk_c), 
            .Q(\registers[12] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[26__800 .GSR = "DISABLED";
    FD1S3AX \registers_12[[25__801  (.D(\registers[12] [29]), .CK(clk_c), 
            .Q(\registers[12] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[25__801 .GSR = "DISABLED";
    FD1S3AX \registers_12[[24__802  (.D(\registers[12] [28]), .CK(clk_c), 
            .Q(\registers[12] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[24__802 .GSR = "DISABLED";
    FD1S3AX \registers_12[[23__803  (.D(\registers[12] [27]), .CK(clk_c), 
            .Q(\registers[12] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[23__803 .GSR = "DISABLED";
    FD1S3AX \registers_12[[22__804  (.D(\registers[12] [26]), .CK(clk_c), 
            .Q(\registers[12] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[22__804 .GSR = "DISABLED";
    FD1S3AX \registers_12[[21__805  (.D(\registers[12] [25]), .CK(clk_c), 
            .Q(\registers[12] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[21__805 .GSR = "DISABLED";
    FD1S3AX \registers_12[[20__806  (.D(\registers[12] [24]), .CK(clk_c), 
            .Q(\registers[12] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[20__806 .GSR = "DISABLED";
    FD1S3AX \registers_12[[19__807  (.D(\registers[12] [23]), .CK(clk_c), 
            .Q(\registers[12] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[19__807 .GSR = "DISABLED";
    FD1S3AX \registers_12[[18__808  (.D(\registers[12] [22]), .CK(clk_c), 
            .Q(\registers[12] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[18__808 .GSR = "DISABLED";
    FD1S3AX \registers_12[[17__809  (.D(\registers[12] [21]), .CK(clk_c), 
            .Q(\registers[12] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[17__809 .GSR = "DISABLED";
    FD1S3AX \registers_12[[16__810  (.D(\registers[12] [20]), .CK(clk_c), 
            .Q(\registers[12] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[16__810 .GSR = "DISABLED";
    FD1S3AX \registers_12[[15__811  (.D(\registers[12] [19]), .CK(clk_c), 
            .Q(\registers[12] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[15__811 .GSR = "DISABLED";
    FD1S3AX \registers_12[[14__812  (.D(\registers[12] [18]), .CK(clk_c), 
            .Q(\registers[12] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[14__812 .GSR = "DISABLED";
    FD1S3AX \registers_12[[13__813  (.D(\registers[12] [17]), .CK(clk_c), 
            .Q(\registers[12] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[13__813 .GSR = "DISABLED";
    FD1S3AX \registers_12[[12__814  (.D(\registers[12] [16]), .CK(clk_c), 
            .Q(\registers[12] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[12__814 .GSR = "DISABLED";
    FD1S3AX \registers_12[[11__815  (.D(\registers[12] [15]), .CK(clk_c), 
            .Q(\registers[12] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[11__815 .GSR = "DISABLED";
    FD1S3AX \registers_12[[10__816  (.D(\registers[12] [14]), .CK(clk_c), 
            .Q(\registers[12] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[10__816 .GSR = "DISABLED";
    FD1S3AX \registers_12[[9__817  (.D(\registers[12] [13]), .CK(clk_c), 
            .Q(\registers[12] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[9__817 .GSR = "DISABLED";
    FD1S3AX \registers_12[[8__818  (.D(\registers[12] [12]), .CK(clk_c), 
            .Q(\registers[12] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[8__818 .GSR = "DISABLED";
    FD1S3AX \registers_12[[7__819  (.D(\registers[12] [11]), .CK(clk_c), 
            .Q(\registers[12] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[7__819 .GSR = "DISABLED";
    FD1S3AX \registers_12[[6__820  (.D(\registers[12] [10]), .CK(clk_c), 
            .Q(\registers[12] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[6__820 .GSR = "DISABLED";
    FD1S3AX \registers_12[[5__821  (.D(\registers[12] [9]), .CK(clk_c), 
            .Q(\registers[12] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[5__821 .GSR = "DISABLED";
    FD1S3AX \registers_12[[4__822  (.D(\registers[12] [8]), .CK(clk_c), 
            .Q(\registers[12] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_12[[4__822 .GSR = "DISABLED";
    FD1S3AX \registers_13[[3__823  (.D(registers_13__3__N_1813), .CK(clk_c), 
            .Q(\registers[13] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[3__823 .GSR = "DISABLED";
    FD1S3AX \registers_13[[2__824  (.D(registers_13__2__N_1816), .CK(clk_c), 
            .Q(\registers[13] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[2__824 .GSR = "DISABLED";
    FD1S3AX \registers_13[[1__825  (.D(registers_13__1__N_1817), .CK(clk_c), 
            .Q(\registers[13] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[1__825 .GSR = "DISABLED";
    FD1S3AX \registers_13[[0__826  (.D(registers_13__0__N_1818), .CK(clk_c), 
            .Q(\registers[13] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_13[[0__826 .GSR = "DISABLED";
    FD1S3AX \registers_13[[31__827  (.D(\registers[13] [3]), .CK(clk_c), 
            .Q(\registers[13] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[31__827 .GSR = "DISABLED";
    FD1S3AX \registers_13[[30__828  (.D(\registers[13] [2]), .CK(clk_c), 
            .Q(\registers[13] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[30__828 .GSR = "DISABLED";
    FD1S3AX \registers_13[[29__829  (.D(\registers[13] [1]), .CK(clk_c), 
            .Q(\registers[13] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[29__829 .GSR = "DISABLED";
    FD1S3AX \registers_13[[28__830  (.D(\registers[13] [0]), .CK(clk_c), 
            .Q(\registers[13] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[28__830 .GSR = "DISABLED";
    FD1S3AX \registers_13[[27__831  (.D(\registers[13] [31]), .CK(clk_c), 
            .Q(\registers[13] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[27__831 .GSR = "DISABLED";
    FD1S3AX \registers_13[[26__832  (.D(\registers[13] [30]), .CK(clk_c), 
            .Q(\registers[13] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[26__832 .GSR = "DISABLED";
    FD1S3AX \registers_13[[25__833  (.D(\registers[13] [29]), .CK(clk_c), 
            .Q(\registers[13] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[25__833 .GSR = "DISABLED";
    FD1S3AX \registers_13[[24__834  (.D(\registers[13] [28]), .CK(clk_c), 
            .Q(\registers[13] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[24__834 .GSR = "DISABLED";
    FD1S3AX \registers_13[[23__835  (.D(\registers[13] [27]), .CK(clk_c), 
            .Q(\registers[13] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[23__835 .GSR = "DISABLED";
    FD1S3AX \registers_13[[22__836  (.D(\registers[13] [26]), .CK(clk_c), 
            .Q(\registers[13] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[22__836 .GSR = "DISABLED";
    FD1S3AX \registers_13[[21__837  (.D(\registers[13] [25]), .CK(clk_c), 
            .Q(\registers[13] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[21__837 .GSR = "DISABLED";
    FD1S3AX \registers_13[[20__838  (.D(\registers[13] [24]), .CK(clk_c), 
            .Q(\registers[13] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[20__838 .GSR = "DISABLED";
    FD1S3AX \registers_13[[19__839  (.D(\registers[13] [23]), .CK(clk_c), 
            .Q(\registers[13] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[19__839 .GSR = "DISABLED";
    FD1S3AX \registers_13[[18__840  (.D(\registers[13] [22]), .CK(clk_c), 
            .Q(\registers[13] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[18__840 .GSR = "DISABLED";
    FD1S3AX \registers_13[[17__841  (.D(\registers[13] [21]), .CK(clk_c), 
            .Q(\registers[13] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[17__841 .GSR = "DISABLED";
    FD1S3AX \registers_13[[16__842  (.D(\registers[13] [20]), .CK(clk_c), 
            .Q(\registers[13] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[16__842 .GSR = "DISABLED";
    FD1S3AX \registers_13[[15__843  (.D(\registers[13] [19]), .CK(clk_c), 
            .Q(\registers[13] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[15__843 .GSR = "DISABLED";
    FD1S3AX \registers_13[[14__844  (.D(\registers[13] [18]), .CK(clk_c), 
            .Q(\registers[13] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[14__844 .GSR = "DISABLED";
    FD1S3AX \registers_13[[13__845  (.D(\registers[13] [17]), .CK(clk_c), 
            .Q(\registers[13] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[13__845 .GSR = "DISABLED";
    FD1S3AX \registers_13[[12__846  (.D(\registers[13] [16]), .CK(clk_c), 
            .Q(\registers[13] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[12__846 .GSR = "DISABLED";
    FD1S3AX \registers_13[[11__847  (.D(\registers[13] [15]), .CK(clk_c), 
            .Q(\registers[13] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[11__847 .GSR = "DISABLED";
    FD1S3AX \registers_13[[10__848  (.D(\registers[13] [14]), .CK(clk_c), 
            .Q(\registers[13] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[10__848 .GSR = "DISABLED";
    FD1S3AX \registers_13[[9__849  (.D(\registers[13] [13]), .CK(clk_c), 
            .Q(\registers[13] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[9__849 .GSR = "DISABLED";
    FD1S3AX \registers_13[[8__850  (.D(\registers[13] [12]), .CK(clk_c), 
            .Q(\registers[13] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[8__850 .GSR = "DISABLED";
    FD1S3AX \registers_13[[7__851  (.D(\registers[13] [11]), .CK(clk_c), 
            .Q(\registers[13] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[7__851 .GSR = "DISABLED";
    FD1S3AX \registers_13[[6__852  (.D(\registers[13] [10]), .CK(clk_c), 
            .Q(\registers[13] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[6__852 .GSR = "DISABLED";
    FD1S3AX \registers_13[[5__853  (.D(\registers[13] [9]), .CK(clk_c), 
            .Q(\registers[13] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[5__853 .GSR = "DISABLED";
    FD1S3AX \registers_13[[4__854  (.D(\registers[13] [8]), .CK(clk_c), 
            .Q(\registers[13] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_13[[4__854 .GSR = "DISABLED";
    FD1S3AX \registers_14[[3__855  (.D(registers_14__3__N_1819), .CK(clk_c), 
            .Q(\registers[14] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[3__855 .GSR = "DISABLED";
    FD1S3AX \registers_14[[2__856  (.D(registers_14__2__N_1822), .CK(clk_c), 
            .Q(\registers[14] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[2__856 .GSR = "DISABLED";
    FD1S3AX \registers_14[[1__857  (.D(registers_14__1__N_1823), .CK(clk_c), 
            .Q(\registers[14] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[1__857 .GSR = "DISABLED";
    FD1S3AX \registers_14[[0__858  (.D(registers_14__0__N_1824), .CK(clk_c), 
            .Q(\registers[14] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_14[[0__858 .GSR = "DISABLED";
    FD1S3AX \registers_14[[31__859  (.D(\registers[14] [3]), .CK(clk_c), 
            .Q(\registers[14] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[31__859 .GSR = "DISABLED";
    FD1S3AX \registers_14[[30__860  (.D(\registers[14] [2]), .CK(clk_c), 
            .Q(\registers[14] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[30__860 .GSR = "DISABLED";
    FD1S3AX \registers_14[[29__861  (.D(\registers[14] [1]), .CK(clk_c), 
            .Q(\registers[14] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[29__861 .GSR = "DISABLED";
    FD1S3AX \registers_14[[28__862  (.D(\registers[14] [0]), .CK(clk_c), 
            .Q(\registers[14] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[28__862 .GSR = "DISABLED";
    FD1S3AX \registers_14[[27__863  (.D(\registers[14] [31]), .CK(clk_c), 
            .Q(\registers[14] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[27__863 .GSR = "DISABLED";
    FD1S3AX \registers_14[[26__864  (.D(\registers[14] [30]), .CK(clk_c), 
            .Q(\registers[14] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[26__864 .GSR = "DISABLED";
    FD1S3AX \registers_14[[25__865  (.D(\registers[14] [29]), .CK(clk_c), 
            .Q(\registers[14] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[25__865 .GSR = "DISABLED";
    FD1S3AX \registers_14[[24__866  (.D(\registers[14] [28]), .CK(clk_c), 
            .Q(\registers[14] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[24__866 .GSR = "DISABLED";
    FD1S3AX \registers_14[[23__867  (.D(\registers[14] [27]), .CK(clk_c), 
            .Q(\registers[14] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[23__867 .GSR = "DISABLED";
    FD1S3AX \registers_14[[22__868  (.D(\registers[14] [26]), .CK(clk_c), 
            .Q(\registers[14] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[22__868 .GSR = "DISABLED";
    FD1S3AX \registers_14[[21__869  (.D(\registers[14] [25]), .CK(clk_c), 
            .Q(\registers[14] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[21__869 .GSR = "DISABLED";
    FD1S3AX \registers_14[[20__870  (.D(\registers[14] [24]), .CK(clk_c), 
            .Q(\registers[14] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[20__870 .GSR = "DISABLED";
    FD1S3AX \registers_14[[19__871  (.D(\registers[14] [23]), .CK(clk_c), 
            .Q(\registers[14] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[19__871 .GSR = "DISABLED";
    FD1S3AX \registers_14[[18__872  (.D(\registers[14] [22]), .CK(clk_c), 
            .Q(\registers[14] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[18__872 .GSR = "DISABLED";
    FD1S3AX \registers_14[[17__873  (.D(\registers[14] [21]), .CK(clk_c), 
            .Q(\registers[14] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[17__873 .GSR = "DISABLED";
    FD1S3AX \registers_14[[16__874  (.D(\registers[14] [20]), .CK(clk_c), 
            .Q(\registers[14] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[16__874 .GSR = "DISABLED";
    FD1S3AX \registers_14[[15__875  (.D(\registers[14] [19]), .CK(clk_c), 
            .Q(\registers[14] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[15__875 .GSR = "DISABLED";
    FD1S3AX \registers_14[[14__876  (.D(\registers[14] [18]), .CK(clk_c), 
            .Q(\registers[14] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[14__876 .GSR = "DISABLED";
    FD1S3AX \registers_14[[13__877  (.D(\registers[14] [17]), .CK(clk_c), 
            .Q(\registers[14] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[13__877 .GSR = "DISABLED";
    FD1S3AX \registers_14[[12__878  (.D(\registers[14] [16]), .CK(clk_c), 
            .Q(\registers[14] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[12__878 .GSR = "DISABLED";
    FD1S3AX \registers_14[[11__879  (.D(\registers[14] [15]), .CK(clk_c), 
            .Q(\registers[14] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[11__879 .GSR = "DISABLED";
    FD1S3AX \registers_14[[10__880  (.D(\registers[14] [14]), .CK(clk_c), 
            .Q(\registers[14] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[10__880 .GSR = "DISABLED";
    FD1S3AX \registers_14[[9__881  (.D(\registers[14] [13]), .CK(clk_c), 
            .Q(\registers[14] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[9__881 .GSR = "DISABLED";
    FD1S3AX \registers_14[[8__882  (.D(\registers[14] [12]), .CK(clk_c), 
            .Q(\registers[14] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[8__882 .GSR = "DISABLED";
    FD1S3AX \registers_14[[7__883  (.D(\registers[14] [11]), .CK(clk_c), 
            .Q(\registers[14] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[7__883 .GSR = "DISABLED";
    FD1S3AX \registers_14[[6__884  (.D(\registers[14] [10]), .CK(clk_c), 
            .Q(\registers[14] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[6__884 .GSR = "DISABLED";
    FD1S3AX \registers_14[[5__885  (.D(\registers[14] [9]), .CK(clk_c), 
            .Q(\registers[14] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[5__885 .GSR = "DISABLED";
    FD1S3AX \registers_14[[4__886  (.D(\registers[14] [8]), .CK(clk_c), 
            .Q(\registers[14] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_14[[4__886 .GSR = "DISABLED";
    FD1S3AX \registers_15[[3__887  (.D(registers_15__3__N_1825), .CK(clk_c), 
            .Q(\registers[15] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[3__887 .GSR = "DISABLED";
    FD1S3AX \registers_15[[2__888  (.D(registers_15__2__N_1828), .CK(clk_c), 
            .Q(\registers[15] [2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[2__888 .GSR = "DISABLED";
    FD1S3AX \registers_15[[1__889  (.D(registers_15__1__N_1829), .CK(clk_c), 
            .Q(\registers[15] [1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[1__889 .GSR = "DISABLED";
    FD1S3AX \registers_15[[0__890  (.D(registers_15__0__N_1830), .CK(clk_c), 
            .Q(\registers[15] [0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_15[[0__890 .GSR = "DISABLED";
    FD1S3AX \registers_15[[31__891  (.D(\registers[15] [3]), .CK(clk_c), 
            .Q(\registers[15] [31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[31__891 .GSR = "DISABLED";
    FD1S3AX \registers_15[[30__892  (.D(\registers[15] [2]), .CK(clk_c), 
            .Q(\registers[15] [30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[30__892 .GSR = "DISABLED";
    FD1S3AX \registers_15[[29__893  (.D(\registers[15] [1]), .CK(clk_c), 
            .Q(\registers[15] [29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[29__893 .GSR = "DISABLED";
    FD1S3AX \registers_15[[28__894  (.D(\registers[15] [0]), .CK(clk_c), 
            .Q(\registers[15] [28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[28__894 .GSR = "DISABLED";
    FD1S3AX \registers_15[[27__895  (.D(\registers[15] [31]), .CK(clk_c), 
            .Q(\registers[15] [27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[27__895 .GSR = "DISABLED";
    FD1S3AX \registers_15[[26__896  (.D(\registers[15] [30]), .CK(clk_c), 
            .Q(\registers[15] [26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[26__896 .GSR = "DISABLED";
    FD1S3AX \registers_15[[25__897  (.D(\registers[15] [29]), .CK(clk_c), 
            .Q(\registers[15] [25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[25__897 .GSR = "DISABLED";
    FD1S3AX \registers_15[[24__898  (.D(\registers[15] [28]), .CK(clk_c), 
            .Q(\registers[15] [24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[24__898 .GSR = "DISABLED";
    FD1S3AX \registers_15[[23__899  (.D(\registers[15] [27]), .CK(clk_c), 
            .Q(\registers[15] [23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[23__899 .GSR = "DISABLED";
    FD1S3AX \registers_15[[22__900  (.D(\registers[15] [26]), .CK(clk_c), 
            .Q(\registers[15] [22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[22__900 .GSR = "DISABLED";
    FD1S3AX \registers_15[[21__901  (.D(\registers[15] [25]), .CK(clk_c), 
            .Q(\registers[15] [21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[21__901 .GSR = "DISABLED";
    FD1S3AX \registers_15[[20__902  (.D(\registers[15] [24]), .CK(clk_c), 
            .Q(\registers[15] [20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[20__902 .GSR = "DISABLED";
    FD1S3AX \registers_15[[19__903  (.D(\registers[15] [23]), .CK(clk_c), 
            .Q(\registers[15] [19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[19__903 .GSR = "DISABLED";
    FD1S3AX \registers_15[[18__904  (.D(\registers[15] [22]), .CK(clk_c), 
            .Q(\registers[15] [18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[18__904 .GSR = "DISABLED";
    FD1S3AX \registers_15[[17__905  (.D(\registers[15] [21]), .CK(clk_c), 
            .Q(\registers[15] [17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[17__905 .GSR = "DISABLED";
    FD1S3AX \registers_15[[16__906  (.D(\registers[15] [20]), .CK(clk_c), 
            .Q(\registers[15] [16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[16__906 .GSR = "DISABLED";
    FD1S3AX \registers_15[[15__907  (.D(\registers[15] [19]), .CK(clk_c), 
            .Q(\registers[15] [15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[15__907 .GSR = "DISABLED";
    FD1S3AX \registers_15[[14__908  (.D(\registers[15] [18]), .CK(clk_c), 
            .Q(\registers[15] [14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[14__908 .GSR = "DISABLED";
    FD1S3AX \registers_15[[13__909  (.D(\registers[15] [17]), .CK(clk_c), 
            .Q(\registers[15] [13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[13__909 .GSR = "DISABLED";
    FD1S3AX \registers_15[[12__910  (.D(\registers[15] [16]), .CK(clk_c), 
            .Q(\registers[15] [12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[12__910 .GSR = "DISABLED";
    FD1S3AX \registers_15[[11__911  (.D(\registers[15] [15]), .CK(clk_c), 
            .Q(\registers[15] [11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[11__911 .GSR = "DISABLED";
    FD1S3AX \registers_15[[10__912  (.D(\registers[15] [14]), .CK(clk_c), 
            .Q(\registers[15] [10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[10__912 .GSR = "DISABLED";
    FD1S3AX \registers_15[[9__913  (.D(\registers[15] [13]), .CK(clk_c), 
            .Q(\registers[15] [9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[9__913 .GSR = "DISABLED";
    FD1S3AX \registers_15[[8__914  (.D(\registers[15] [12]), .CK(clk_c), 
            .Q(\registers[15] [8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[8__914 .GSR = "DISABLED";
    FD1S3AX \registers_15[[7__915  (.D(\registers[15] [11]), .CK(clk_c), 
            .Q(\registers[15] [7])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[7__915 .GSR = "DISABLED";
    FD1S3AX \registers_15[[6__916  (.D(\registers[15] [10]), .CK(clk_c), 
            .Q(\registers[15] [6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[6__916 .GSR = "DISABLED";
    FD1S3AX \registers_15[[5__917  (.D(\registers[15] [9]), .CK(clk_c), 
            .Q(\registers[15] [5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[5__917 .GSR = "DISABLED";
    FD1S3AX \registers_15[[4__918  (.D(\registers[15] [8]), .CK(clk_c), 
            .Q(\registers[15] [4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(64[24:69])
    defparam \registers_15[[4__918 .GSR = "DISABLED";
    FD1S3AX \registers_1[[3__503  (.D(registers_1__3__N_1753), .CK(clk_c), 
            .Q(\registers[1] [3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=9, LSE_RCOL=103, LSE_LLINE=91, LSE_RLINE=91 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(42[24] 47[20])
    defparam \registers_1[[3__503 .GSR = "DISABLED";
    LUT4 registers_15__7__I_0_3_lut_4_lut (.A(n31984), .B(n31750), .C(debug_rd[3]), 
         .D(\registers[15] [7]), .Z(registers_15__3__N_1825)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_543), .C(mstatus_mie), 
         .D(interrupt_pending_N_1671), .Z(n27480)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h2000;
    LUT4 registers_15__6__I_0_3_lut_4_lut (.A(n31984), .B(n31750), .C(debug_rd[2]), 
         .D(\registers[15] [6]), .Z(registers_15__2__N_1828)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_15__5__I_0_3_lut_4_lut (.A(n31984), .B(n31750), .C(debug_rd[1]), 
         .D(\registers[15] [5]), .Z(registers_15__1__N_1829)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 debug_branch_N_441_I_0_2_lut_rep_542_3_lut_4_lut (.A(counter_hi[2]), 
         .B(clk_c_enable_543), .C(was_early_branch), .D(n26597), .Z(n31747)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam debug_branch_N_441_I_0_2_lut_rep_542_3_lut_4_lut.init = 16'hfdff;
    LUT4 registers_15__4__I_0_3_lut_4_lut (.A(n31984), .B(n31750), .C(debug_rd[0]), 
         .D(\registers[15] [4]), .Z(registers_15__0__N_1830)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_15__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i27681_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_543), 
         .C(rst_reg_n), .D(n18086), .Z(clk_c_enable_348)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;
    defparam i27681_2_lut_3_lut_4_lut.init = 16'h2f0f;
    LUT4 i1_3_lut_4_lut_adj_275 (.A(counter_hi[2]), .B(clk_c_enable_543), 
         .C(mstatus_mie), .D(no_write_in_progress), .Z(n27534)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_275.init = 16'h2000;
    LUT4 registers_14__7__I_0_3_lut_4_lut (.A(n31984), .B(n31751), .C(debug_rd[3]), 
         .D(\registers[14] [7]), .Z(registers_14__3__N_1819)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 cycle_count_wide_6__I_0_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_543), 
         .C(time_hi[2]), .D(\cycle_count_wide[6] ), .Z(\time_count[3] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam cycle_count_wide_6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_14__6__I_0_3_lut_4_lut (.A(n31984), .B(n31751), .C(debug_rd[2]), 
         .D(\registers[14] [6]), .Z(registers_14__2__N_1822)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 cycle_count_wide_4__I_0_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_543), 
         .C(time_hi[0]), .D(\cycle_count_wide[4] ), .Z(\time_count[1] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam cycle_count_wide_4__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_14__5__I_0_3_lut_4_lut (.A(n31984), .B(n31751), .C(debug_rd[1]), 
         .D(\registers[14] [5]), .Z(registers_14__1__N_1823)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_543), 
         .C(n28150), .D(n26597), .Z(n27762)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hd0f0;
    LUT4 cycle_count_wide_5__I_0_3_lut_4_lut (.A(counter_hi[2]), .B(clk_c_enable_543), 
         .C(time_hi[1]), .D(\cycle_count_wide[5] ), .Z(\time_count[2] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam cycle_count_wide_5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_14__4__I_0_3_lut_4_lut (.A(n31984), .B(n31751), .C(debug_rd[0]), 
         .D(\registers[14] [4]), .Z(registers_14__0__N_1824)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_14__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__7__I_0_3_lut_4_lut (.A(n31984), .B(n31752), .C(debug_rd[3]), 
         .D(\registers[13] [7]), .Z(registers_13__3__N_1813)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__6__I_0_3_lut_4_lut (.A(n31984), .B(n31752), .C(debug_rd[2]), 
         .D(\registers[13] [6]), .Z(registers_13__2__N_1816)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_13__5__I_0_3_lut_4_lut (.A(n31984), .B(n31752), .C(debug_rd[1]), 
         .D(\registers[13] [5]), .Z(registers_13__1__N_1817)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_3_lut_4_lut_adj_276 (.A(counter_hi[2]), .B(clk_c_enable_543), 
         .C(n27018), .D(n26597), .Z(n28182)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (C))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_276.init = 16'h2f0f;
    LUT4 registers_13__4__I_0_3_lut_4_lut (.A(n31984), .B(n31752), .C(debug_rd[0]), 
         .D(\registers[13] [4]), .Z(registers_13__0__N_1818)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_13__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__7__I_0_3_lut_4_lut (.A(n31984), .B(n31749), .C(debug_rd[3]), 
         .D(\registers[12] [7]), .Z(registers_12__3__N_1807)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__7__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__6__I_0_3_lut_4_lut (.A(n31984), .B(n31749), .C(debug_rd[2]), 
         .D(\registers[12] [6]), .Z(registers_12__2__N_1810)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__6__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__5__I_0_3_lut_4_lut (.A(n31984), .B(n31749), .C(debug_rd[1]), 
         .D(\registers[12] [5]), .Z(registers_12__1__N_1811)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__5__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_12__4__I_0_3_lut_4_lut (.A(n31984), .B(n31749), .C(debug_rd[0]), 
         .D(\registers[12] [4]), .Z(registers_12__0__N_1812)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam registers_12__4__I_0_3_lut_4_lut.init = 16'hf780;
    LUT4 registers_11__7__I_0_3_lut_4_lut (.A(n31985), .B(n31750), .C(debug_rd[3]), 
         .D(\registers[11] [7]), .Z(registers_11__3__N_1801)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__6__I_0_3_lut_4_lut (.A(n31985), .B(n31750), .C(debug_rd[2]), 
         .D(\registers[11] [6]), .Z(registers_11__2__N_1804)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__5__I_0_3_lut_4_lut (.A(n31985), .B(n31750), .C(debug_rd[1]), 
         .D(\registers[11] [5]), .Z(registers_11__1__N_1805)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_11__4__I_0_3_lut_4_lut (.A(n31985), .B(n31750), .C(debug_rd[0]), 
         .D(\registers[11] [4]), .Z(registers_11__0__N_1806)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_11__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__7__I_0_3_lut_4_lut (.A(n31985), .B(n31751), .C(debug_rd[3]), 
         .D(\registers[10] [7]), .Z(registers_10__3__N_1795)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__6__I_0_3_lut_4_lut (.A(n31985), .B(n31751), .C(debug_rd[2]), 
         .D(\registers[10] [6]), .Z(registers_10__2__N_1798)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__5__I_0_3_lut_4_lut (.A(n31985), .B(n31751), .C(debug_rd[1]), 
         .D(\registers[10] [5]), .Z(registers_10__1__N_1799)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_10__4__I_0_3_lut_4_lut (.A(n31985), .B(n31751), .C(debug_rd[0]), 
         .D(\registers[10] [4]), .Z(registers_10__0__N_1800)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_10__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__7__I_0_3_lut_4_lut (.A(n31985), .B(n31752), .C(debug_rd[3]), 
         .D(\registers[9] [7]), .Z(registers_9__3__N_1789)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__6__I_0_3_lut_4_lut (.A(n31985), .B(n31752), .C(debug_rd[2]), 
         .D(\registers[9] [6]), .Z(registers_9__2__N_1792)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 i27144_4_lut_4_lut (.A(\registers[2] [5]), .B(rs2[0]), .C(rs2[1]), 
         .D(\registers[1] [5]), .Z(n29761)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i27144_4_lut_4_lut.init = 16'h2c20;
    LUT4 registers_9__5__I_0_3_lut_4_lut (.A(n31985), .B(n31752), .C(debug_rd[1]), 
         .D(\registers[9] [5]), .Z(registers_9__1__N_1793)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_9__4__I_0_3_lut_4_lut (.A(n31985), .B(n31752), .C(debug_rd[0]), 
         .D(\registers[9] [4]), .Z(registers_9__0__N_1794)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_9__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__7__I_0_3_lut_4_lut (.A(n31985), .B(n31749), .C(debug_rd[3]), 
         .D(\registers[8] [7]), .Z(registers_8__3__N_1783)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__6__I_0_3_lut_4_lut (.A(n31985), .B(n31749), .C(debug_rd[2]), 
         .D(\registers[8] [6]), .Z(registers_8__2__N_1786)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__5__I_0_3_lut_4_lut (.A(n31985), .B(n31749), .C(debug_rd[1]), 
         .D(\registers[8] [5]), .Z(registers_8__1__N_1787)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_8__4__I_0_3_lut_4_lut (.A(n31985), .B(n31749), .C(debug_rd[0]), 
         .D(\registers[8] [4]), .Z(registers_8__0__N_1788)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_8__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__7__I_0_3_lut_4_lut (.A(n31986), .B(n31750), .C(debug_rd[3]), 
         .D(\registers[7][7] ), .Z(registers_7__3__N_1777)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__6__I_0_3_lut_4_lut (.A(n31986), .B(n31750), .C(debug_rd[2]), 
         .D(\registers[7] [6]), .Z(registers_7__2__N_1780)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__5__I_0_3_lut_4_lut (.A(n31986), .B(n31750), .C(debug_rd[1]), 
         .D(\registers[7] [5]), .Z(registers_7__1__N_1781)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_7__4__I_0_3_lut_4_lut (.A(n31986), .B(n31750), .C(debug_rd[0]), 
         .D(\registers[7] [4]), .Z(registers_7__0__N_1782)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_7__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__7__I_0_3_lut_4_lut (.A(n31986), .B(n31751), .C(debug_rd[3]), 
         .D(\registers[6][7] ), .Z(registers_6__3__N_1771)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__6__I_0_3_lut_4_lut (.A(n31986), .B(n31751), .C(debug_rd[2]), 
         .D(\registers[6] [6]), .Z(registers_6__2__N_1774)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_6__5__I_0_3_lut_4_lut (.A(n31986), .B(n31751), .C(debug_rd[1]), 
         .D(\registers[6] [5]), .Z(registers_6__1__N_1775)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 i27050_3_lut (.A(\registers[2] [4]), .B(n15604), .C(rs1[0]), 
         .Z(n29667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27050_3_lut.init = 16'hcaca;
    LUT4 i27049_3_lut (.A(\registers[1] [4]), .B(rs1[0]), .Z(n29666)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27049_3_lut.init = 16'h8888;
    LUT4 registers_6__4__I_0_3_lut_4_lut (.A(n31986), .B(n31751), .C(debug_rd[0]), 
         .D(\registers[6] [4]), .Z(registers_6__0__N_1776)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_6__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__4__I_0_3_lut_4_lut (.A(n31986), .B(n31752), .C(debug_rd[0]), 
         .D(\registers[5] [4]), .Z(registers_5__0__N_1770)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__4__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__5__I_0_3_lut_4_lut (.A(n31986), .B(n31752), .C(debug_rd[1]), 
         .D(\registers[5] [5]), .Z(registers_5__1__N_1769)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__5__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__6__I_0_3_lut_4_lut (.A(n31986), .B(n31752), .C(debug_rd[2]), 
         .D(\registers[5] [6]), .Z(registers_5__2__N_1768)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__6__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_5__7__I_0_3_lut_4_lut (.A(n31986), .B(n31752), .C(debug_rd[3]), 
         .D(\registers[5][7] ), .Z(registers_5__3__N_1765)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam registers_5__7__I_0_3_lut_4_lut.init = 16'hfb40;
    LUT4 registers_2__6__I_0_3_lut_4_lut (.A(n31751), .B(n31989), .C(debug_rd[2]), 
         .D(\registers[2] [6]), .Z(registers_2__2__N_1762)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_2__4__I_0_3_lut_4_lut (.A(n31751), .B(n31989), .C(debug_rd[0]), 
         .D(\registers[2] [4]), .Z(registers_2__0__N_1764)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__4__I_0_3_lut_4_lut.init = 16'hfd20;
    PFUMX i27094 (.BLUT(n29703), .ALUT(n29704), .C0(rs1[1]), .Z(n29711));
    LUT4 registers_2__5__I_0_3_lut_4_lut (.A(n31751), .B(n31989), .C(debug_rd[1]), 
         .D(\registers[2] [5]), .Z(registers_2__1__N_1763)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 i15375_2_lut_rep_779 (.A(rd[2]), .B(rd[3]), .Z(n31984)) /* synthesis lut_function=(A (B)) */ ;
    defparam i15375_2_lut_rep_779.init = 16'h8888;
    LUT4 registers_2__7__I_0_3_lut_4_lut (.A(n31751), .B(n31989), .C(debug_rd[3]), 
         .D(\registers[2] [7]), .Z(registers_2__3__N_1759)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_2__7__I_0_3_lut_4_lut.init = 16'hfd20;
    PFUMX i27109 (.BLUT(n29718), .ALUT(n29719), .C0(rs2[1]), .Z(n29726));
    LUT4 registers_1__5__I_0_3_lut_4_lut (.A(n31752), .B(n31989), .C(debug_rd[1]), 
         .D(\registers[1] [5]), .Z(registers_1__1__N_1757)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__5__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 equal_147_i6_2_lut_rep_780 (.A(rd[2]), .B(rd[3]), .Z(n31985)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam equal_147_i6_2_lut_rep_780.init = 16'hbbbb;
    LUT4 registers_1__7__I_0_3_lut_4_lut (.A(n31752), .B(n31989), .C(debug_rd[3]), 
         .D(\registers[1] [7]), .Z(registers_1__3__N_1753)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__7__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 registers_1__4__I_0_3_lut_4_lut (.A(n31752), .B(n31989), .C(debug_rd[0]), 
         .D(\registers[1] [4]), .Z(registers_1__0__N_1758)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__4__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 equal_142_i6_2_lut_rep_781 (.A(rd[2]), .B(rd[3]), .Z(n31986)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(43[34:41])
    defparam equal_142_i6_2_lut_rep_781.init = 16'hdddd;
    LUT4 registers_1__6__I_0_3_lut_4_lut (.A(n31752), .B(n31989), .C(debug_rd[2]), 
         .D(\registers[1] [6]), .Z(registers_1__2__N_1756)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;
    defparam registers_1__6__I_0_3_lut_4_lut.init = 16'hfd20;
    LUT4 i15852_2_lut_rep_784 (.A(rd[3]), .B(rd[2]), .Z(n31989)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i15852_2_lut_rep_784.init = 16'heeee;
    PFUMX i27148 (.BLUT(n29761), .ALUT(n29762), .C0(rs2[2]), .Z(n29765));
    L6MUX21 i27149 (.D0(n29763), .D1(n29764), .SD(rs2[2]), .Z(n29766));
    PFUMX i27155 (.BLUT(n29768), .ALUT(n29769), .C0(rs1[2]), .Z(n29772));
    L6MUX21 i27156 (.D0(n29770), .D1(n29771), .SD(rs1[2]), .Z(n29773));
    LUT4 rs1_3__I_0_Mux_1_i12_3_lut (.A(\registers[14] [5]), .B(\registers[15] [5]), 
         .C(rs1[0]), .Z(n12_adj_3095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i12_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i11_3_lut (.A(\registers[12] [5]), .B(\registers[13] [5]), 
         .C(rs1[0]), .Z(n11_adj_3096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i11_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i9_3_lut (.A(\registers[10] [5]), .B(\registers[11] [5]), 
         .C(rs1[0]), .Z(n9_adj_3097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 i27130_4_lut_4_lut (.A(\registers[2] [7]), .B(rs2[0]), .C(rs2[1]), 
         .D(\registers[1] [7]), .Z(n29747)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i27130_4_lut_4_lut.init = 16'h2c20;
    LUT4 i27123_4_lut_4_lut (.A(\registers[2] [7]), .B(rs1[0]), .C(rs1[1]), 
         .D(\registers[1] [7]), .Z(n29740)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i27123_4_lut_4_lut.init = 16'h2c20;
    LUT4 rs1_3__I_0_Mux_1_i8_3_lut (.A(\registers[8] [5]), .B(\registers[9] [5]), 
         .C(rs1[0]), .Z(n8_adj_3098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i8_3_lut.init = 16'hcaca;
    LUT4 rs1_3__I_0_Mux_1_i5_3_lut (.A(\registers[6] [5]), .B(\registers[7] [5]), 
         .C(rs1[0]), .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i12_3_lut (.A(\registers[14] [5]), .B(\registers[15] [5]), 
         .C(rs2[0]), .Z(n12_adj_3099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i12_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i11_3_lut (.A(\registers[12] [5]), .B(\registers[13] [5]), 
         .C(rs2[0]), .Z(n11_adj_3100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i11_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i9_3_lut (.A(\registers[10] [5]), .B(\registers[11] [5]), 
         .C(rs2[0]), .Z(n9_adj_3101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i9_3_lut.init = 16'hcaca;
    LUT4 rs2_3__I_0_Mux_1_i8_3_lut (.A(\registers[8] [5]), .B(\registers[9] [5]), 
         .C(rs2[0]), .Z(n8_adj_3102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i8_3_lut.init = 16'hcaca;
    PFUMX i27028 (.BLUT(n29637), .ALUT(n29638), .C0(rs2[1]), .Z(n29645));
    LUT4 rs2_3__I_0_Mux_1_i5_3_lut (.A(\registers[6] [5]), .B(\registers[7] [5]), 
         .C(rs2[0]), .Z(n5_adj_3103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam rs2_3__I_0_Mux_1_i5_3_lut.init = 16'hcaca;
    LUT4 i27021_3_lut (.A(\registers[2] [4]), .B(n15604), .C(rs2[0]), 
         .Z(n29638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27021_3_lut.init = 16'hcaca;
    L6MUX21 i27033 (.D0(n29647), .D1(n29648), .SD(rs2[2]), .Z(n29650));
    L6MUX21 i27062 (.D0(n29676), .D1(n29677), .SD(rs1[2]), .Z(n29679));
    LUT4 i27020_3_lut (.A(\registers[1] [4]), .B(rs2[0]), .Z(n29637)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27020_3_lut.init = 16'h8888;
    L6MUX21 i27099 (.D0(n29713), .D1(n29714), .SD(rs1[2]), .Z(n29716));
    L6MUX21 i27114 (.D0(n29728), .D1(n29729), .SD(rs2[2]), .Z(n29731));
    L6MUX21 i27128 (.D0(n29742), .D1(n29743), .SD(rs1[2]), .Z(n29745));
    PFUMX i27146 (.BLUT(n8_adj_3102), .ALUT(n9_adj_3101), .C0(rs2[1]), 
          .Z(n29763));
    PFUMX i27147 (.BLUT(n11_adj_3100), .ALUT(n12_adj_3099), .C0(rs2[1]), 
          .Z(n29764));
    LUT4 i27250_3_lut_4_lut (.A(\registers[5] [5]), .B(rs2[0]), .C(rs2[1]), 
         .D(n5_adj_3103), .Z(n29762)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(72[34:37])
    defparam i27250_3_lut_4_lut.init = 16'hf808;
    PFUMX i27153 (.BLUT(n8_adj_3098), .ALUT(n9_adj_3097), .C0(rs1[1]), 
          .Z(n29770));
    LUT4 i27247_3_lut_4_lut (.A(\registers[5] [5]), .B(rs1[0]), .C(rs1[1]), 
         .D(n5), .Z(n29769)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i27247_3_lut_4_lut.init = 16'hf808;
    PFUMX i27154 (.BLUT(n11_adj_3096), .ALUT(n12_adj_3095), .C0(rs1[1]), 
          .Z(n29771));
    LUT4 rs1_3__I_0_Mux_3_i5_3_lut (.A(\registers[6][7] ), .B(\registers[7][7] ), 
         .C(rs1[0]), .Z(n5_adj_3104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam rs1_3__I_0_Mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 i27150_3_lut (.A(n29765), .B(n29766), .C(rs2[3]), .Z(\data_rs2[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27150_3_lut.init = 16'hcaca;
    LUT4 i27300_3_lut (.A(n4), .B(n5_adj_3104), .C(rs1[1]), .Z(n29741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27300_3_lut.init = 16'hcaca;
    LUT4 i27102_3_lut (.A(\registers[2] [6]), .B(\reg_access[3][2] ), .C(rs2[0]), 
         .Z(n29719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27102_3_lut.init = 16'hcaca;
    LUT4 i27101_3_lut (.A(\registers[1] [6]), .B(rs2[0]), .Z(n29718)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27101_3_lut.init = 16'h8888;
    LUT4 i27808_2_lut_rep_843 (.A(counter_hi[3]), .B(n33484), .Z(clk_c_enable_543)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i27808_2_lut_rep_843.init = 16'h7777;
    LUT4 i1_2_lut_3_lut_4_lut_adj_277 (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(\mcause[5] ), .D(counter_hi[2]), .Z(n28520)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_277.init = 16'h8000;
    LUT4 i23992_rep_126_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n26597), .D(counter_hi[2]), .Z(n30165)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i23992_rep_126_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23992_rep_127_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n26597), .D(counter_hi[2]), .Z(n30166)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i23992_rep_127_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23992_rep_130_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n26597), .D(counter_hi[2]), .Z(n30169)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i23992_rep_130_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23992_2_lut_rep_543_3_lut_4_lut (.A(n33486), .B(n33484), .C(n26597), 
         .D(counter_hi[2]), .Z(n31748)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i23992_2_lut_rep_543_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_712_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n32046), .D(counter_hi[2]), .Z(n31917)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_712_3_lut_4_lut.init = 16'h8000;
    LUT4 i23992_rep_128_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n26597), .D(counter_hi[2]), .Z(n30167)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i23992_rep_128_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_738_3_lut_4_lut (.A(n33486), .B(n33484), .C(n32046), 
         .D(counter_hi[2]), .Z(n31943)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_738_3_lut_4_lut.init = 16'h0800;
    PFUMX i27057 (.BLUT(n29666), .ALUT(n29667), .C0(rs1[1]), .Z(n29674));
    LUT4 i16084_2_lut_rep_769_3_lut (.A(n33486), .B(n33484), .C(counter_hi[2]), 
         .Z(clk_c_enable_36)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i16084_2_lut_rep_769_3_lut.init = 16'h8080;
    LUT4 i15355_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), .C(\mepc[0] ), 
         .Z(\csr_read_3__N_1451[0] )) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i15355_2_lut_3_lut.init = 16'h7070;
    LUT4 i23992_rep_129_2_lut_3_lut_4_lut (.A(counter_hi[3]), .B(counter_hi[4]), 
         .C(n26597), .D(counter_hi[2]), .Z(n30168)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i23992_rep_129_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i27769_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), .C(rst_reg_n), 
         .Z(n11559)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam i27769_2_lut_3_lut.init = 16'h0707;
    LUT4 i1_2_lut_3_lut (.A(counter_hi[3]), .B(counter_hi[4]), .C(\imm[6] ), 
         .Z(n26121)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h7070;
    LUT4 csr_read_3__N_1447_3__bdd_3_lut_4_lut (.A(n33486), .B(n33484), 
         .C(\imm[6] ), .D(\mepc[3] ), .Z(n31171)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;
    defparam csr_read_3__N_1447_3__bdd_3_lut_4_lut.init = 16'h7000;
    LUT4 i27157_3_lut (.A(n29772), .B(n29773), .C(rs1[3]), .Z(data_rs1[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27157_3_lut.init = 16'hcaca;
    LUT4 i27129_3_lut (.A(n29744), .B(n29745), .C(rs1[3]), .Z(data_rs1[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27129_3_lut.init = 16'hcaca;
    LUT4 i27087_3_lut (.A(\registers[2] [6]), .B(\reg_access[3][2] ), .C(rs1[0]), 
         .Z(n29704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27087_3_lut.init = 16'hcaca;
    LUT4 i27086_3_lut (.A(\registers[1] [6]), .B(rs1[0]), .Z(n29703)) /* synthesis lut_function=(A (B)) */ ;
    defparam i27086_3_lut.init = 16'h8888;
    LUT4 i27151_4_lut_4_lut (.A(\registers[2] [5]), .B(rs1[0]), .C(rs1[1]), 
         .D(\registers[1] [5]), .Z(n29768)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(71[34:37])
    defparam i27151_4_lut_4_lut.init = 16'h2c20;
    LUT4 i27715_3_lut (.A(counter_hi[2]), .B(n33486), .C(n33484), .Z(\reg_access[3][2] )) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(38[47:61])
    defparam i27715_3_lut.init = 16'h0404;
    LUT4 i27656_3_lut (.A(n33484), .B(n33486), .C(counter_hi[2]), .Z(n15604)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/register.v(40[41:55])
    defparam i27656_3_lut.init = 16'h0808;
    PFUMX i27029 (.BLUT(n29639), .ALUT(n29640), .C0(rs2[1]), .Z(n29646));
    PFUMX i27030 (.BLUT(n29641), .ALUT(n29642), .C0(rs2[1]), .Z(n29647));
    PFUMX i27031 (.BLUT(n29643), .ALUT(n29644), .C0(rs2[1]), .Z(n29648));
    PFUMX i27058 (.BLUT(n29668), .ALUT(n29669), .C0(rs1[1]), .Z(n29675));
    LUT4 i27063_3_lut (.A(n29678), .B(n29679), .C(rs1[3]), .Z(data_rs1[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27063_3_lut.init = 16'hcaca;
    PFUMX i27059 (.BLUT(n29670), .ALUT(n29671), .C0(rs1[1]), .Z(n29676));
    PFUMX i27060 (.BLUT(n29672), .ALUT(n29673), .C0(rs1[1]), .Z(n29677));
    PFUMX i27095 (.BLUT(n29705), .ALUT(n29706), .C0(rs1[1]), .Z(n29712));
    L6MUX21 i27034 (.D0(n29649), .D1(n29650), .SD(rs2[3]), .Z(\data_rs2[0] ));
    PFUMX i27096 (.BLUT(n29707), .ALUT(n29708), .C0(rs1[1]), .Z(n29713));
    PFUMX i27097 (.BLUT(n29709), .ALUT(n29710), .C0(rs1[1]), .Z(n29714));
    PFUMX i27110 (.BLUT(n29720), .ALUT(n29721), .C0(rs2[1]), .Z(n29727));
    L6MUX21 i27100 (.D0(n29715), .D1(n29716), .SD(rs1[3]), .Z(data_rs1[2]));
    L6MUX21 i27115 (.D0(n29730), .D1(n29731), .SD(rs2[3]), .Z(\data_rs2[2] ));
    PFUMX i27111 (.BLUT(n29722), .ALUT(n29723), .C0(rs2[1]), .Z(n29728));
    LUT4 i27063_3_lut_rep_865 (.A(n29678), .B(n29679), .C(rs1[3]), .Z(n33494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i27063_3_lut_rep_865.init = 16'hcaca;
    PFUMX i27112 (.BLUT(n29724), .ALUT(n29725), .C0(rs2[1]), .Z(n29729));
    L6MUX21 i27032 (.D0(n29645), .D1(n29646), .SD(rs2[2]), .Z(n29649));
    L6MUX21 i27061 (.D0(n29674), .D1(n29675), .SD(rs1[2]), .Z(n29678));
    L6MUX21 i27098 (.D0(n29711), .D1(n29712), .SD(rs1[2]), .Z(n29715));
    L6MUX21 i27113 (.D0(n29726), .D1(n29727), .SD(rs2[2]), .Z(n29730));
    PFUMX i27127 (.BLUT(n29740), .ALUT(n29741), .C0(rs1[2]), .Z(n29744));
    PFUMX i27125 (.BLUT(n8_adj_3094), .ALUT(n9_adj_3093), .C0(rs1[1]), 
          .Z(n29742));
    PFUMX i27126 (.BLUT(n11_adj_3092), .ALUT(n12_adj_3091), .C0(rs1[1]), 
          .Z(n29743));
    
endmodule
//
// Verilog Description of module tinyqv_counter_U0
//

module tinyqv_counter_U0 (cy, clk_c, n31980, \increment_result_3__N_1925[0] , 
            instrret_count, n31873, n31890) /* synthesis syn_module_defined=1 */ ;
    output cy;
    input clk_c;
    input n31980;
    input \increment_result_3__N_1925[0] ;
    output [3:0]instrret_count;
    input n31873;
    input n31890;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [4:0]increment_result_3__N_1925;
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    
    FD1S3IX cy_51 (.D(increment_result_3__N_1925[4]), .CK(clk_c), .CD(n31980), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3IX register_2__48 (.D(increment_result_3__N_1925[2]), .CK(clk_c), 
            .CD(n31980), .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result_3__N_1925[1]), .CK(clk_c), 
            .CD(n31980), .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(\increment_result_3__N_1925[0] ), .CK(clk_c), 
            .CD(n31980), .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(register[10])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(register[9])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(register[8])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(instrret_count[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(register[10]), .CK(clk_c), .Q(instrret_count[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(register[9]), .CK(clk_c), .Q(instrret_count[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(register[8]), .CK(clk_c), .Q(instrret_count[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result_3__N_1925[3]), .CK(clk_c), 
            .CD(n31980), .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=307, LSE_RLINE=315 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 i4803_2_lut_3_lut_4_lut (.A(instrret_count[1]), .B(n31873), .C(instrret_count[3]), 
         .D(instrret_count[2]), .Z(increment_result_3__N_1925[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4803_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4805_2_lut_3_lut_4_lut (.A(instrret_count[1]), .B(n31873), .C(instrret_count[3]), 
         .D(instrret_count[2]), .Z(increment_result_3__N_1925[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4805_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4789_2_lut_3_lut (.A(instrret_count[0]), .B(n31890), .C(instrret_count[1]), 
         .Z(increment_result_3__N_1925[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4789_2_lut_3_lut.init = 16'h7878;
    LUT4 i4796_2_lut_3_lut_4_lut (.A(instrret_count[0]), .B(n31890), .C(instrret_count[2]), 
         .D(instrret_count[1]), .Z(increment_result_3__N_1925[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4796_2_lut_3_lut_4_lut.init = 16'h78f0;
    
endmodule
//
// Verilog Description of module \tinyqv_counter(OUTPUT_WIDTH=7) 
//

module \tinyqv_counter(OUTPUT_WIDTH=7)  (cy, clk_c, n31980, \increment_result_3__N_1911[0] , 
            cycle_count_wide, n31912, n31945, n31870, n31949) /* synthesis syn_module_defined=1 */ ;
    output cy;
    input clk_c;
    input n31980;
    input \increment_result_3__N_1911[0] ;
    output [6:0]cycle_count_wide;
    input n31912;
    input n31945;
    output n31870;
    input n31949;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    wire [4:0]increment_result_3__N_1911;
    wire [31:0]register;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(17[16:24])
    
    FD1S3IX cy_51 (.D(increment_result_3__N_1911[4]), .CK(clk_c), .CD(n31980), 
            .Q(cy)) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam cy_51.GSR = "DISABLED";
    FD1S3IX register_2__48 (.D(increment_result_3__N_1911[2]), .CK(clk_c), 
            .CD(n31980), .Q(register[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_2__48.GSR = "DISABLED";
    FD1S3IX register_1__49 (.D(increment_result_3__N_1911[1]), .CK(clk_c), 
            .CD(n31980), .Q(register[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_1__49.GSR = "DISABLED";
    FD1S3IX register_0__50 (.D(\increment_result_3__N_1911[0] ), .CK(clk_c), 
            .CD(n31980), .Q(register[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_0__50.GSR = "DISABLED";
    FD1S3AX register_31__52 (.D(register[3]), .CK(clk_c), .Q(register[31])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_31__52.GSR = "DISABLED";
    FD1S3AX register_30__53 (.D(register[2]), .CK(clk_c), .Q(register[30])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_30__53.GSR = "DISABLED";
    FD1S3AX register_29__54 (.D(register[1]), .CK(clk_c), .Q(register[29])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_29__54.GSR = "DISABLED";
    FD1S3AX register_28__55 (.D(register[0]), .CK(clk_c), .Q(register[28])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_28__55.GSR = "DISABLED";
    FD1S3AX register_27__56 (.D(register[31]), .CK(clk_c), .Q(register[27])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_27__56.GSR = "DISABLED";
    FD1S3AX register_26__57 (.D(register[30]), .CK(clk_c), .Q(register[26])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_26__57.GSR = "DISABLED";
    FD1S3AX register_25__58 (.D(register[29]), .CK(clk_c), .Q(register[25])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_25__58.GSR = "DISABLED";
    FD1S3AX register_24__59 (.D(register[28]), .CK(clk_c), .Q(register[24])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_24__59.GSR = "DISABLED";
    FD1S3AX register_23__60 (.D(register[27]), .CK(clk_c), .Q(register[23])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_23__60.GSR = "DISABLED";
    FD1S3AX register_22__61 (.D(register[26]), .CK(clk_c), .Q(register[22])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_22__61.GSR = "DISABLED";
    FD1S3AX register_21__62 (.D(register[25]), .CK(clk_c), .Q(register[21])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_21__62.GSR = "DISABLED";
    FD1S3AX register_20__63 (.D(register[24]), .CK(clk_c), .Q(register[20])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_20__63.GSR = "DISABLED";
    FD1S3AX register_19__64 (.D(register[23]), .CK(clk_c), .Q(register[19])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_19__64.GSR = "DISABLED";
    FD1S3AX register_18__65 (.D(register[22]), .CK(clk_c), .Q(register[18])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_18__65.GSR = "DISABLED";
    FD1S3AX register_17__66 (.D(register[21]), .CK(clk_c), .Q(register[17])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_17__66.GSR = "DISABLED";
    FD1S3AX register_16__67 (.D(register[20]), .CK(clk_c), .Q(register[16])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_16__67.GSR = "DISABLED";
    FD1S3AX register_15__68 (.D(register[19]), .CK(clk_c), .Q(register[15])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_15__68.GSR = "DISABLED";
    FD1S3AX register_14__69 (.D(register[18]), .CK(clk_c), .Q(register[14])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_14__69.GSR = "DISABLED";
    FD1S3AX register_13__70 (.D(register[17]), .CK(clk_c), .Q(register[13])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_13__70.GSR = "DISABLED";
    FD1S3AX register_12__71 (.D(register[16]), .CK(clk_c), .Q(register[12])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_12__71.GSR = "DISABLED";
    FD1S3AX register_11__72 (.D(register[15]), .CK(clk_c), .Q(register[11])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_11__72.GSR = "DISABLED";
    FD1S3AX register_10__73 (.D(register[14]), .CK(clk_c), .Q(cycle_count_wide[6])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_10__73.GSR = "DISABLED";
    FD1S3AX register_9__74 (.D(register[13]), .CK(clk_c), .Q(cycle_count_wide[5])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_9__74.GSR = "DISABLED";
    FD1S3AX register_8__75 (.D(register[12]), .CK(clk_c), .Q(cycle_count_wide[4])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_8__75.GSR = "DISABLED";
    FD1S3AX register_7__76 (.D(register[11]), .CK(clk_c), .Q(cycle_count_wide[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_7__76.GSR = "DISABLED";
    FD1S3AX register_6__77 (.D(cycle_count_wide[6]), .CK(clk_c), .Q(cycle_count_wide[2])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_6__77.GSR = "DISABLED";
    FD1S3AX register_5__78 (.D(cycle_count_wide[5]), .CK(clk_c), .Q(cycle_count_wide[1])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_5__78.GSR = "DISABLED";
    FD1S3AX register_4__79 (.D(cycle_count_wide[4]), .CK(clk_c), .Q(cycle_count_wide[0])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(45[12:53])
    defparam register_4__79.GSR = "DISABLED";
    FD1S3IX register_3__47 (.D(increment_result_3__N_1911[3]), .CK(clk_c), 
            .CD(n31980), .Q(register[3])) /* synthesis LSE_LINE_FILE_ID=5, LSE_LCOL=40, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=290 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(21[12] 28[8])
    defparam register_3__47.GSR = "DISABLED";
    LUT4 i4777_2_lut_3_lut_4_lut (.A(cycle_count_wide[1]), .B(n31912), .C(cycle_count_wide[3]), 
         .D(cycle_count_wide[2]), .Z(increment_result_3__N_1911[4])) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4777_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i4775_2_lut_3_lut_4_lut (.A(cycle_count_wide[1]), .B(n31912), .C(cycle_count_wide[3]), 
         .D(cycle_count_wide[2]), .Z(increment_result_3__N_1911[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4775_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4770_2_lut_rep_665_3_lut_4_lut (.A(cycle_count_wide[0]), .B(n31945), 
         .C(cycle_count_wide[2]), .D(cycle_count_wide[1]), .Z(n31870)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4770_2_lut_rep_665_3_lut_4_lut.init = 16'h8000;
    LUT4 i4768_2_lut_3_lut_4_lut (.A(cycle_count_wide[0]), .B(n31945), .C(cycle_count_wide[2]), 
         .D(cycle_count_wide[1]), .Z(increment_result_3__N_1911[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[59:119])
    defparam i4768_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i4761_2_lut_3_lut_4_lut (.A(cy), .B(n31949), .C(cycle_count_wide[1]), 
         .D(cycle_count_wide[0]), .Z(increment_result_3__N_1911[1])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/counter.v(20[93:118])
    defparam i4761_2_lut_3_lut_4_lut.init = 16'h4bf0;
    
endmodule
//
// Verilog Description of module tinyqv_alu
//

module tinyqv_alu (alu_a_in, n31826, n31827, n30868, n28436, alu_b_in, 
            \alu_op_in[2] , n31959, n31924, n31787, n31856, cy_out, 
            n27558, n4913, n31979, n30870, n31825, n31960, alu_out) /* synthesis syn_module_defined=1 */ ;
    input [3:0]alu_a_in;
    input n31826;
    input n31827;
    output n30868;
    input n28436;
    input [3:0]alu_b_in;
    input \alu_op_in[2] ;
    input n31959;
    input n31924;
    input n31787;
    input n31856;
    output cy_out;
    input n27558;
    input [3:0]n4913;
    input n31979;
    output n30870;
    input n31825;
    input n31960;
    output [3:0]alu_out;
    
    
    wire n33478, n31759, n33477, n31753, n30869, n6, n28891, n31788, 
        n31767, n28342, n28308, n28370, n31859;
    wire [3:0]n4923;
    
    wire n31756;
    wire [3:0]a_xor_b;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[16:23])
    
    wire cmp_res_N_1855;
    wire [3:0]n4932;
    
    LUT4 i5371_4_lut_rep_853 (.A(alu_a_in[2]), .B(n33478), .C(n31759), 
         .D(n31826), .Z(n33477)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i5371_4_lut_rep_853.init = 16'haaa8;
    LUT4 n7026_bdd_4_lut (.A(n31753), .B(n33477), .C(n31827), .D(alu_a_in[3]), 
         .Z(n30869)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+(D)))) */ ;
    defparam n7026_bdd_4_lut.init = 16'hf110;
    LUT4 alu_op_in_0__bdd_4_lut (.A(n31753), .B(n33477), .C(n31827), .D(alu_a_in[3]), 
         .Z(n30868)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C (D))))) */ ;
    defparam alu_op_in_0__bdd_4_lut.init = 16'h011f;
    LUT4 i4745_2_lut_3_lut_4_lut_4_lut (.A(alu_a_in[2]), .B(n33478), .C(n31759), 
         .D(n31826), .Z(n6)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4745_2_lut_3_lut_4_lut_4_lut.init = 16'hfea8;
    LUT4 i26333_4_lut (.A(alu_a_in[0]), .B(n28436), .C(alu_b_in[0]), .D(\alu_op_in[2] ), 
         .Z(n28891)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A !(B (C+!(D))+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam i26333_4_lut.init = 16'h5a66;
    LUT4 i5449_3_lut_rep_583_4_lut (.A(alu_b_in[0]), .B(n31959), .C(n31924), 
         .D(alu_a_in[0]), .Z(n31788)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i5449_3_lut_rep_583_4_lut.init = 16'hf600;
    LUT4 i4731_2_lut_rep_562_3_lut_3_lut_4_lut (.A(alu_b_in[0]), .B(n31959), 
         .C(n31924), .D(alu_a_in[0]), .Z(n31767)) /* synthesis lut_function=(A (B (C (D))+!B (C+(D)))+!A (B (C+(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i4731_2_lut_rep_562_3_lut_3_lut_4_lut.init = 16'hf660;
    LUT4 i1_2_lut_3_lut (.A(alu_b_in[2]), .B(n31959), .C(alu_a_in[2]), 
         .Z(n28342)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut.init = 16'h9696;
    LUT4 i1_2_lut_3_lut_adj_273 (.A(alu_b_in[3]), .B(n31959), .C(alu_a_in[3]), 
         .Z(n28308)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut_adj_273.init = 16'h9696;
    LUT4 i5412_4_lut_rep_854 (.A(alu_a_in[1]), .B(n31787), .C(n31788), 
         .D(n31856), .Z(n33478)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i5412_4_lut_rep_854.init = 16'haaa8;
    LUT4 mux_3042_i2_4_lut (.A(n28370), .B(n31859), .C(\alu_op_in[2] ), 
         .D(n31767), .Z(n4923[1])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_3042_i2_4_lut.init = 16'hc5ca;
    LUT4 i4738_2_lut_rep_551_3_lut_4_lut_4_lut (.A(alu_a_in[1]), .B(n31787), 
         .C(n31788), .D(n31856), .Z(n31756)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4738_2_lut_rep_551_3_lut_4_lut_4_lut.init = 16'hfea8;
    LUT4 mux_3042_i3_4_lut (.A(n28342), .B(a_xor_b[2]), .C(\alu_op_in[2] ), 
         .D(n31756), .Z(n4923[2])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_3042_i3_4_lut.init = 16'hc5ca;
    LUT4 i4752_4_lut_4_lut (.A(alu_a_in[3]), .B(n31753), .C(n33477), .D(n31827), 
         .Z(cy_out)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B (D)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4752_4_lut_4_lut.init = 16'hfea8;
    LUT4 a_3__I_0_29_i3_2_lut (.A(alu_a_in[2]), .B(alu_b_in[2]), .Z(a_xor_b[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i3_2_lut.init = 16'h6666;
    LUT4 a_3__I_0_29_i4_2_lut (.A(alu_a_in[3]), .B(alu_b_in[3]), .Z(a_xor_b[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i4_2_lut.init = 16'h6666;
    LUT4 a_3__I_0_29_i1_2_lut (.A(alu_a_in[0]), .B(alu_b_in[0]), .Z(a_xor_b[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i1_2_lut.init = 16'h6666;
    LUT4 mux_3042_i4_4_lut (.A(n28308), .B(a_xor_b[3]), .C(\alu_op_in[2] ), 
         .D(n6), .Z(n4923[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(42[9] 48[16])
    defparam mux_3042_i4_4_lut.init = 16'hc5ca;
    LUT4 i1_4_lut (.A(a_xor_b[2]), .B(a_xor_b[3]), .C(a_xor_b[0]), .D(n27558), 
         .Z(cmp_res_N_1855)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    LUT4 i4743_2_lut_rep_548_3_lut_4_lut (.A(n31856), .B(n31767), .C(n31826), 
         .D(n33478), .Z(n31753)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4743_2_lut_rep_548_3_lut_4_lut.init = 16'hf080;
    PFUMX mux_3047_i4 (.BLUT(n4923[3]), .ALUT(n4913[3]), .C0(n31979), 
          .Z(n4932[3]));
    LUT4 i1_2_lut_3_lut_adj_274 (.A(alu_b_in[1]), .B(n31959), .C(alu_a_in[1]), 
         .Z(n28370)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(37[35:60])
    defparam i1_2_lut_3_lut_adj_274.init = 16'h9696;
    PFUMX mux_3047_i3 (.BLUT(n4923[2]), .ALUT(n4913[2]), .C0(n31979), 
          .Z(n4932[2]));
    LUT4 a_3__I_0_29_i2_2_lut_rep_654 (.A(alu_a_in[1]), .B(alu_b_in[1]), 
         .Z(n31859)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(39[26:31])
    defparam a_3__I_0_29_i2_2_lut_rep_654.init = 16'h6666;
    PFUMX mux_3047_i2 (.BLUT(n4923[1]), .ALUT(n4913[1]), .C0(n31979), 
          .Z(n4932[1]));
    PFUMX mux_3047_i1 (.BLUT(n28891), .ALUT(n4913[0]), .C0(n31979), .Z(n4932[0]));
    PFUMX i28113 (.BLUT(cmp_res_N_1855), .ALUT(n30869), .C0(n31979), .Z(n30870));
    LUT4 i4736_2_lut_rep_554_3_lut_4_lut_4_lut (.A(alu_a_in[0]), .B(n31825), 
         .C(n31924), .D(n31856), .Z(n31759)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/alu.v(38[22:43])
    defparam i4736_2_lut_rep_554_3_lut_4_lut_4_lut.init = 16'he800;
    LUT4 i15408_2_lut_4_lut (.A(n31960), .B(\alu_op_in[2] ), .C(n31979), 
         .D(n4932[0]), .Z(alu_out[0])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i15408_2_lut_4_lut.init = 16'hc500;
    LUT4 i15698_2_lut_4_lut (.A(n31960), .B(\alu_op_in[2] ), .C(n31979), 
         .D(n4932[1]), .Z(alu_out[1])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i15698_2_lut_4_lut.init = 16'hc500;
    LUT4 i15700_2_lut_4_lut (.A(n31960), .B(\alu_op_in[2] ), .C(n31979), 
         .D(n4932[3]), .Z(alu_out[3])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i15700_2_lut_4_lut.init = 16'hc500;
    LUT4 i15699_2_lut_4_lut (.A(n31960), .B(\alu_op_in[2] ), .C(n31979), 
         .D(n4932[2]), .Z(alu_out[2])) /* synthesis lut_function=(A (B (C (D)))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i15699_2_lut_4_lut.init = 16'hc500;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module tqvp_uart_tx_U1
//

module tqvp_uart_tx_U1 (cycle_counter, clk_c, clk_c_enable_376, n6210, 
            n72, debug_uart_txd, clk_c_enable_445, fsm_state, n32013, 
            debug_uart_tx_start, n31828, n26116, rst_reg_n, \data_to_write[7] , 
            next_bit, clk_c_enable_534, n31961, \data_to_write[1] , 
            \data_to_write[2] , \data_to_write[3] , \data_to_write[0] , 
            \data_to_write[4] , \data_to_write[5] , \data_to_write[6] , 
            uart_txd_N_2974) /* synthesis syn_module_defined=1 */ ;
    output [12:0]cycle_counter;
    input clk_c;
    input clk_c_enable_376;
    input n6210;
    input [12:0]n72;
    output debug_uart_txd;
    input clk_c_enable_445;
    output [3:0]fsm_state;
    output n32013;
    input debug_uart_tx_start;
    output n31828;
    output n26116;
    input rst_reg_n;
    input \data_to_write[7] ;
    output next_bit;
    input clk_c_enable_534;
    output n31961;
    input \data_to_write[1] ;
    input \data_to_write[2] ;
    input \data_to_write[3] ;
    input \data_to_write[0] ;
    input \data_to_write[4] ;
    input \data_to_write[5] ;
    input \data_to_write[6] ;
    output uart_txd_N_2974;
    
    wire clk_c /* synthesis SET_AS_NETWORK=clk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/top.v(9[20:23])
    
    wire uart_txd_N_2972, clk_c_enable_44, n31829, n32096;
    wire [3:0]fsm_state_c;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(47[11:20])
    
    wire n26117, n9337, n30569, n30568;
    wire [3:0]n162;
    wire [7:0]data_to_send;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(39[24:36])
    wire [7:0]data_to_send_7__N_2944;
    
    wire n28836, n28832, n28830, n28820;
    
    FD1P3IX cycle_counter__i0 (.D(n72[0]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i0.GSR = "DISABLED";
    FD1S3JX txd_reg_46 (.D(uart_txd_N_2972), .CK(clk_c), .PD(clk_c_enable_445), 
            .Q(debug_uart_txd)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(123[8] 133[4])
    defparam txd_reg_46.GSR = "DISABLED";
    FD1P3IX fsm_state__i0 (.D(n32096), .SP(clk_c_enable_44), .CD(n31829), 
            .CK(clk_c), .Q(fsm_state[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i0.GSR = "DISABLED";
    LUT4 fsm_state_0__bdd_4_lut (.A(fsm_state[0]), .B(fsm_state_c[2]), .C(fsm_state_c[1]), 
         .D(fsm_state_c[3]), .Z(n32096)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;
    defparam fsm_state_0__bdd_4_lut.init = 16'h4555;
    LUT4 i201_2_lut_rep_623_3_lut (.A(fsm_state[0]), .B(n32013), .C(debug_uart_tx_start), 
         .Z(n31828)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i201_2_lut_rep_623_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_4_lut (.A(fsm_state[0]), .B(n32013), .C(n26116), 
         .D(debug_uart_tx_start), .Z(n26117)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i27737_3_lut_rep_624_4_lut (.A(fsm_state[0]), .B(n32013), .C(debug_uart_tx_start), 
         .D(rst_reg_n), .Z(n31829)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i27737_3_lut_rep_624_4_lut.init = 16'h01ff;
    LUT4 i6737_2_lut_3_lut_2_lut_3_lut (.A(fsm_state[0]), .B(n32013), .C(rst_reg_n), 
         .Z(n9337)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i6737_2_lut_3_lut_2_lut_3_lut.init = 16'h1f1f;
    LUT4 i1_2_lut (.A(rst_reg_n), .B(\data_to_write[7] ), .Z(n26116)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    FD1P3IX fsm_state__i3 (.D(n30569), .SP(next_bit), .CD(n9337), .CK(clk_c), 
            .Q(fsm_state_c[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i3.GSR = "DISABLED";
    FD1P3IX fsm_state__i2 (.D(n30568), .SP(next_bit), .CD(n9337), .CK(clk_c), 
            .Q(fsm_state_c[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i2.GSR = "DISABLED";
    FD1P3IX fsm_state__i1 (.D(n162[1]), .SP(next_bit), .CD(n9337), .CK(clk_c), 
            .Q(fsm_state_c[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(112[8] 118[4])
    defparam fsm_state__i1.GSR = "DISABLED";
    LUT4 fsm_state_2__bdd_3_lut (.A(fsm_state_c[2]), .B(fsm_state_c[1]), 
         .C(fsm_state[0]), .Z(n30568)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam fsm_state_2__bdd_3_lut.init = 16'h6a6a;
    FD1P3IX cycle_counter__i12 (.D(n72[12]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i12.GSR = "DISABLED";
    FD1P3IX cycle_counter__i11 (.D(n72[11]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i11.GSR = "DISABLED";
    FD1P3IX cycle_counter__i10 (.D(n72[10]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i10.GSR = "DISABLED";
    FD1P3IX cycle_counter__i9 (.D(n72[9]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i9.GSR = "DISABLED";
    FD1P3IX cycle_counter__i8 (.D(n72[8]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i8.GSR = "DISABLED";
    FD1P3IX cycle_counter__i7 (.D(n72[7]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i7.GSR = "DISABLED";
    FD1P3IX cycle_counter__i6 (.D(n72[6]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i6.GSR = "DISABLED";
    FD1P3IX cycle_counter__i5 (.D(n72[5]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i5.GSR = "DISABLED";
    FD1P3IX cycle_counter__i4 (.D(n72[4]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i4.GSR = "DISABLED";
    FD1P3IX cycle_counter__i3 (.D(n72[3]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i3.GSR = "DISABLED";
    FD1P3IX cycle_counter__i2 (.D(n72[2]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i2.GSR = "DISABLED";
    FD1P3IX cycle_counter__i1 (.D(n72[1]), .SP(clk_c_enable_376), .CD(n6210), 
            .CK(clk_c), .Q(cycle_counter[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(99[8] 107[4])
    defparam cycle_counter__i1.GSR = "DISABLED";
    FD1P3IX data_to_send__i1 (.D(data_to_send_7__N_2944[1]), .SP(clk_c_enable_534), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i1.GSR = "DISABLED";
    LUT4 mux_13_i2_3_lut_4_lut (.A(n31961), .B(debug_uart_tx_start), .C(\data_to_write[1] ), 
         .D(data_to_send[2]), .Z(data_to_send_7__N_2944[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i3_3_lut_4_lut (.A(n31961), .B(debug_uart_tx_start), .C(\data_to_write[2] ), 
         .D(data_to_send[3]), .Z(data_to_send_7__N_2944[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i4_3_lut_4_lut (.A(n31961), .B(debug_uart_tx_start), .C(\data_to_write[3] ), 
         .D(data_to_send[4]), .Z(data_to_send_7__N_2944[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i4_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i1_3_lut_4_lut (.A(n31961), .B(debug_uart_tx_start), .C(\data_to_write[0] ), 
         .D(data_to_send[1]), .Z(data_to_send_7__N_2944[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i5_3_lut_4_lut (.A(n31961), .B(debug_uart_tx_start), .C(\data_to_write[4] ), 
         .D(data_to_send[5]), .Z(data_to_send_7__N_2944[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i6_3_lut_4_lut (.A(n31961), .B(debug_uart_tx_start), .C(\data_to_write[5] ), 
         .D(data_to_send[6]), .Z(data_to_send_7__N_2944[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 mux_13_i7_3_lut_4_lut (.A(n31961), .B(debug_uart_tx_start), .C(\data_to_write[6] ), 
         .D(data_to_send[7]), .Z(data_to_send_7__N_2944[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(89[17:52])
    defparam mux_13_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_3_lut_4_lut_3_lut (.A(n31961), .B(rst_reg_n), .C(next_bit), 
         .Z(clk_c_enable_44)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'hf7f7;
    FD1P3IX data_to_send__i2 (.D(data_to_send_7__N_2944[2]), .SP(clk_c_enable_534), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i2.GSR = "DISABLED";
    FD1P3IX data_to_send__i3 (.D(data_to_send_7__N_2944[3]), .SP(clk_c_enable_534), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i3.GSR = "DISABLED";
    FD1P3IX data_to_send__i0 (.D(data_to_send_7__N_2944[0]), .SP(clk_c_enable_534), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i0.GSR = "DISABLED";
    FD1P3IX data_to_send__i4 (.D(data_to_send_7__N_2944[4]), .SP(clk_c_enable_534), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i4.GSR = "DISABLED";
    FD1P3IX data_to_send__i5 (.D(data_to_send_7__N_2944[5]), .SP(clk_c_enable_534), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i5.GSR = "DISABLED";
    LUT4 i15414_3_lut_3_lut_4_lut (.A(fsm_state_c[3]), .B(fsm_state_c[1]), 
         .C(fsm_state_c[2]), .D(fsm_state[0]), .Z(n162[1])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(D)))) */ ;
    defparam i15414_3_lut_3_lut_4_lut.init = 16'h33c4;
    LUT4 i1_3_lut_rep_808 (.A(fsm_state_c[1]), .B(fsm_state_c[2]), .C(fsm_state_c[3]), 
         .Z(n32013)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i1_3_lut_rep_808.init = 16'hfefe;
    LUT4 i1_2_lut_rep_756_4_lut (.A(fsm_state_c[1]), .B(fsm_state_c[2]), 
         .C(fsm_state_c[3]), .D(fsm_state[0]), .Z(n31961)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam i1_2_lut_rep_756_4_lut.init = 16'hfffe;
    LUT4 uart_txd_I_254_4_lut_3_lut (.A(fsm_state_c[1]), .B(fsm_state_c[2]), 
         .C(fsm_state_c[3]), .Z(uart_txd_N_2974)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(126[17:39])
    defparam uart_txd_I_254_4_lut_3_lut.init = 16'h1e1e;
    FD1P3IX data_to_send__i6 (.D(data_to_send_7__N_2944[6]), .SP(clk_c_enable_534), 
            .CD(clk_c_enable_445), .CK(clk_c), .Q(data_to_send[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i6.GSR = "DISABLED";
    FD1P3AX data_to_send__i7 (.D(n26117), .SP(clk_c_enable_534), .CK(clk_c), 
            .Q(data_to_send[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=228, LSE_RLINE=236 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(86[8] 94[4])
    defparam data_to_send__i7.GSR = "DISABLED";
    LUT4 i15226_4_lut (.A(data_to_send[0]), .B(fsm_state[0]), .C(uart_txd_N_2974), 
         .D(n32013), .Z(uart_txd_N_2972)) /* synthesis lut_function=(A ((D)+!B)+!A !(B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/uart_tx.v(128[14] 132[8])
    defparam i15226_4_lut.init = 16'haf23;
    LUT4 i1_4_lut (.A(n28836), .B(n28832), .C(n28830), .D(cycle_counter[1]), 
         .Z(next_bit)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut.init = 16'hfefc;
    LUT4 i1_2_lut_adj_269 (.A(cycle_counter[3]), .B(cycle_counter[2]), .Z(n28836)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_269.init = 16'h8888;
    LUT4 i1_4_lut_adj_270 (.A(cycle_counter[8]), .B(n28820), .C(cycle_counter[10]), 
         .D(cycle_counter[6]), .Z(n28832)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_270.init = 16'hfffe;
    LUT4 i1_4_lut_adj_271 (.A(cycle_counter[11]), .B(cycle_counter[12]), 
         .C(cycle_counter[5]), .D(cycle_counter[7]), .Z(n28830)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_271.init = 16'hfffe;
    LUT4 i1_2_lut_adj_272 (.A(cycle_counter[9]), .B(cycle_counter[4]), .Z(n28820)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_272.init = 16'heeee;
    LUT4 fsm_state_3__bdd_4_lut (.A(fsm_state_c[3]), .B(fsm_state_c[1]), 
         .C(fsm_state_c[2]), .D(fsm_state[0]), .Z(n30569)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A !(B (C (D))))) */ ;
    defparam fsm_state_3__bdd_4_lut.init = 16'h6aa2;
    
endmodule
//
// Verilog Description of module sim_qspi_pmod
//

module sim_qspi_pmod (\addr[2] , qspi_clk_N_56, qspi_data_in, spi_clk_pos_derived_59, 
            qspi_data_in_3__N_1, \addr[1] , VCC_net, \addr[14] , \addr_24__N_228[14] , 
            \addr[13] , \addr[12] , \addr[11] , \addr[10] , \addr[9] , 
            \addr[8] , \addr[7] , \addr[6] , \addr[5] , \addr[4] , 
            \addr[3] , qspi_ram_a_select, qspi_ram_b_select, \addr[0] , 
            \addr_24__N_228[0] , \writing_N_164[3] , GND_net, \addr_24__N_228[9] , 
            \addr_24__N_228[7] , \addr_24__N_228[8] , \addr_24__N_228[6] , 
            \addr_24__N_228[5] , \addr_24__N_228[4] , \addr_24__N_228[3] , 
            \addr_24__N_228[2] , \addr_24__N_228[10] , \addr_24__N_228[11] , 
            \addr_24__N_228[12] , \addr_24__N_228[13] , \addr_24__N_228[1] , 
            n32031) /* synthesis syn_module_defined=1 */ ;
    output \addr[2] ;
    input qspi_clk_N_56;
    output [3:0]qspi_data_in;
    input spi_clk_pos_derived_59;
    input [3:0]qspi_data_in_3__N_1;
    output \addr[1] ;
    input VCC_net;
    output \addr[14] ;
    input \addr_24__N_228[14] ;
    output \addr[13] ;
    output \addr[12] ;
    output \addr[11] ;
    output \addr[10] ;
    output \addr[9] ;
    output \addr[8] ;
    output \addr[7] ;
    output \addr[6] ;
    output \addr[5] ;
    output \addr[4] ;
    output \addr[3] ;
    input qspi_ram_a_select;
    input qspi_ram_b_select;
    output \addr[0] ;
    input \addr_24__N_228[0] ;
    input \writing_N_164[3] ;
    input GND_net;
    input \addr_24__N_228[9] ;
    input \addr_24__N_228[7] ;
    input \addr_24__N_228[8] ;
    input \addr_24__N_228[6] ;
    input \addr_24__N_228[5] ;
    input \addr_24__N_228[4] ;
    input \addr_24__N_228[3] ;
    input \addr_24__N_228[2] ;
    input \addr_24__N_228[10] ;
    input \addr_24__N_228[11] ;
    input \addr_24__N_228[12] ;
    input \addr_24__N_228[13] ;
    input \addr_24__N_228[1] ;
    output n32031;
    
    wire qspi_clk_N_56 /* synthesis is_inv_clock=1, is_clock=1, SET_AS_NETWORK=\i_qspi/qspi_clk_N_56 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(8[22:35])
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    wire [24:0]addr_24__N_89;
    wire [3:0]qspi_data_out_3__N_51;
    wire [3:0]data_buff_in;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(29[15:27])
    
    wire spi_clk_pos_derived_59_enable_4, reading_dummy, qspi_clk_N_56_enable_1, 
        reading_dummy_N_262, error, qspi_clk_N_56_enable_2;
    wire [5:0]start_count;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(24[15:26])
    wire [5:0]n29;
    
    wire reading, writing, error_N_160, reading_N_139, n32082, n17761, 
        writing_N_151, n32081, n6579, n6587, n6595, n29094, n6583, 
        n6591, n29093;
    wire [12:0]n6481;
    wire [31:0]cmd;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(22[16:19])
    
    wire cmd_31__N_132, qspi_clk_N_56_enable_3, n29202, n29203, qspi_clk_N_56_enable_4;
    wire [3:0]qspi_data_out_3__N_257;
    wire [7:0]rom_buff_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(30[16:28])
    wire [3:0]qspi_data_out_3__N_253;
    
    wire n29174, n29175, n29177, n29178, n29180, n29181, n29183, 
        n29184, n6541, n6549, n6574, n30997, n6561, n6569, n30996, 
        n6538, n6546, n31008, n6558, n6566, n31007, n6580, n6588, 
        n29139, n6540, n6548, n31028, n6584, n6592, n29138, n6560, 
        n6568, n31027, n6581, n6589, n29133, n6585, n6593, n29132, 
        n6582, n6590, n29130, n6586, n6594, n29129;
    wire [7:0]ram_b_buff_out;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(32[16:30])
    
    wire n29208, n6559, n6567, n31078, n6539, n6547, n31079, qspi_clk_N_56_enable_5, 
        n11519;
    wire [11:0]n6497;
    
    wire ram_a_buff_out_7__N_127, n26312, n28596, n28592, n23673, 
        n23672, ram_b_buff_out_7__N_131, n26168, n26167, ram_b_buff_out_7__N_128, 
        addr_24__N_208, addr_24__N_212, addr_24__N_210, addr_24__N_214, 
        addr_24__N_216, addr_24__N_218, addr_24__N_220, n10521, addr_24__N_222, 
        addr_24__N_206, addr_24__N_204, addr_24__N_202, addr_24__N_200, 
        addr_24__N_224, n23671, n6532, n28702, n28704, n28660, n26016, 
        n28564, n28566, n26156, rom_buff_out_7__N_118;
    
    FD1S3AX addr_i2 (.D(addr_24__N_89[2]), .CK(qspi_clk_N_56), .Q(\addr[2] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i2.GSR = "ENABLED";
    FD1S3AX qspi_data_out_i0 (.D(qspi_data_out_3__N_51[0]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i0.GSR = "DISABLED";
    FD1P3AX data_buff_in_i0_i0 (.D(qspi_data_in_3__N_1[0]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i0.GSR = "DISABLED";
    FD1S3AX addr_i1 (.D(addr_24__N_89[1]), .CK(qspi_clk_N_56), .Q(\addr[1] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i1.GSR = "ENABLED";
    FD1P3AX data_buff_in_i0_i3 (.D(qspi_data_in_3__N_1[3]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i3.GSR = "DISABLED";
    FD1P3AX data_buff_in_i0_i2 (.D(qspi_data_in_3__N_1[2]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i2.GSR = "DISABLED";
    FD1P3AX data_buff_in_i0_i1 (.D(qspi_data_in_3__N_1[1]), .SP(spi_clk_pos_derived_59_enable_4), 
            .CK(spi_clk_pos_derived_59), .Q(data_buff_in[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam data_buff_in_i0_i1.GSR = "DISABLED";
    FD1P3AX reading_dummy_116 (.D(reading_dummy_N_262), .SP(qspi_clk_N_56_enable_1), 
            .CK(qspi_clk_N_56), .Q(reading_dummy)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam reading_dummy_116.GSR = "ENABLED";
    FD1P3AX error_118 (.D(VCC_net), .SP(qspi_clk_N_56_enable_2), .CK(qspi_clk_N_56), 
            .Q(error)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam error_118.GSR = "ENABLED";
    FD1S3AX start_count_3562__i0 (.D(n29[0]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562__i0.GSR = "ENABLED";
    LUT4 i27759_4_lut_then_3_lut_4_lut (.A(reading), .B(writing), .C(error_N_160), 
         .D(reading_N_139), .Z(n32082)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i27759_4_lut_then_3_lut_4_lut.init = 16'h1110;
    LUT4 i27759_4_lut_else_3_lut_4_lut (.A(reading), .B(writing), .C(n17761), 
         .D(writing_N_151), .Z(n32081)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i27759_4_lut_else_3_lut_4_lut.init = 16'h0100;
    LUT4 i26477_3_lut (.A(n6579), .B(n6587), .C(n6595), .Z(n29094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26477_3_lut.init = 16'hcaca;
    LUT4 i26476_3_lut (.A(n6583), .B(n6591), .C(n6595), .Z(n29093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26476_3_lut.init = 16'hcaca;
    FD1S3AX addr_res1_i0_i0 (.D(addr_24__N_89[1]), .CK(qspi_clk_N_56), .Q(n6481[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i0.GSR = "ENABLED";
    FD1S3AX qspi_data_out_i3 (.D(qspi_data_out_3__N_51[3]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i3.GSR = "DISABLED";
    FD1S3AX qspi_data_out_i2 (.D(qspi_data_out_3__N_51[2]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i2.GSR = "DISABLED";
    FD1S3AX qspi_data_out_i1 (.D(qspi_data_out_3__N_51[1]), .CK(qspi_clk_N_56), 
            .Q(qspi_data_in[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(110[12] 114[8])
    defparam qspi_data_out_i1.GSR = "DISABLED";
    FD1P3AX cmd_i0_i0 (.D(qspi_data_in_3__N_1[0]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i0.GSR = "ENABLED";
    FD1P3AX writing_117 (.D(n29202), .SP(qspi_clk_N_56_enable_3), .CK(qspi_clk_N_56), 
            .Q(writing)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam writing_117.GSR = "ENABLED";
    FD1P3AX reading_115 (.D(n29203), .SP(reading_N_139), .CK(qspi_clk_N_56), 
            .Q(reading)) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam reading_115.GSR = "ENABLED";
    FD1P3AX addr_i14 (.D(\addr_24__N_228[14] ), .SP(qspi_clk_N_56_enable_4), 
            .CK(qspi_clk_N_56), .Q(\addr[14] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i14.GSR = "ENABLED";
    FD1S3AX addr_i13 (.D(addr_24__N_89[13]), .CK(qspi_clk_N_56), .Q(\addr[13] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i13.GSR = "ENABLED";
    FD1S3AX addr_i12 (.D(addr_24__N_89[12]), .CK(qspi_clk_N_56), .Q(\addr[12] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i12.GSR = "ENABLED";
    FD1S3AX addr_i11 (.D(addr_24__N_89[11]), .CK(qspi_clk_N_56), .Q(\addr[11] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i11.GSR = "ENABLED";
    FD1S3AX addr_i10 (.D(addr_24__N_89[10]), .CK(qspi_clk_N_56), .Q(\addr[10] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i10.GSR = "ENABLED";
    FD1S3AX addr_i9 (.D(addr_24__N_89[9]), .CK(qspi_clk_N_56), .Q(\addr[9] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i9.GSR = "ENABLED";
    FD1S3AX addr_i8 (.D(addr_24__N_89[8]), .CK(qspi_clk_N_56), .Q(\addr[8] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i8.GSR = "ENABLED";
    FD1S3AX addr_i7 (.D(addr_24__N_89[7]), .CK(qspi_clk_N_56), .Q(\addr[7] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i7.GSR = "ENABLED";
    FD1S3AX addr_i6 (.D(addr_24__N_89[6]), .CK(qspi_clk_N_56), .Q(\addr[6] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i6.GSR = "ENABLED";
    FD1S3AX addr_i5 (.D(addr_24__N_89[5]), .CK(qspi_clk_N_56), .Q(\addr[5] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i5.GSR = "ENABLED";
    FD1S3AX addr_i4 (.D(addr_24__N_89[4]), .CK(qspi_clk_N_56), .Q(\addr[4] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i4.GSR = "ENABLED";
    FD1S3AX addr_i3 (.D(addr_24__N_89[3]), .CK(qspi_clk_N_56), .Q(\addr[3] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i3.GSR = "ENABLED";
    LUT4 i26562_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[0]), 
         .C(rom_buff_out[4]), .Z(qspi_data_out_3__N_253[0])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i26562_3_lut_3_lut.init = 16'he4e4;
    LUT4 i26559_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[3]), 
         .C(rom_buff_out[7]), .Z(qspi_data_out_3__N_253[3])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i26559_3_lut_3_lut.init = 16'he4e4;
    LUT4 i26565_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[2]), 
         .C(rom_buff_out[6]), .Z(qspi_data_out_3__N_253[2])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i26565_3_lut_3_lut.init = 16'he4e4;
    LUT4 i26568_3_lut_3_lut (.A(qspi_ram_a_select), .B(qspi_data_out_3__N_257[1]), 
         .C(rom_buff_out[5]), .Z(qspi_data_out_3__N_253[1])) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26:44])
    defparam i26568_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27275_3_lut_3_lut (.A(qspi_ram_b_select), .B(n29174), .C(rom_buff_out[3]), 
         .Z(n29175)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i27275_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27252_3_lut_3_lut (.A(qspi_ram_b_select), .B(n29177), .C(rom_buff_out[0]), 
         .Z(n29178)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i27252_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27277_3_lut_3_lut (.A(qspi_ram_b_select), .B(n29180), .C(rom_buff_out[2]), 
         .Z(n29181)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i27277_3_lut_3_lut.init = 16'he4e4;
    LUT4 i27279_3_lut_3_lut (.A(qspi_ram_b_select), .B(n29183), .C(rom_buff_out[1]), 
         .Z(n29184)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(112[26:44])
    defparam i27279_3_lut_3_lut.init = 16'he4e4;
    LUT4 n6561_bdd_3_lut (.A(n6541), .B(n6549), .C(n6574), .Z(n30997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n6561_bdd_3_lut.init = 16'hcaca;
    LUT4 n6561_bdd_3_lut_28191 (.A(n6561), .B(n6574), .C(n6569), .Z(n30996)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6561_bdd_3_lut_28191.init = 16'he2e2;
    LUT4 n6558_bdd_3_lut (.A(n6538), .B(n6546), .C(n6574), .Z(n31008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n6558_bdd_3_lut.init = 16'hcaca;
    LUT4 n6558_bdd_3_lut_28197 (.A(n6558), .B(n6574), .C(n6566), .Z(n31007)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6558_bdd_3_lut_28197.init = 16'he2e2;
    LUT4 i26522_3_lut (.A(n6580), .B(n6588), .C(n6595), .Z(n29139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26522_3_lut.init = 16'hcaca;
    FD1S3AX start_count_3562__i1 (.D(n29[1]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562__i1.GSR = "ENABLED";
    LUT4 n6560_bdd_3_lut (.A(n6540), .B(n6548), .C(n6574), .Z(n31028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n6560_bdd_3_lut.init = 16'hcaca;
    LUT4 i26521_3_lut (.A(n6584), .B(n6592), .C(n6595), .Z(n29138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26521_3_lut.init = 16'hcaca;
    LUT4 n6560_bdd_3_lut_28209 (.A(n6560), .B(n6574), .C(n6568), .Z(n31027)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6560_bdd_3_lut_28209.init = 16'he2e2;
    LUT4 i26516_3_lut (.A(n6581), .B(n6589), .C(n6595), .Z(n29133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26516_3_lut.init = 16'hcaca;
    LUT4 i26515_3_lut (.A(n6585), .B(n6593), .C(n6595), .Z(n29132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26515_3_lut.init = 16'hcaca;
    LUT4 i26513_3_lut (.A(n6582), .B(n6590), .C(n6595), .Z(n29130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26513_3_lut.init = 16'hcaca;
    LUT4 i26512_3_lut (.A(n6586), .B(n6594), .C(n6595), .Z(n29129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26512_3_lut.init = 16'hcaca;
    LUT4 i26560_3_lut (.A(ram_b_buff_out[4]), .B(ram_b_buff_out[0]), .C(\addr[0] ), 
         .Z(n29177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26560_3_lut.init = 16'hcaca;
    FD1S3AX start_count_3562__i2 (.D(n29[2]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562__i2.GSR = "ENABLED";
    FD1S3AX start_count_3562__i3 (.D(n29[3]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562__i3.GSR = "ENABLED";
    FD1S3AX start_count_3562__i4 (.D(n29[4]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562__i4.GSR = "ENABLED";
    FD1S3AX start_count_3562__i5 (.D(n29[5]), .CK(spi_clk_pos_derived_59), 
            .Q(start_count[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562__i5.GSR = "ENABLED";
    LUT4 i27861_3_lut (.A(reading), .B(writing), .C(error), .Z(cmd_31__N_132)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i27861_3_lut.init = 16'h0101;
    LUT4 i26566_3_lut (.A(ram_b_buff_out[5]), .B(ram_b_buff_out[1]), .C(\addr[0] ), 
         .Z(n29183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26566_3_lut.init = 16'hcaca;
    LUT4 i26563_3_lut (.A(ram_b_buff_out[6]), .B(ram_b_buff_out[2]), .C(\addr[0] ), 
         .Z(n29180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26563_3_lut.init = 16'hcaca;
    LUT4 i26557_3_lut (.A(ram_b_buff_out[7]), .B(ram_b_buff_out[3]), .C(\addr[0] ), 
         .Z(n29174)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26557_3_lut.init = 16'hcaca;
    PFUMX qspi_data_out_3__I_0_i1 (.BLUT(n29178), .ALUT(qspi_data_out_3__N_253[0]), 
          .C0(n29208), .Z(qspi_data_out_3__N_51[0])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    LUT4 n6559_bdd_3_lut_28240 (.A(n6559), .B(n6574), .C(n6567), .Z(n31078)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n6559_bdd_3_lut_28240.init = 16'he2e2;
    LUT4 n6559_bdd_3_lut (.A(n6539), .B(n6547), .C(n6574), .Z(n31079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n6559_bdd_3_lut.init = 16'hcaca;
    FD1P3IX addr_i0 (.D(\addr_24__N_228[0] ), .SP(qspi_clk_N_56_enable_5), 
            .CD(n11519), .CK(qspi_clk_N_56), .Q(\addr[0] )) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_i0.GSR = "ENABLED";
    FD1S3AX addr_res2_i0_i11 (.D(addr_24__N_89[12]), .CK(qspi_clk_N_56), 
            .Q(n6497[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res2_i0_i11.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i1 (.D(addr_24__N_89[2]), .CK(qspi_clk_N_56), .Q(n6481[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i1.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i2 (.D(addr_24__N_89[3]), .CK(qspi_clk_N_56), .Q(n6481[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i2.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i3 (.D(addr_24__N_89[4]), .CK(qspi_clk_N_56), .Q(n6481[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i3.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i4 (.D(addr_24__N_89[5]), .CK(qspi_clk_N_56), .Q(n6481[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i4.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i5 (.D(addr_24__N_89[6]), .CK(qspi_clk_N_56), .Q(n6481[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i5.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i6 (.D(addr_24__N_89[7]), .CK(qspi_clk_N_56), .Q(n6481[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i6.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i7 (.D(addr_24__N_89[8]), .CK(qspi_clk_N_56), .Q(n6481[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i7.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i8 (.D(addr_24__N_89[9]), .CK(qspi_clk_N_56), .Q(n6481[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i8.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i9 (.D(addr_24__N_89[10]), .CK(qspi_clk_N_56), 
            .Q(n6481[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i9.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i10 (.D(addr_24__N_89[11]), .CK(qspi_clk_N_56), 
            .Q(n6481[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i10.GSR = "ENABLED";
    FD1S3AX addr_res1_i0_i12 (.D(addr_24__N_89[13]), .CK(qspi_clk_N_56), 
            .Q(n6481[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam addr_res1_i0_i12.GSR = "ENABLED";
    LUT4 i27643_2_lut (.A(\addr[0] ), .B(qspi_ram_a_select), .Z(ram_a_buff_out_7__N_127)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i27643_2_lut.init = 16'h1111;
    LUT4 i1_4_lut (.A(start_count[3]), .B(n26312), .C(n28596), .D(\writing_N_164[3] ), 
         .Z(writing_N_151)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h2010;
    LUT4 i1_4_lut_adj_259 (.A(start_count[0]), .B(n28592), .C(start_count[1]), 
         .D(\writing_N_164[3] ), .Z(n28596)) /* synthesis lut_function=(!(A+((C (D)+!C !(D))+!B))) */ ;
    defparam i1_4_lut_adj_259.init = 16'h0440;
    LUT4 i1_3_lut (.A(start_count[2]), .B(error), .C(\writing_N_164[3] ), 
         .Z(n28592)) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(C)))) */ ;
    defparam i1_3_lut.init = 16'h1212;
    CCU2C start_count_3562_add_4_7 (.A0(start_count[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n23673), .S0(n29[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562_add_4_7.INIT0 = 16'haaa0;
    defparam start_count_3562_add_4_7.INIT1 = 16'h0000;
    defparam start_count_3562_add_4_7.INJECT1_0 = "NO";
    defparam start_count_3562_add_4_7.INJECT1_1 = "NO";
    CCU2C start_count_3562_add_4_5 (.A0(start_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(start_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23672), .COUT(n23673), .S0(n29[3]), .S1(n29[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562_add_4_5.INIT0 = 16'haaa0;
    defparam start_count_3562_add_4_5.INIT1 = 16'haaa0;
    defparam start_count_3562_add_4_5.INJECT1_0 = "NO";
    defparam start_count_3562_add_4_5.INJECT1_1 = "NO";
    FD1P3AX cmd_i0_i1 (.D(qspi_data_in_3__N_1[1]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i1.GSR = "ENABLED";
    LUT4 i23814_2_lut (.A(start_count[4]), .B(start_count[5]), .Z(n26312)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23814_2_lut.init = 16'heeee;
    FD1P3AX cmd_i0_i2 (.D(qspi_data_in_3__N_1[2]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i2.GSR = "ENABLED";
    FD1P3AX cmd_i0_i3 (.D(qspi_data_in_3__N_1[3]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i3.GSR = "ENABLED";
    FD1P3AX cmd_i0_i4 (.D(cmd[0]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[4])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i4.GSR = "ENABLED";
    FD1P3AX cmd_i0_i5 (.D(cmd[1]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[5])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i5.GSR = "ENABLED";
    FD1P3AX cmd_i0_i6 (.D(cmd[2]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[6])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i6.GSR = "ENABLED";
    FD1P3AX cmd_i0_i7 (.D(cmd[3]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[7])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i7.GSR = "ENABLED";
    FD1P3AX cmd_i0_i8 (.D(cmd[4]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[8])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i8.GSR = "ENABLED";
    FD1P3AX cmd_i0_i9 (.D(cmd[5]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[9])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i9.GSR = "ENABLED";
    FD1P3AX cmd_i0_i10 (.D(cmd[6]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[10])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i10.GSR = "ENABLED";
    FD1P3AX cmd_i0_i11 (.D(cmd[7]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[11])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i11.GSR = "ENABLED";
    FD1P3AX cmd_i0_i12 (.D(cmd[8]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[12])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i12.GSR = "ENABLED";
    FD1P3AX cmd_i0_i13 (.D(cmd[9]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[13])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i13.GSR = "ENABLED";
    FD1P3AX cmd_i0_i14 (.D(cmd[10]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[14])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i14.GSR = "ENABLED";
    FD1P3AX cmd_i0_i15 (.D(cmd[11]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[15])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i15.GSR = "ENABLED";
    FD1P3AX cmd_i0_i16 (.D(cmd[12]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[16])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i16.GSR = "ENABLED";
    FD1P3AX cmd_i0_i17 (.D(cmd[13]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[17])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i17.GSR = "ENABLED";
    FD1P3AX cmd_i0_i18 (.D(cmd[14]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[18])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i18.GSR = "ENABLED";
    FD1P3AX cmd_i0_i19 (.D(cmd[15]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[19])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i19.GSR = "ENABLED";
    FD1P3AX cmd_i0_i20 (.D(cmd[16]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[20])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i20.GSR = "ENABLED";
    FD1P3AX cmd_i0_i21 (.D(cmd[17]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[21])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i21.GSR = "ENABLED";
    FD1P3AX cmd_i0_i22 (.D(cmd[18]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[22])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i22.GSR = "ENABLED";
    FD1P3AX cmd_i0_i23 (.D(cmd[19]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[23])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i23.GSR = "ENABLED";
    FD1P3AX cmd_i0_i24 (.D(cmd[20]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[24])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i24.GSR = "ENABLED";
    FD1P3AX cmd_i0_i25 (.D(cmd[21]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[25])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i25.GSR = "ENABLED";
    FD1P3AX cmd_i0_i26 (.D(cmd[22]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[26])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i26.GSR = "ENABLED";
    FD1P3AX cmd_i0_i27 (.D(cmd[23]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[27])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i27.GSR = "ENABLED";
    FD1P3AX cmd_i0_i28 (.D(cmd[24]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[28])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i28.GSR = "ENABLED";
    FD1P3AX cmd_i0_i29 (.D(cmd[25]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[29])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i29.GSR = "ENABLED";
    FD1P3AX cmd_i0_i30 (.D(cmd[26]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[30])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i30.GSR = "ENABLED";
    FD1P3AX cmd_i0_i31 (.D(cmd[27]), .SP(cmd_31__N_132), .CK(spi_clk_pos_derived_59), 
            .Q(cmd[31])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(67[18] 75[12])
    defparam cmd_i0_i31.GSR = "ENABLED";
    LUT4 i27646_2_lut (.A(\addr[0] ), .B(qspi_ram_b_select), .Z(ram_b_buff_out_7__N_131)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i27646_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_4_lut (.A(writing), .B(\addr[0] ), .C(\addr[12] ), 
         .D(qspi_ram_a_select), .Z(n26168)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(49[14:31])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_260 (.A(writing), .B(\addr[0] ), .C(\addr[12] ), 
         .D(qspi_ram_a_select), .Z(n26167)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(49[14:31])
    defparam i1_2_lut_3_lut_4_lut_adj_260.init = 16'h0008;
    LUT4 ram_a_buff_out_7__N_124_I_0_2_lut_3_lut (.A(writing), .B(\addr[0] ), 
         .C(qspi_ram_b_select), .Z(ram_b_buff_out_7__N_128)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(49[14:31])
    defparam ram_a_buff_out_7__N_124_I_0_2_lut_3_lut.init = 16'h0808;
    LUT4 addr_24__I_0_i10_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[9] ), 
         .D(addr_24__N_208), .Z(addr_24__N_89[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i8_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[7] ), 
         .D(addr_24__N_212), .Z(addr_24__N_89[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i9_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[8] ), 
         .D(addr_24__N_210), .Z(addr_24__N_89[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i7_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[6] ), 
         .D(addr_24__N_214), .Z(addr_24__N_89[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i6_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[5] ), 
         .D(addr_24__N_216), .Z(addr_24__N_89[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i5_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[4] ), 
         .D(addr_24__N_218), .Z(addr_24__N_89[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i4_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[3] ), 
         .D(addr_24__N_220), .Z(addr_24__N_89[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i8893_2_lut_3_lut_4_lut (.A(reading), .B(writing), .C(reading_dummy), 
         .D(writing_N_151), .Z(n11519)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i8893_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i26585_4_lut_4_lut_4_lut (.A(reading), .B(writing), .C(n10521), 
         .D(reading_dummy), .Z(n29202)) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i26585_4_lut_4_lut_4_lut.init = 16'hcccd;
    LUT4 addr_24__I_0_i3_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[2] ), 
         .D(addr_24__N_222), .Z(addr_24__N_89[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i11_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[10] ), 
         .D(addr_24__N_206), .Z(addr_24__N_89[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i12_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[11] ), 
         .D(addr_24__N_204), .Z(addr_24__N_89[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i13_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[12] ), 
         .D(addr_24__N_202), .Z(addr_24__N_89[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 addr_24__I_0_i14_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[13] ), 
         .D(addr_24__N_200), .Z(addr_24__N_89[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_261 (.A(reading), .B(writing), .C(reading_dummy), 
         .D(writing_N_151), .Z(qspi_clk_N_56_enable_5)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i1_2_lut_3_lut_4_lut_adj_261.init = 16'hefee;
    LUT4 i26586_4_lut_3_lut (.A(reading), .B(writing), .C(reading_dummy), 
         .Z(n29203)) /* synthesis lut_function=(A+!(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam i26586_4_lut_3_lut.init = 16'hbaba;
    LUT4 addr_24__I_0_i2_3_lut_4_lut (.A(reading), .B(writing), .C(\addr_24__N_228[1] ), 
         .D(addr_24__N_224), .Z(addr_24__N_89[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam addr_24__I_0_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i27744_3_lut_rep_826 (.A(\writing_N_164[3] ), .B(qspi_ram_b_select), 
         .C(qspi_ram_a_select), .Z(n32031)) /* synthesis lut_function=(!(A (B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(34[23:82])
    defparam i27744_3_lut_rep_826.init = 16'h7f7f;
    LUT4 i27740_2_lut_4_lut (.A(\writing_N_164[3] ), .B(qspi_ram_b_select), 
         .C(qspi_ram_a_select), .D(\addr[0] ), .Z(spi_clk_pos_derived_59_enable_4)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(34[23:82])
    defparam i27740_2_lut_4_lut.init = 16'h007f;
    CCU2C start_count_3562_add_4_3 (.A0(start_count[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(start_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n23671), .COUT(n23672), .S0(n29[1]), .S1(n29[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562_add_4_3.INIT0 = 16'haaa0;
    defparam start_count_3562_add_4_3.INIT1 = 16'haaa0;
    defparam start_count_3562_add_4_3.INJECT1_0 = "NO";
    defparam start_count_3562_add_4_3.INJECT1_1 = "NO";
    CCU2C start_count_3562_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(start_count[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n23671), .S1(n29[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(61[35:50])
    defparam start_count_3562_add_4_1.INIT0 = 16'h0000;
    defparam start_count_3562_add_4_1.INIT1 = 16'h555f;
    defparam start_count_3562_add_4_1.INJECT1_0 = "NO";
    defparam start_count_3562_add_4_1.INJECT1_1 = "NO";
    PFUMX qspi_data_out_3__I_0_i2 (.BLUT(n29184), .ALUT(qspi_data_out_3__N_253[1]), 
          .C0(n29208), .Z(qspi_data_out_3__N_51[1])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    PFUMX i28241 (.BLUT(n31079), .ALUT(n31078), .C0(n6532), .Z(rom_buff_out[1]));
    PFUMX qspi_data_out_3__I_0_i3 (.BLUT(n29181), .ALUT(qspi_data_out_3__N_253[2]), 
          .C0(n29208), .Z(qspi_data_out_3__N_51[2])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    PFUMX i26514 (.BLUT(n29129), .ALUT(n29130), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[3]));
    LUT4 i27775_3_lut (.A(qspi_ram_a_select), .B(qspi_ram_b_select), .C(\addr[0] ), 
         .Z(n29208)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(111[26] 113[96])
    defparam i27775_3_lut.init = 16'h5d5d;
    PFUMX i28210 (.BLUT(n31028), .ALUT(n31027), .C0(n6532), .Z(rom_buff_out[2]));
    LUT4 i27705_4_lut (.A(n28702), .B(n28704), .C(start_count[2]), .D(start_count[1]), 
         .Z(reading_N_139)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(93[21:38])
    defparam i27705_4_lut.init = 16'h0010;
    LUT4 i1_2_lut (.A(start_count[3]), .B(start_count[4]), .Z(n28702)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(93[21:38])
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_adj_262 (.A(start_count[0]), .B(start_count[5]), .Z(n28704)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(93[21:38])
    defparam i1_2_lut_adj_262.init = 16'heeee;
    LUT4 i1_4_lut_adj_263 (.A(n28660), .B(n26312), .C(start_count[3]), 
         .D(cmd[3]), .Z(error_N_160)) /* synthesis lut_function=(!(A (B+(C))+!A (B+(C+(D))))) */ ;
    defparam i1_4_lut_adj_263.init = 16'h0203;
    LUT4 i1_3_lut_adj_264 (.A(cmd[1]), .B(cmd[2]), .C(cmd[0]), .Z(n28660)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_3_lut_adj_264.init = 16'hfdfd;
    LUT4 i15196_4_lut (.A(\writing_N_164[3] ), .B(cmd[27]), .C(n26016), 
         .D(cmd[24]), .Z(n17761)) /* synthesis lut_function=(A ((C+!(D))+!B)) */ ;
    defparam i15196_4_lut.init = 16'ha2aa;
    LUT4 i1_4_lut_adj_265 (.A(n28564), .B(cmd[25]), .C(n28566), .D(cmd[26]), 
         .Z(n26016)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(102[26:45])
    defparam i1_4_lut_adj_265.init = 16'hfffb;
    LUT4 i1_2_lut_adj_266 (.A(cmd[29]), .B(cmd[30]), .Z(n28564)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(102[26:45])
    defparam i1_2_lut_adj_266.init = 16'heeee;
    LUT4 i1_2_lut_adj_267 (.A(cmd[31]), .B(cmd[28]), .Z(n28566)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(102[26:45])
    defparam i1_2_lut_adj_267.init = 16'heeee;
    PFUMX i26517 (.BLUT(n29132), .ALUT(n29133), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[2]));
    PFUMX i26523 (.BLUT(n29138), .ALUT(n29139), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[1]));
    PFUMX i28198 (.BLUT(n31008), .ALUT(n31007), .C0(n6532), .Z(rom_buff_out[0]));
    PFUMX qspi_data_out_3__I_0_i4 (.BLUT(n29175), .ALUT(qspi_data_out_3__N_253[3]), 
          .C0(n29208), .Z(qspi_data_out_3__N_51[3])) /* synthesis LSE_LINE_FILE_ID=17, LSE_LCOL=19, LSE_RCOL=6, LSE_LLINE=42, LSE_RLINE=50 */ ;
    PFUMX i28192 (.BLUT(n30997), .ALUT(n30996), .C0(n6532), .Z(rom_buff_out[3]));
    LUT4 reading_I_0_126_2_lut_rep_856 (.A(reading), .B(writing), .Z(qspi_clk_N_56_enable_4)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(86[17:35])
    defparam reading_I_0_126_2_lut_rep_856.init = 16'heeee;
    LUT4 i27734_4_lut (.A(n26156), .B(qspi_clk_N_56_enable_4), .C(error_N_160), 
         .D(reading_dummy), .Z(qspi_clk_N_56_enable_2)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(85[18] 107[12])
    defparam i27734_4_lut.init = 16'h3022;
    LUT4 i1_3_lut_adj_268 (.A(cmd[27]), .B(n26016), .C(cmd[24]), .Z(n10521)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(102[26:45])
    defparam i1_3_lut_adj_268.init = 16'hfefe;
    LUT4 i1_2_lut_rep_692 (.A(writing_N_151), .B(n17761), .Z(qspi_clk_N_56_enable_3)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_692.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(writing_N_151), .B(n17761), .C(n10521), .Z(n26156)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i8807_2_lut_3_lut (.A(n17761), .B(writing_N_151), .C(reading_dummy), 
         .Z(reading_dummy_N_262)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i8807_2_lut_3_lut.init = 16'h0404;
    LUT4 i27640_2_lut (.A(\addr[0] ), .B(\writing_N_164[3] ), .Z(rom_buff_out_7__N_118)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i27640_2_lut.init = 16'h1111;
    LUT4 i5288_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[0]), 
         .D(\addr[1] ), .Z(addr_24__N_224)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5288_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5286_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[1]), 
         .D(\addr[2] ), .Z(addr_24__N_222)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5286_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5264_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[12]), 
         .D(\addr[13] ), .Z(addr_24__N_200)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5264_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5266_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[11]), 
         .D(\addr[12] ), .Z(addr_24__N_202)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5266_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5268_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[10]), 
         .D(\addr[11] ), .Z(addr_24__N_204)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5268_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5270_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[9]), 
         .D(\addr[10] ), .Z(addr_24__N_206)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5270_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5272_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[8]), 
         .D(\addr[9] ), .Z(addr_24__N_208)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5272_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5274_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[7]), 
         .D(\addr[8] ), .Z(addr_24__N_210)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5274_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5276_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[6]), 
         .D(\addr[7] ), .Z(addr_24__N_212)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5276_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5278_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[5]), 
         .D(\addr[6] ), .Z(addr_24__N_214)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5278_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5280_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[4]), 
         .D(\addr[5] ), .Z(addr_24__N_216)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5280_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5282_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[3]), 
         .D(\addr[4] ), .Z(addr_24__N_218)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5282_3_lut_4_lut.init = 16'hfd20;
    LUT4 i5284_3_lut_4_lut (.A(writing_N_151), .B(reading_dummy), .C(cmd[2]), 
         .D(\addr[3] ), .Z(addr_24__N_220)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(97[22] 106[16])
    defparam i5284_3_lut_4_lut.init = 16'hfd20;
    PFUMX i26478 (.BLUT(n29093), .ALUT(n29094), .C0(\addr[0] ), .Z(qspi_data_out_3__N_257[0]));
    PFUMX i28624 (.BLUT(n32081), .ALUT(n32082), .C0(reading_dummy), .Z(qspi_clk_N_56_enable_1));
    \BRAM(ADDR_WIDTH=13)  rom (.n6574(n6574), .\addr[1] (\addr[1] ), .\addr[2] (\addr[2] ), 
            .\addr[3] (\addr[3] ), .\addr[4] (\addr[4] ), .\addr[5] (\addr[5] ), 
            .\addr[6] (\addr[6] ), .\addr[7] (\addr[7] ), .\addr[8] (\addr[8] ), 
            .\addr[9] (\addr[9] ), .\addr[10] (\addr[10] ), .\addr[11] (\addr[11] ), 
            .n6485(n6481[0]), .n6480(n6481[1]), .n6479(n6481[2]), .n6478(n6481[3]), 
            .n6477(n6481[4]), .n6476(n6481[5]), .n6475(n6481[6]), .n6474(n6481[7]), 
            .n6473(n6481[8]), .n6472(n6481[9]), .n6471(n6481[10]), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .data_buff_in({data_buff_in}), .n6566(n6566), .n6567(n6567), 
            .n6568(n6568), .n6569(n6569), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .GND_net(GND_net), .rom_buff_out_7__N_118(rom_buff_out_7__N_118), 
            .VCC_net(VCC_net), .n6558(n6558), .n6559(n6559), .n6560(n6560), 
            .n6561(n6561), .n6486(n6497[11]), .n6538(n6538), .n6539(n6539), 
            .n6540(n6540), .n6541(n6541), .n6546(n6546), .n6547(n6547), 
            .n6548(n6548), .n6549(n6549), .n6532(n6532), .n6469(n6481[12]), 
            .\rom_buff_out[6] (rom_buff_out[6]), .\rom_buff_out[5] (rom_buff_out[5]), 
            .\rom_buff_out[4] (rom_buff_out[4]), .\rom_buff_out[7] (rom_buff_out[7])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(36[58] 43[6])
    \BRAM(ADDR_WIDTH=11)  ram_b (.\addr[1] (\addr[1] ), .\addr[2] (\addr[2] ), 
            .\addr[3] (\addr[3] ), .\addr[4] (\addr[4] ), .\addr[5] (\addr[5] ), 
            .\addr[6] (\addr[6] ), .\addr[7] (\addr[7] ), .\addr[8] (\addr[8] ), 
            .\addr[9] (\addr[9] ), .\addr[10] (\addr[10] ), .\addr[11] (\addr[11] ), 
            .n6485(n6481[0]), .n6480(n6481[1]), .n6479(n6481[2]), .n6478(n6481[3]), 
            .n6477(n6481[4]), .n6476(n6481[5]), .n6475(n6481[6]), .n6474(n6481[7]), 
            .n6473(n6481[8]), .n6472(n6481[9]), .n6471(n6481[10]), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .data_buff_in({data_buff_in}), .ram_b_buff_out({ram_b_buff_out}), 
            .spi_clk_pos_derived_59(spi_clk_pos_derived_59), .ram_b_buff_out_7__N_128(ram_b_buff_out_7__N_128), 
            .ram_b_buff_out_7__N_131(ram_b_buff_out_7__N_131), .GND_net(GND_net), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(52[37] 59[6])
    \BRAM(ADDR_WIDTH=12)  ram_a (.\addr[1] (\addr[1] ), .\addr[2] (\addr[2] ), 
            .\addr[3] (\addr[3] ), .\addr[4] (\addr[4] ), .\addr[5] (\addr[5] ), 
            .\addr[6] (\addr[6] ), .\addr[7] (\addr[7] ), .\addr[8] (\addr[8] ), 
            .\addr[9] (\addr[9] ), .\addr[10] (\addr[10] ), .\addr[11] (\addr[11] ), 
            .n6485(n6481[0]), .n6480(n6481[1]), .n6479(n6481[2]), .n6478(n6481[3]), 
            .n6477(n6481[4]), .n6476(n6481[5]), .n6475(n6481[6]), .n6474(n6481[7]), 
            .n6473(n6481[8]), .n6472(n6481[9]), .n6471(n6481[10]), .qspi_data_in_3__N_1({qspi_data_in_3__N_1}), 
            .data_buff_in({data_buff_in}), .n6587(n6587), .n6588(n6588), 
            .n6589(n6589), .n6590(n6590), .n6591(n6591), .n6592(n6592), 
            .n6593(n6593), .n6594(n6594), .spi_clk_pos_derived_59(spi_clk_pos_derived_59), 
            .n26168(n26168), .ram_a_buff_out_7__N_127(ram_a_buff_out_7__N_127), 
            .GND_net(GND_net), .VCC_net(VCC_net), .n6579(n6579), .n6580(n6580), 
            .n6581(n6581), .n6582(n6582), .n6583(n6583), .n6584(n6584), 
            .n6585(n6585), .n6586(n6586), .n26167(n26167), .n6595(n6595), 
            .n6486(n6497[11])) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/sim_qspi.v(44[37] 51[6])
    
endmodule
//
// Verilog Description of module \BRAM(ADDR_WIDTH=13) 
//

module \BRAM(ADDR_WIDTH=13)  (n6574, \addr[1] , \addr[2] , \addr[3] , 
            \addr[4] , \addr[5] , \addr[6] , \addr[7] , \addr[8] , 
            \addr[9] , \addr[10] , \addr[11] , n6485, n6480, n6479, 
            n6478, n6477, n6476, n6475, n6474, n6473, n6472, n6471, 
            qspi_data_in_3__N_1, data_buff_in, n6566, n6567, n6568, 
            n6569, spi_clk_pos_derived_59, GND_net, rom_buff_out_7__N_118, 
            VCC_net, n6558, n6559, n6560, n6561, n6486, n6538, 
            n6539, n6540, n6541, n6546, n6547, n6548, n6549, n6532, 
            n6469, \rom_buff_out[6] , \rom_buff_out[5] , \rom_buff_out[4] , 
            \rom_buff_out[7] ) /* synthesis syn_module_defined=1 */ ;
    output n6574;
    input \addr[1] ;
    input \addr[2] ;
    input \addr[3] ;
    input \addr[4] ;
    input \addr[5] ;
    input \addr[6] ;
    input \addr[7] ;
    input \addr[8] ;
    input \addr[9] ;
    input \addr[10] ;
    input \addr[11] ;
    input n6485;
    input n6480;
    input n6479;
    input n6478;
    input n6477;
    input n6476;
    input n6475;
    input n6474;
    input n6473;
    input n6472;
    input n6471;
    input [3:0]qspi_data_in_3__N_1;
    input [3:0]data_buff_in;
    output n6566;
    output n6567;
    output n6568;
    output n6569;
    input spi_clk_pos_derived_59;
    input GND_net;
    input rom_buff_out_7__N_118;
    input VCC_net;
    output n6558;
    output n6559;
    output n6560;
    output n6561;
    input n6486;
    output n6538;
    output n6539;
    output n6540;
    output n6541;
    output n6546;
    output n6547;
    output n6548;
    output n6549;
    output n6532;
    input n6469;
    output \rom_buff_out[6] ;
    output \rom_buff_out[5] ;
    output \rom_buff_out[4] ;
    output \rom_buff_out[7] ;
    
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    wire n6565, n6573, n29106, n6545, n6553, n29105, n6570, n6571, 
        n6572, n6562, n6563, n6564, n6542, n6543, n6544, n6550, 
        n6551, n6552, n29115, n29114, n29112, n29111, n29109, 
        n29108;
    
    LUT4 i26489_3_lut (.A(n6565), .B(n6573), .C(n6574), .Z(n29106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26489_3_lut.init = 16'hcaca;
    LUT4 i26488_3_lut (.A(n6545), .B(n6553), .C(n6574), .Z(n29105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26488_3_lut.init = 16'hcaca;
    DP16KD mem3 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6485), .ADB4(n6480), 
           .ADB5(n6479), .ADB6(n6478), .ADB7(n6477), .ADB8(n6476), .ADB9(n6475), 
           .ADB10(n6474), .ADB11(n6473), .ADB12(n6472), .ADB13(n6471), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6566), .DOB1(n6567), .DOB2(n6568), 
           .DOB3(n6569), .DOB4(n6570), .DOB5(n6571), .DOB6(n6572), .DOB7(n6573));
    defparam mem3.DATA_WIDTH_A = 9;
    defparam mem3.DATA_WIDTH_B = 9;
    defparam mem3.REGMODE_A = "NOREG";
    defparam mem3.REGMODE_B = "NOREG";
    defparam mem3.RESETMODE = "SYNC";
    defparam mem3.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem3.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem3.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem3.CSDECODE_A = "0b000";
    defparam mem3.CSDECODE_B = "0b000";
    defparam mem3.GSR = "DISABLED";
    defparam mem3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem3.INIT_DATA = "STATIC";
    DP16KD mem1 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6485), .ADB4(n6480), 
           .ADB5(n6479), .ADB6(n6478), .ADB7(n6477), .ADB8(n6476), .ADB9(n6475), 
           .ADB10(n6474), .ADB11(n6473), .ADB12(n6472), .ADB13(n6471), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6558), .DOB1(n6559), .DOB2(n6560), 
           .DOB3(n6561), .DOB4(n6562), .DOB5(n6563), .DOB6(n6564), .DOB7(n6565));
    defparam mem1.DATA_WIDTH_A = 9;
    defparam mem1.DATA_WIDTH_B = 9;
    defparam mem1.REGMODE_A = "NOREG";
    defparam mem1.REGMODE_B = "NOREG";
    defparam mem1.RESETMODE = "SYNC";
    defparam mem1.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem1.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem1.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem1.CSDECODE_A = "0b000";
    defparam mem1.CSDECODE_B = "0b000";
    defparam mem1.GSR = "DISABLED";
    defparam mem1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INIT_DATA = "STATIC";
    FD1P3AX i4305 (.D(n6486), .SP(rom_buff_out_7__N_118), .CK(spi_clk_pos_derived_59), 
            .Q(n6574));
    defparam i4305.GSR = "DISABLED";
    DP16KD mem0 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6485), .ADB4(n6480), 
           .ADB5(n6479), .ADB6(n6478), .ADB7(n6477), .ADB8(n6476), .ADB9(n6475), 
           .ADB10(n6474), .ADB11(n6473), .ADB12(n6472), .ADB13(n6471), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6538), .DOB1(n6539), .DOB2(n6540), 
           .DOB3(n6541), .DOB4(n6542), .DOB5(n6543), .DOB6(n6544), .DOB7(n6545));
    defparam mem0.DATA_WIDTH_A = 9;
    defparam mem0.DATA_WIDTH_B = 9;
    defparam mem0.REGMODE_A = "NOREG";
    defparam mem0.REGMODE_B = "NOREG";
    defparam mem0.RESETMODE = "SYNC";
    defparam mem0.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem0.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem0.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem0.CSDECODE_A = "0b000";
    defparam mem0.CSDECODE_B = "0b000";
    defparam mem0.GSR = "DISABLED";
    defparam mem0.INITVAL_00 = "0x00000000000000000004108E7080840088A002F50E8930682004A731E02400C800006F00A000006F";
    defparam mem0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_02 = "0x00280002170100000437080011029300200002B7000000024A000000008000000000700000000070";
    defparam mem0.INITVAL_03 = "0x0602000073068820684416073000A4128B30888506020000731400105079004C0000EF1F44100213";
    defparam mem0.INITVAL_04 = "0x1D80110E93000E61F2631D80110E131D80110C930602000073068820604416073000A4128B308885";
    defparam mem0.INITVAL_05 = "0x11C911FEF710C93004F60EA630008710E931800110C130020000EB71FCE71DAE300EC1000071C023";
    defparam mem0.INITVAL_06 = "0x1FCD7136E31FCC705C2300E1100E91086900382000E9312CB21800110E1300C910382000C13134F1";
    defparam mem0.INITVAL_07 = "0x00EC100E41000A71E023000070EA03040A000E131D80110E93000670FC631D801106131D80110E13";
    defparam mem0.INITVAL_08 = "0x08E92184021849008C05022F700E130400610C93022610000714E371000000CB7100821FC671D4E3";
    defparam mem0.INITVAL_09 = "0x00E8508E821FCF7082E308E821800200006140231FCF70B8E308E921843E00E8508E92000F709063";
    defparam mem0.INITVAL_0A = "0x0009500E63188811089300A051D026102040049500263180011688317EC91FCF70B8E308E821803E";
    defparam mem0.INITVAL_0B = "0x10E1306020000730688206045060730000800A3717ECD1808110A13060200007306882180A114423";
    defparam mem0.INITVAL_0C = "0x0000800AB7180B114023000B601C63000E511A6300A85112881800116A83060061607308CA118881";
    defparam mem0.INITVAL_0D = "0x06006160731FCE601CE31804114E03060061407316EDD1808110A931008206006140730604514073";
    defparam mem0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000020000008002000000817EE1";
    defparam mem0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INIT_DATA = "STATIC";
    DP16KD mem2 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(GND_net), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6485), .ADB4(n6480), 
           .ADB5(n6479), .ADB6(n6478), .ADB7(n6477), .ADB8(n6476), .ADB9(n6475), 
           .ADB10(n6474), .ADB11(n6473), .ADB12(n6472), .ADB13(n6471), 
           .CEB(rom_buff_out_7__N_118), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6546), .DOB1(n6547), .DOB2(n6548), 
           .DOB3(n6549), .DOB4(n6550), .DOB5(n6551), .DOB6(n6552), .DOB7(n6553));
    defparam mem2.DATA_WIDTH_A = 9;
    defparam mem2.DATA_WIDTH_B = 9;
    defparam mem2.REGMODE_A = "NOREG";
    defparam mem2.REGMODE_B = "NOREG";
    defparam mem2.RESETMODE = "SYNC";
    defparam mem2.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem2.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem2.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem2.CSDECODE_A = "0b000";
    defparam mem2.CSDECODE_B = "0b000";
    defparam mem2.GSR = "DISABLED";
    defparam mem2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem2.INIT_DATA = "STATIC";
    FD1P3AX i4287 (.D(n6469), .SP(rom_buff_out_7__N_118), .CK(spi_clk_pos_derived_59), 
            .Q(n6532));
    defparam i4287.GSR = "DISABLED";
    LUT4 i26498_3_lut (.A(n6562), .B(n6570), .C(n6574), .Z(n29115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26498_3_lut.init = 16'hcaca;
    LUT4 i26497_3_lut (.A(n6542), .B(n6550), .C(n6574), .Z(n29114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26497_3_lut.init = 16'hcaca;
    LUT4 i26495_3_lut (.A(n6563), .B(n6571), .C(n6574), .Z(n29112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26495_3_lut.init = 16'hcaca;
    LUT4 i26494_3_lut (.A(n6543), .B(n6551), .C(n6574), .Z(n29111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26494_3_lut.init = 16'hcaca;
    LUT4 i26492_3_lut (.A(n6564), .B(n6572), .C(n6574), .Z(n29109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26492_3_lut.init = 16'hcaca;
    LUT4 i26491_3_lut (.A(n6544), .B(n6552), .C(n6574), .Z(n29108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i26491_3_lut.init = 16'hcaca;
    PFUMX i26493 (.BLUT(n29108), .ALUT(n29109), .C0(n6532), .Z(\rom_buff_out[6] ));
    PFUMX i26496 (.BLUT(n29111), .ALUT(n29112), .C0(n6532), .Z(\rom_buff_out[5] ));
    PFUMX i26499 (.BLUT(n29114), .ALUT(n29115), .C0(n6532), .Z(\rom_buff_out[4] ));
    PFUMX i26490 (.BLUT(n29105), .ALUT(n29106), .C0(n6532), .Z(\rom_buff_out[7] ));
    
endmodule
//
// Verilog Description of module \BRAM(ADDR_WIDTH=11) 
//

module \BRAM(ADDR_WIDTH=11)  (\addr[1] , \addr[2] , \addr[3] , \addr[4] , 
            \addr[5] , \addr[6] , \addr[7] , \addr[8] , \addr[9] , 
            \addr[10] , \addr[11] , n6485, n6480, n6479, n6478, 
            n6477, n6476, n6475, n6474, n6473, n6472, n6471, qspi_data_in_3__N_1, 
            data_buff_in, ram_b_buff_out, spi_clk_pos_derived_59, ram_b_buff_out_7__N_128, 
            ram_b_buff_out_7__N_131, GND_net, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input \addr[1] ;
    input \addr[2] ;
    input \addr[3] ;
    input \addr[4] ;
    input \addr[5] ;
    input \addr[6] ;
    input \addr[7] ;
    input \addr[8] ;
    input \addr[9] ;
    input \addr[10] ;
    input \addr[11] ;
    input n6485;
    input n6480;
    input n6479;
    input n6478;
    input n6477;
    input n6476;
    input n6475;
    input n6474;
    input n6473;
    input n6472;
    input n6471;
    input [3:0]qspi_data_in_3__N_1;
    input [3:0]data_buff_in;
    output [7:0]ram_b_buff_out;
    input spi_clk_pos_derived_59;
    input ram_b_buff_out_7__N_128;
    input ram_b_buff_out_7__N_131;
    input GND_net;
    input VCC_net;
    
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    DP16KD mem0 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(ram_b_buff_out_7__N_128), .CSA0(GND_net), .CSA1(GND_net), 
           .CSA2(GND_net), .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), 
           .DIB2(GND_net), .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), 
           .DIB6(GND_net), .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), 
           .DIB10(GND_net), .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), 
           .DIB14(GND_net), .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), 
           .ADB0(GND_net), .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6485), 
           .ADB4(n6480), .ADB5(n6479), .ADB6(n6478), .ADB7(n6477), .ADB8(n6476), 
           .ADB9(n6475), .ADB10(n6474), .ADB11(n6473), .ADB12(n6472), 
           .ADB13(n6471), .CEB(ram_b_buff_out_7__N_131), .OCEB(VCC_net), 
           .CLKB(spi_clk_pos_derived_59), .WEB(GND_net), .CSB0(GND_net), 
           .CSB1(GND_net), .CSB2(GND_net), .RSTB(GND_net), .DOB0(ram_b_buff_out[0]), 
           .DOB1(ram_b_buff_out[1]), .DOB2(ram_b_buff_out[2]), .DOB3(ram_b_buff_out[3]), 
           .DOB4(ram_b_buff_out[4]), .DOB5(ram_b_buff_out[5]), .DOB6(ram_b_buff_out[6]), 
           .DOB7(ram_b_buff_out[7]));
    defparam mem0.DATA_WIDTH_A = 9;
    defparam mem0.DATA_WIDTH_B = 9;
    defparam mem0.REGMODE_A = "NOREG";
    defparam mem0.REGMODE_B = "NOREG";
    defparam mem0.RESETMODE = "SYNC";
    defparam mem0.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem0.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem0.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem0.CSDECODE_A = "0b000";
    defparam mem0.CSDECODE_B = "0b000";
    defparam mem0.GSR = "DISABLED";
    defparam mem0.INITVAL_00 = "0x00000000000000000004108E7080840088A002F50E8930682004A731E02400C800006F00A000006F";
    defparam mem0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_02 = "0x00280002170100000437080011029300200002B7000000024A000000008000000000700000000070";
    defparam mem0.INITVAL_03 = "0x0602000073068820684416073000A4128B30888506020000731400105079004C0000EF1F44100213";
    defparam mem0.INITVAL_04 = "0x1D80110E93000E61F2631D80110E131D80110C930602000073068820604416073000A4128B308885";
    defparam mem0.INITVAL_05 = "0x11C911FEF710C93004F60EA630008710E931800110C130020000EB71FCE71DAE300EC1000071C023";
    defparam mem0.INITVAL_06 = "0x1FCD7136E31FCC705C2300E1100E91086900382000E9312CB21800110E1300C910382000C13134F1";
    defparam mem0.INITVAL_07 = "0x00EC100E41000A71E023000070EA03040A000E131D80110E93000670FC631D801106131D80110E13";
    defparam mem0.INITVAL_08 = "0x08E92184021849008C05022F700E130400610C93022610000714E371000000CB7100821FC671D4E3";
    defparam mem0.INITVAL_09 = "0x00E8508E821FCF7082E308E821800200006140231FCF70B8E308E921843E00E8508E92000F709063";
    defparam mem0.INITVAL_0A = "0x0009500E63188811089300A051D026102040049500263180011688317EC91FCF70B8E308E821803E";
    defparam mem0.INITVAL_0B = "0x10E1306020000730688206045060730000800A3717ECD1808110A13060200007306882180A114423";
    defparam mem0.INITVAL_0C = "0x0000800AB7180B114023000B601C63000E511A6300A85112881800116A83060061607308CA118881";
    defparam mem0.INITVAL_0D = "0x06006160731FCE601CE31804114E03060061407316EDD1808110A931008206006140730604514073";
    defparam mem0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000020000008002000000817EE1";
    defparam mem0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INIT_DATA = "STATIC";
    
endmodule
//
// Verilog Description of module \BRAM(ADDR_WIDTH=12) 
//

module \BRAM(ADDR_WIDTH=12)  (\addr[1] , \addr[2] , \addr[3] , \addr[4] , 
            \addr[5] , \addr[6] , \addr[7] , \addr[8] , \addr[9] , 
            \addr[10] , \addr[11] , n6485, n6480, n6479, n6478, 
            n6477, n6476, n6475, n6474, n6473, n6472, n6471, qspi_data_in_3__N_1, 
            data_buff_in, n6587, n6588, n6589, n6590, n6591, n6592, 
            n6593, n6594, spi_clk_pos_derived_59, n26168, ram_a_buff_out_7__N_127, 
            GND_net, VCC_net, n6579, n6580, n6581, n6582, n6583, 
            n6584, n6585, n6586, n26167, n6595, n6486) /* synthesis syn_module_defined=1 */ ;
    input \addr[1] ;
    input \addr[2] ;
    input \addr[3] ;
    input \addr[4] ;
    input \addr[5] ;
    input \addr[6] ;
    input \addr[7] ;
    input \addr[8] ;
    input \addr[9] ;
    input \addr[10] ;
    input \addr[11] ;
    input n6485;
    input n6480;
    input n6479;
    input n6478;
    input n6477;
    input n6476;
    input n6475;
    input n6474;
    input n6473;
    input n6472;
    input n6471;
    input [3:0]qspi_data_in_3__N_1;
    input [3:0]data_buff_in;
    output n6587;
    output n6588;
    output n6589;
    output n6590;
    output n6591;
    output n6592;
    output n6593;
    output n6594;
    input spi_clk_pos_derived_59;
    input n26168;
    input ram_a_buff_out_7__N_127;
    input GND_net;
    input VCC_net;
    output n6579;
    output n6580;
    output n6581;
    output n6582;
    output n6583;
    output n6584;
    output n6585;
    output n6586;
    input n26167;
    output n6595;
    input n6486;
    
    wire spi_clk_pos_derived_59 /* synthesis is_clock=1, SET_AS_NETWORK=\i_tinyqv/mem/q_ctrl/spi_clk_pos_derived_59 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase3/projetotinyqv/projetotinyqv/impl1/source/qspi_ctrl.v(89[15:26])
    
    DP16KD mem1 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(n26168), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6485), .ADB4(n6480), 
           .ADB5(n6479), .ADB6(n6478), .ADB7(n6477), .ADB8(n6476), .ADB9(n6475), 
           .ADB10(n6474), .ADB11(n6473), .ADB12(n6472), .ADB13(n6471), 
           .CEB(ram_a_buff_out_7__N_127), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6587), .DOB1(n6588), .DOB2(n6589), 
           .DOB3(n6590), .DOB4(n6591), .DOB5(n6592), .DOB6(n6593), .DOB7(n6594));
    defparam mem1.DATA_WIDTH_A = 9;
    defparam mem1.DATA_WIDTH_B = 9;
    defparam mem1.REGMODE_A = "NOREG";
    defparam mem1.REGMODE_B = "NOREG";
    defparam mem1.RESETMODE = "SYNC";
    defparam mem1.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem1.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem1.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem1.CSDECODE_A = "0b000";
    defparam mem1.CSDECODE_B = "0b000";
    defparam mem1.GSR = "DISABLED";
    defparam mem1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem1.INIT_DATA = "STATIC";
    DP16KD mem0 (.DIA0(qspi_data_in_3__N_1[0]), .DIA1(qspi_data_in_3__N_1[1]), 
           .DIA2(qspi_data_in_3__N_1[2]), .DIA3(qspi_data_in_3__N_1[3]), 
           .DIA4(data_buff_in[0]), .DIA5(data_buff_in[1]), .DIA6(data_buff_in[2]), 
           .DIA7(data_buff_in[3]), .DIA8(GND_net), .DIA9(GND_net), .DIA10(GND_net), 
           .DIA11(GND_net), .DIA12(GND_net), .DIA13(GND_net), .DIA14(GND_net), 
           .DIA15(GND_net), .DIA16(GND_net), .DIA17(GND_net), .ADA0(GND_net), 
           .ADA1(GND_net), .ADA2(GND_net), .ADA3(\addr[1] ), .ADA4(\addr[2] ), 
           .ADA5(\addr[3] ), .ADA6(\addr[4] ), .ADA7(\addr[5] ), .ADA8(\addr[6] ), 
           .ADA9(\addr[7] ), .ADA10(\addr[8] ), .ADA11(\addr[9] ), .ADA12(\addr[10] ), 
           .ADA13(\addr[11] ), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(spi_clk_pos_derived_59), 
           .WEA(n26167), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
           .RSTA(GND_net), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
           .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
           .DIB7(GND_net), .DIB8(GND_net), .DIB9(GND_net), .DIB10(GND_net), 
           .DIB11(GND_net), .DIB12(GND_net), .DIB13(GND_net), .DIB14(GND_net), 
           .DIB15(GND_net), .DIB16(GND_net), .DIB17(GND_net), .ADB0(GND_net), 
           .ADB1(GND_net), .ADB2(GND_net), .ADB3(n6485), .ADB4(n6480), 
           .ADB5(n6479), .ADB6(n6478), .ADB7(n6477), .ADB8(n6476), .ADB9(n6475), 
           .ADB10(n6474), .ADB11(n6473), .ADB12(n6472), .ADB13(n6471), 
           .CEB(ram_a_buff_out_7__N_127), .OCEB(VCC_net), .CLKB(spi_clk_pos_derived_59), 
           .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), .CSB2(GND_net), 
           .RSTB(GND_net), .DOB0(n6579), .DOB1(n6580), .DOB2(n6581), 
           .DOB3(n6582), .DOB4(n6583), .DOB5(n6584), .DOB6(n6585), .DOB7(n6586));
    defparam mem0.DATA_WIDTH_A = 9;
    defparam mem0.DATA_WIDTH_B = 9;
    defparam mem0.REGMODE_A = "NOREG";
    defparam mem0.REGMODE_B = "NOREG";
    defparam mem0.RESETMODE = "SYNC";
    defparam mem0.ASYNC_RESET_RELEASE = "SYNC";
    defparam mem0.WRITEMODE_A = "READBEFOREWRITE";
    defparam mem0.WRITEMODE_B = "READBEFOREWRITE";
    defparam mem0.CSDECODE_A = "0b000";
    defparam mem0.CSDECODE_B = "0b000";
    defparam mem0.GSR = "DISABLED";
    defparam mem0.INITVAL_00 = "0x00000000000000000004108E7080840088A002F50E8930682004A731E02400C800006F00A000006F";
    defparam mem0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_02 = "0x00280002170100000437080011029300200002B7000000024A000000008000000000700000000070";
    defparam mem0.INITVAL_03 = "0x0602000073068820684416073000A4128B30888506020000731400105079004C0000EF1F44100213";
    defparam mem0.INITVAL_04 = "0x1D80110E93000E61F2631D80110E131D80110C930602000073068820604416073000A4128B308885";
    defparam mem0.INITVAL_05 = "0x11C911FEF710C93004F60EA630008710E931800110C130020000EB71FCE71DAE300EC1000071C023";
    defparam mem0.INITVAL_06 = "0x1FCD7136E31FCC705C2300E1100E91086900382000E9312CB21800110E1300C910382000C13134F1";
    defparam mem0.INITVAL_07 = "0x00EC100E41000A71E023000070EA03040A000E131D80110E93000670FC631D801106131D80110E13";
    defparam mem0.INITVAL_08 = "0x08E92184021849008C05022F700E130400610C93022610000714E371000000CB7100821FC671D4E3";
    defparam mem0.INITVAL_09 = "0x00E8508E821FCF7082E308E821800200006140231FCF70B8E308E921843E00E8508E92000F709063";
    defparam mem0.INITVAL_0A = "0x0009500E63188811089300A051D026102040049500263180011688317EC91FCF70B8E308E821803E";
    defparam mem0.INITVAL_0B = "0x10E1306020000730688206045060730000800A3717ECD1808110A13060200007306882180A114423";
    defparam mem0.INITVAL_0C = "0x0000800AB7180B114023000B601C63000E511A6300A85112881800116A83060061607308CA118881";
    defparam mem0.INITVAL_0D = "0x06006160731FCE601CE31804114E03060061407316EDD1808110A931008206006140730604514073";
    defparam mem0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000020000008002000000817EE1";
    defparam mem0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mem0.INIT_DATA = "STATIC";
    FD1P3AX i4312 (.D(n6486), .SP(ram_a_buff_out_7__N_127), .CK(spi_clk_pos_derived_59), 
            .Q(n6595));
    defparam i4312.GSR = "DISABLED";
    
endmodule
